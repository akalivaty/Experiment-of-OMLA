

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U559 ( .A(n749), .B(n748), .ZN(n762) );
  NOR2_X1 U560 ( .A1(n664), .A2(G651), .ZN(n675) );
  NOR2_X1 U561 ( .A1(n747), .A2(G2084), .ZN(n749) );
  NOR2_X1 U562 ( .A1(n664), .A2(n569), .ZN(n681) );
  XOR2_X1 U563 ( .A(n532), .B(KEYINPUT23), .Z(n526) );
  NOR2_X1 U564 ( .A1(n726), .A2(n1009), .ZN(n725) );
  AND2_X1 U565 ( .A1(n723), .A2(n722), .ZN(n726) );
  BUF_X1 U566 ( .A(n720), .Z(n747) );
  OR2_X1 U567 ( .A1(n720), .A2(n718), .ZN(n719) );
  XNOR2_X1 U568 ( .A(n542), .B(KEYINPUT64), .ZN(n720) );
  AND2_X1 U569 ( .A1(n548), .A2(n547), .ZN(n817) );
  OR2_X1 U570 ( .A1(n549), .A2(n580), .ZN(n544) );
  OR2_X1 U571 ( .A1(n564), .A2(n563), .ZN(n548) );
  AND2_X1 U572 ( .A1(n555), .A2(G2104), .ZN(n640) );
  INV_X1 U573 ( .A(G2105), .ZN(n555) );
  AND2_X1 U574 ( .A1(n762), .A2(G8), .ZN(n533) );
  NOR2_X1 U575 ( .A1(n750), .A2(G168), .ZN(n751) );
  XNOR2_X1 U576 ( .A(n535), .B(KEYINPUT30), .ZN(n750) );
  INV_X1 U577 ( .A(KEYINPUT98), .ZN(n538) );
  AND2_X1 U578 ( .A1(n817), .A2(G40), .ZN(n543) );
  AND2_X1 U579 ( .A1(G2104), .A2(G2105), .ZN(n912) );
  NAND2_X1 U580 ( .A1(n555), .A2(n560), .ZN(n554) );
  NAND2_X1 U581 ( .A1(n640), .A2(G101), .ZN(n532) );
  INV_X1 U582 ( .A(KEYINPUT90), .ZN(n748) );
  XNOR2_X1 U583 ( .A(n536), .B(KEYINPUT31), .ZN(n769) );
  XNOR2_X1 U584 ( .A(n751), .B(n538), .ZN(n537) );
  INV_X1 U585 ( .A(KEYINPUT29), .ZN(n736) );
  NAND2_X1 U586 ( .A1(n747), .A2(G8), .ZN(n795) );
  INV_X1 U587 ( .A(G1384), .ZN(n547) );
  XNOR2_X1 U588 ( .A(n540), .B(n546), .ZN(n539) );
  INV_X1 U589 ( .A(KEYINPUT102), .ZN(n546) );
  NOR2_X1 U590 ( .A1(n836), .A2(n556), .ZN(n837) );
  NAND2_X1 U591 ( .A1(n526), .A2(n581), .ZN(n549) );
  XOR2_X1 U592 ( .A(n717), .B(n716), .Z(n527) );
  OR2_X1 U593 ( .A1(G299), .A2(n734), .ZN(n528) );
  XOR2_X1 U594 ( .A(KEYINPUT99), .B(n753), .Z(n529) );
  XOR2_X1 U595 ( .A(KEYINPUT93), .B(n729), .Z(n530) );
  INV_X1 U596 ( .A(G2104), .ZN(n560) );
  XOR2_X1 U597 ( .A(n736), .B(KEYINPUT97), .Z(n531) );
  NAND2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n535) );
  INV_X1 U599 ( .A(n764), .ZN(n534) );
  NAND2_X1 U600 ( .A1(n537), .A2(n529), .ZN(n536) );
  NAND2_X1 U601 ( .A1(n539), .A2(n838), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n541), .A2(n837), .ZN(n540) );
  XNOR2_X1 U603 ( .A(n805), .B(KEYINPUT101), .ZN(n541) );
  NAND2_X1 U604 ( .A1(G160), .A2(n543), .ZN(n542) );
  XNOR2_X2 U605 ( .A(n544), .B(KEYINPUT65), .ZN(G160) );
  NAND2_X1 U606 ( .A1(n545), .A2(n852), .ZN(n853) );
  INV_X1 U607 ( .A(n548), .ZN(G164) );
  XNOR2_X1 U608 ( .A(n550), .B(n531), .ZN(n761) );
  NAND2_X1 U609 ( .A1(n551), .A2(n527), .ZN(n550) );
  XNOR2_X1 U610 ( .A(n552), .B(KEYINPUT96), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n553), .A2(n528), .ZN(n552) );
  INV_X1 U612 ( .A(n735), .ZN(n553) );
  NAND2_X1 U613 ( .A1(n916), .A2(G137), .ZN(n578) );
  XNOR2_X2 U614 ( .A(n554), .B(KEYINPUT17), .ZN(n916) );
  AND2_X1 U615 ( .A1(n849), .A2(n953), .ZN(n556) );
  NOR2_X1 U616 ( .A1(n721), .A2(n998), .ZN(n722) );
  INV_X1 U617 ( .A(KEYINPUT94), .ZN(n724) );
  INV_X1 U618 ( .A(n994), .ZN(n797) );
  INV_X1 U619 ( .A(G651), .ZN(n569) );
  NAND2_X1 U620 ( .A1(n593), .A2(n592), .ZN(n998) );
  NAND2_X1 U621 ( .A1(n640), .A2(G102), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n557), .B(KEYINPUT84), .ZN(n559) );
  NAND2_X1 U623 ( .A1(G138), .A2(n916), .ZN(n558) );
  NAND2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n564) );
  AND2_X1 U625 ( .A1(n560), .A2(G2105), .ZN(n633) );
  NAND2_X1 U626 ( .A1(G126), .A2(n633), .ZN(n562) );
  NAND2_X1 U627 ( .A1(G114), .A2(n912), .ZN(n561) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U629 ( .A1(G543), .A2(G651), .ZN(n677) );
  NAND2_X1 U630 ( .A1(n677), .A2(G89), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT4), .ZN(n567) );
  XOR2_X1 U632 ( .A(KEYINPUT0), .B(G543), .Z(n664) );
  NAND2_X1 U633 ( .A1(G76), .A2(n681), .ZN(n566) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(KEYINPUT5), .ZN(n576) );
  NAND2_X1 U636 ( .A1(n675), .A2(G51), .ZN(n573) );
  NOR2_X1 U637 ( .A1(G543), .A2(n569), .ZN(n570) );
  XOR2_X1 U638 ( .A(KEYINPUT1), .B(n570), .Z(n571) );
  XNOR2_X2 U639 ( .A(KEYINPUT66), .B(n571), .ZN(n678) );
  NAND2_X1 U640 ( .A1(G63), .A2(n678), .ZN(n572) );
  NAND2_X1 U641 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U642 ( .A(KEYINPUT6), .B(n574), .Z(n575) );
  NAND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n577), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U645 ( .A1(G113), .A2(n912), .ZN(n581) );
  NAND2_X1 U646 ( .A1(G125), .A2(n633), .ZN(n579) );
  NAND2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n580) );
  AND2_X1 U648 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U649 ( .A(G132), .ZN(G219) );
  INV_X1 U650 ( .A(G82), .ZN(G220) );
  INV_X1 U651 ( .A(G57), .ZN(G237) );
  XOR2_X1 U652 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U653 ( .A1(G7), .A2(G661), .ZN(n582) );
  XNOR2_X1 U654 ( .A(n582), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U655 ( .A(G223), .ZN(n854) );
  NAND2_X1 U656 ( .A1(n854), .A2(G567), .ZN(n583) );
  XNOR2_X1 U657 ( .A(n583), .B(KEYINPUT69), .ZN(n584) );
  XNOR2_X1 U658 ( .A(KEYINPUT11), .B(n584), .ZN(G234) );
  NAND2_X1 U659 ( .A1(n678), .A2(G56), .ZN(n585) );
  XOR2_X1 U660 ( .A(KEYINPUT14), .B(n585), .Z(n591) );
  NAND2_X1 U661 ( .A1(n677), .A2(G81), .ZN(n586) );
  XNOR2_X1 U662 ( .A(n586), .B(KEYINPUT12), .ZN(n588) );
  NAND2_X1 U663 ( .A1(G68), .A2(n681), .ZN(n587) );
  NAND2_X1 U664 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U665 ( .A(KEYINPUT13), .B(n589), .Z(n590) );
  NOR2_X1 U666 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U667 ( .A1(n675), .A2(G43), .ZN(n592) );
  INV_X1 U668 ( .A(n998), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n594), .A2(G860), .ZN(n595) );
  XNOR2_X1 U670 ( .A(KEYINPUT70), .B(n595), .ZN(G153) );
  NAND2_X1 U671 ( .A1(n675), .A2(G52), .ZN(n597) );
  NAND2_X1 U672 ( .A1(G64), .A2(n678), .ZN(n596) );
  NAND2_X1 U673 ( .A1(n597), .A2(n596), .ZN(n602) );
  NAND2_X1 U674 ( .A1(G90), .A2(n677), .ZN(n599) );
  NAND2_X1 U675 ( .A1(G77), .A2(n681), .ZN(n598) );
  NAND2_X1 U676 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U677 ( .A(KEYINPUT9), .B(n600), .Z(n601) );
  NOR2_X1 U678 ( .A1(n602), .A2(n601), .ZN(G171) );
  INV_X1 U679 ( .A(G868), .ZN(n622) );
  NOR2_X1 U680 ( .A1(n622), .A2(G171), .ZN(n603) );
  XNOR2_X1 U681 ( .A(n603), .B(KEYINPUT71), .ZN(n613) );
  NAND2_X1 U682 ( .A1(n677), .A2(G92), .ZN(n605) );
  NAND2_X1 U683 ( .A1(G66), .A2(n678), .ZN(n604) );
  NAND2_X1 U684 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U685 ( .A1(G79), .A2(n681), .ZN(n607) );
  NAND2_X1 U686 ( .A1(G54), .A2(n675), .ZN(n606) );
  NAND2_X1 U687 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U688 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U689 ( .A(KEYINPUT15), .B(n610), .Z(n611) );
  XNOR2_X2 U690 ( .A(KEYINPUT72), .B(n611), .ZN(n1009) );
  OR2_X1 U691 ( .A1(G868), .A2(n1009), .ZN(n612) );
  NAND2_X1 U692 ( .A1(n613), .A2(n612), .ZN(G284) );
  NAND2_X1 U693 ( .A1(G53), .A2(n675), .ZN(n614) );
  XNOR2_X1 U694 ( .A(n614), .B(KEYINPUT68), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n677), .A2(G91), .ZN(n616) );
  NAND2_X1 U696 ( .A1(G65), .A2(n678), .ZN(n615) );
  NAND2_X1 U697 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U698 ( .A1(G78), .A2(n681), .ZN(n617) );
  XNOR2_X1 U699 ( .A(KEYINPUT67), .B(n617), .ZN(n618) );
  NOR2_X1 U700 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n621), .A2(n620), .ZN(G299) );
  NOR2_X1 U702 ( .A1(G286), .A2(n622), .ZN(n624) );
  NOR2_X1 U703 ( .A1(G868), .A2(G299), .ZN(n623) );
  NOR2_X1 U704 ( .A1(n624), .A2(n623), .ZN(G297) );
  INV_X1 U705 ( .A(G559), .ZN(n625) );
  NOR2_X1 U706 ( .A1(G860), .A2(n625), .ZN(n626) );
  XNOR2_X1 U707 ( .A(KEYINPUT73), .B(n626), .ZN(n627) );
  NAND2_X1 U708 ( .A1(n627), .A2(n1009), .ZN(n628) );
  XNOR2_X1 U709 ( .A(n628), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U710 ( .A1(G868), .A2(n1009), .ZN(n629) );
  NOR2_X1 U711 ( .A1(G559), .A2(n629), .ZN(n630) );
  XNOR2_X1 U712 ( .A(n630), .B(KEYINPUT74), .ZN(n632) );
  NOR2_X1 U713 ( .A1(n998), .A2(G868), .ZN(n631) );
  NOR2_X1 U714 ( .A1(n632), .A2(n631), .ZN(G282) );
  NAND2_X1 U715 ( .A1(n633), .A2(G123), .ZN(n634) );
  XNOR2_X1 U716 ( .A(n634), .B(KEYINPUT18), .ZN(n636) );
  NAND2_X1 U717 ( .A1(G135), .A2(n916), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U719 ( .A(n637), .B(KEYINPUT75), .ZN(n639) );
  NAND2_X1 U720 ( .A1(G111), .A2(n912), .ZN(n638) );
  NAND2_X1 U721 ( .A1(n639), .A2(n638), .ZN(n643) );
  BUF_X1 U722 ( .A(n640), .Z(n915) );
  NAND2_X1 U723 ( .A1(n915), .A2(G99), .ZN(n641) );
  XOR2_X1 U724 ( .A(KEYINPUT76), .B(n641), .Z(n642) );
  NOR2_X1 U725 ( .A1(n643), .A2(n642), .ZN(n948) );
  XNOR2_X1 U726 ( .A(G2096), .B(n948), .ZN(n645) );
  INV_X1 U727 ( .A(G2100), .ZN(n644) );
  NAND2_X1 U728 ( .A1(n645), .A2(n644), .ZN(G156) );
  NAND2_X1 U729 ( .A1(G559), .A2(n1009), .ZN(n695) );
  XNOR2_X1 U730 ( .A(n998), .B(n695), .ZN(n646) );
  NOR2_X1 U731 ( .A1(n646), .A2(G860), .ZN(n653) );
  NAND2_X1 U732 ( .A1(n675), .A2(G55), .ZN(n648) );
  NAND2_X1 U733 ( .A1(G67), .A2(n678), .ZN(n647) );
  NAND2_X1 U734 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U735 ( .A1(G93), .A2(n677), .ZN(n650) );
  NAND2_X1 U736 ( .A1(G80), .A2(n681), .ZN(n649) );
  NAND2_X1 U737 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U738 ( .A1(n652), .A2(n651), .ZN(n690) );
  XNOR2_X1 U739 ( .A(n653), .B(n690), .ZN(G145) );
  AND2_X1 U740 ( .A1(G60), .A2(n678), .ZN(n657) );
  NAND2_X1 U741 ( .A1(G85), .A2(n677), .ZN(n655) );
  NAND2_X1 U742 ( .A1(G72), .A2(n681), .ZN(n654) );
  NAND2_X1 U743 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U744 ( .A1(n657), .A2(n656), .ZN(n659) );
  NAND2_X1 U745 ( .A1(n675), .A2(G47), .ZN(n658) );
  NAND2_X1 U746 ( .A1(n659), .A2(n658), .ZN(G290) );
  NAND2_X1 U747 ( .A1(G49), .A2(n675), .ZN(n661) );
  NAND2_X1 U748 ( .A1(G74), .A2(G651), .ZN(n660) );
  NAND2_X1 U749 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U750 ( .A1(n678), .A2(n662), .ZN(n663) );
  XOR2_X1 U751 ( .A(KEYINPUT77), .B(n663), .Z(n666) );
  NAND2_X1 U752 ( .A1(n664), .A2(G87), .ZN(n665) );
  NAND2_X1 U753 ( .A1(n666), .A2(n665), .ZN(G288) );
  NAND2_X1 U754 ( .A1(G88), .A2(n677), .ZN(n667) );
  XNOR2_X1 U755 ( .A(n667), .B(KEYINPUT80), .ZN(n670) );
  NAND2_X1 U756 ( .A1(G50), .A2(n675), .ZN(n668) );
  XOR2_X1 U757 ( .A(KEYINPUT79), .B(n668), .Z(n669) );
  NAND2_X1 U758 ( .A1(n670), .A2(n669), .ZN(n674) );
  NAND2_X1 U759 ( .A1(n681), .A2(G75), .ZN(n672) );
  NAND2_X1 U760 ( .A1(G62), .A2(n678), .ZN(n671) );
  NAND2_X1 U761 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U762 ( .A1(n674), .A2(n673), .ZN(G166) );
  NAND2_X1 U763 ( .A1(G48), .A2(n675), .ZN(n676) );
  XNOR2_X1 U764 ( .A(n676), .B(KEYINPUT78), .ZN(n686) );
  NAND2_X1 U765 ( .A1(n677), .A2(G86), .ZN(n680) );
  NAND2_X1 U766 ( .A1(G61), .A2(n678), .ZN(n679) );
  NAND2_X1 U767 ( .A1(n680), .A2(n679), .ZN(n684) );
  NAND2_X1 U768 ( .A1(n681), .A2(G73), .ZN(n682) );
  XOR2_X1 U769 ( .A(KEYINPUT2), .B(n682), .Z(n683) );
  NOR2_X1 U770 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U771 ( .A1(n686), .A2(n685), .ZN(G305) );
  NOR2_X1 U772 ( .A1(G868), .A2(n690), .ZN(n687) );
  XNOR2_X1 U773 ( .A(n687), .B(KEYINPUT81), .ZN(n698) );
  XNOR2_X1 U774 ( .A(KEYINPUT19), .B(G290), .ZN(n688) );
  XNOR2_X1 U775 ( .A(n688), .B(n998), .ZN(n689) );
  XNOR2_X1 U776 ( .A(n690), .B(n689), .ZN(n692) );
  XNOR2_X1 U777 ( .A(G288), .B(G166), .ZN(n691) );
  XNOR2_X1 U778 ( .A(n692), .B(n691), .ZN(n693) );
  XOR2_X1 U779 ( .A(n693), .B(G305), .Z(n694) );
  XNOR2_X1 U780 ( .A(G299), .B(n694), .ZN(n926) );
  XNOR2_X1 U781 ( .A(n926), .B(n695), .ZN(n696) );
  NAND2_X1 U782 ( .A1(G868), .A2(n696), .ZN(n697) );
  NAND2_X1 U783 ( .A1(n698), .A2(n697), .ZN(G295) );
  NAND2_X1 U784 ( .A1(G2078), .A2(G2084), .ZN(n699) );
  XOR2_X1 U785 ( .A(KEYINPUT20), .B(n699), .Z(n700) );
  NAND2_X1 U786 ( .A1(G2090), .A2(n700), .ZN(n701) );
  XNOR2_X1 U787 ( .A(KEYINPUT21), .B(n701), .ZN(n702) );
  NAND2_X1 U788 ( .A1(n702), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U789 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U790 ( .A1(G69), .A2(G120), .ZN(n703) );
  NOR2_X1 U791 ( .A1(G237), .A2(n703), .ZN(n704) );
  NAND2_X1 U792 ( .A1(G108), .A2(n704), .ZN(n861) );
  NAND2_X1 U793 ( .A1(n861), .A2(G567), .ZN(n710) );
  NOR2_X1 U794 ( .A1(G220), .A2(G219), .ZN(n705) );
  XOR2_X1 U795 ( .A(KEYINPUT22), .B(n705), .Z(n706) );
  NOR2_X1 U796 ( .A1(G218), .A2(n706), .ZN(n707) );
  NAND2_X1 U797 ( .A1(G96), .A2(n707), .ZN(n862) );
  NAND2_X1 U798 ( .A1(G2106), .A2(n862), .ZN(n708) );
  XNOR2_X1 U799 ( .A(KEYINPUT82), .B(n708), .ZN(n709) );
  NAND2_X1 U800 ( .A1(n710), .A2(n709), .ZN(n864) );
  NAND2_X1 U801 ( .A1(G661), .A2(G483), .ZN(n711) );
  NOR2_X1 U802 ( .A1(n864), .A2(n711), .ZN(n712) );
  XOR2_X1 U803 ( .A(KEYINPUT83), .B(n712), .Z(n859) );
  NAND2_X1 U804 ( .A1(n859), .A2(G36), .ZN(G176) );
  INV_X1 U805 ( .A(G171), .ZN(G301) );
  INV_X1 U806 ( .A(G166), .ZN(G303) );
  XOR2_X1 U807 ( .A(KEYINPUT28), .B(KEYINPUT92), .Z(n717) );
  INV_X1 U808 ( .A(n720), .ZN(n738) );
  NAND2_X1 U809 ( .A1(G2072), .A2(n738), .ZN(n713) );
  XOR2_X1 U810 ( .A(KEYINPUT27), .B(n713), .Z(n715) );
  NAND2_X1 U811 ( .A1(n747), .A2(G1956), .ZN(n714) );
  NAND2_X1 U812 ( .A1(n715), .A2(n714), .ZN(n734) );
  NAND2_X1 U813 ( .A1(n734), .A2(G299), .ZN(n716) );
  INV_X1 U814 ( .A(G1996), .ZN(n718) );
  XNOR2_X1 U815 ( .A(n719), .B(KEYINPUT26), .ZN(n723) );
  AND2_X1 U816 ( .A1(n720), .A2(G1341), .ZN(n721) );
  XNOR2_X1 U817 ( .A(n725), .B(n724), .ZN(n732) );
  NAND2_X1 U818 ( .A1(n726), .A2(n1009), .ZN(n730) );
  NAND2_X1 U819 ( .A1(G2067), .A2(n738), .ZN(n728) );
  NAND2_X1 U820 ( .A1(n747), .A2(G1348), .ZN(n727) );
  NAND2_X1 U821 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U822 ( .A1(n730), .A2(n530), .ZN(n731) );
  NAND2_X1 U823 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U824 ( .A(n733), .B(KEYINPUT95), .ZN(n735) );
  XNOR2_X1 U825 ( .A(KEYINPUT25), .B(G2078), .ZN(n980) );
  NAND2_X1 U826 ( .A1(n738), .A2(n980), .ZN(n737) );
  XNOR2_X1 U827 ( .A(n737), .B(KEYINPUT91), .ZN(n740) );
  NOR2_X1 U828 ( .A1(n738), .A2(G1961), .ZN(n739) );
  NOR2_X1 U829 ( .A1(n740), .A2(n739), .ZN(n752) );
  OR2_X1 U830 ( .A1(n752), .A2(G301), .ZN(n767) );
  NOR2_X1 U831 ( .A1(n747), .A2(G2090), .ZN(n742) );
  NOR2_X1 U832 ( .A1(G1971), .A2(n795), .ZN(n741) );
  NOR2_X1 U833 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U834 ( .A1(G303), .A2(n743), .ZN(n754) );
  INV_X1 U835 ( .A(n754), .ZN(n744) );
  OR2_X1 U836 ( .A1(n744), .A2(G286), .ZN(n745) );
  AND2_X1 U837 ( .A1(n745), .A2(G8), .ZN(n755) );
  AND2_X1 U838 ( .A1(n767), .A2(n755), .ZN(n746) );
  NAND2_X1 U839 ( .A1(n761), .A2(n746), .ZN(n758) );
  NOR2_X1 U840 ( .A1(G1966), .A2(n795), .ZN(n764) );
  NAND2_X1 U841 ( .A1(n752), .A2(G301), .ZN(n753) );
  NAND2_X1 U842 ( .A1(n769), .A2(n754), .ZN(n756) );
  NAND2_X1 U843 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U844 ( .A1(n758), .A2(n757), .ZN(n760) );
  INV_X1 U845 ( .A(KEYINPUT32), .ZN(n759) );
  XNOR2_X1 U846 ( .A(n760), .B(n759), .ZN(n786) );
  INV_X1 U847 ( .A(n762), .ZN(n763) );
  AND2_X1 U848 ( .A1(n763), .A2(G8), .ZN(n765) );
  OR2_X1 U849 ( .A1(n765), .A2(n764), .ZN(n770) );
  INV_X1 U850 ( .A(n770), .ZN(n766) );
  AND2_X1 U851 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U852 ( .A1(n761), .A2(n768), .ZN(n785) );
  OR2_X1 U853 ( .A1(n770), .A2(n769), .ZN(n783) );
  AND2_X1 U854 ( .A1(n785), .A2(n783), .ZN(n771) );
  NAND2_X1 U855 ( .A1(n786), .A2(n771), .ZN(n774) );
  NOR2_X1 U856 ( .A1(G2090), .A2(G303), .ZN(n772) );
  NAND2_X1 U857 ( .A1(G8), .A2(n772), .ZN(n773) );
  NAND2_X1 U858 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U859 ( .A1(n775), .A2(n795), .ZN(n777) );
  INV_X1 U860 ( .A(KEYINPUT100), .ZN(n776) );
  XNOR2_X1 U861 ( .A(n777), .B(n776), .ZN(n804) );
  NOR2_X1 U862 ( .A1(G1981), .A2(G305), .ZN(n778) );
  XNOR2_X1 U863 ( .A(n778), .B(KEYINPUT24), .ZN(n779) );
  XNOR2_X1 U864 ( .A(n779), .B(KEYINPUT89), .ZN(n780) );
  OR2_X1 U865 ( .A1(n780), .A2(n795), .ZN(n802) );
  NAND2_X1 U866 ( .A1(G1976), .A2(G288), .ZN(n1003) );
  INV_X1 U867 ( .A(n795), .ZN(n781) );
  NAND2_X1 U868 ( .A1(n1003), .A2(n781), .ZN(n789) );
  INV_X1 U869 ( .A(n789), .ZN(n782) );
  AND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n784) );
  AND2_X1 U871 ( .A1(n785), .A2(n784), .ZN(n787) );
  AND2_X1 U872 ( .A1(n787), .A2(n786), .ZN(n793) );
  NOR2_X1 U873 ( .A1(G1976), .A2(G288), .ZN(n794) );
  NOR2_X1 U874 ( .A1(G1971), .A2(G303), .ZN(n788) );
  NOR2_X1 U875 ( .A1(n794), .A2(n788), .ZN(n1011) );
  OR2_X1 U876 ( .A1(n789), .A2(n1011), .ZN(n791) );
  INV_X1 U877 ( .A(KEYINPUT33), .ZN(n790) );
  NAND2_X1 U878 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U879 ( .A1(n793), .A2(n792), .ZN(n800) );
  NAND2_X1 U880 ( .A1(n794), .A2(KEYINPUT33), .ZN(n796) );
  NOR2_X1 U881 ( .A1(n796), .A2(n795), .ZN(n798) );
  XOR2_X1 U882 ( .A(G1981), .B(G305), .Z(n994) );
  OR2_X1 U883 ( .A1(n798), .A2(n797), .ZN(n799) );
  OR2_X1 U884 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U885 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U886 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U887 ( .A(G2067), .B(KEYINPUT37), .Z(n806) );
  XNOR2_X1 U888 ( .A(KEYINPUT85), .B(n806), .ZN(n847) );
  NAND2_X1 U889 ( .A1(G104), .A2(n915), .ZN(n808) );
  NAND2_X1 U890 ( .A1(G140), .A2(n916), .ZN(n807) );
  NAND2_X1 U891 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U892 ( .A(KEYINPUT34), .B(n809), .ZN(n814) );
  NAND2_X1 U893 ( .A1(G128), .A2(n633), .ZN(n811) );
  NAND2_X1 U894 ( .A1(G116), .A2(n912), .ZN(n810) );
  NAND2_X1 U895 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U896 ( .A(KEYINPUT35), .B(n812), .Z(n813) );
  NOR2_X1 U897 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U898 ( .A(KEYINPUT36), .B(n815), .ZN(n909) );
  NOR2_X1 U899 ( .A1(n847), .A2(n909), .ZN(n949) );
  NAND2_X1 U900 ( .A1(G160), .A2(G40), .ZN(n816) );
  NOR2_X1 U901 ( .A1(n817), .A2(n816), .ZN(n849) );
  NAND2_X1 U902 ( .A1(n949), .A2(n849), .ZN(n818) );
  XNOR2_X1 U903 ( .A(n818), .B(KEYINPUT86), .ZN(n846) );
  INV_X1 U904 ( .A(n846), .ZN(n836) );
  NAND2_X1 U905 ( .A1(G119), .A2(n633), .ZN(n820) );
  NAND2_X1 U906 ( .A1(G131), .A2(n916), .ZN(n819) );
  NAND2_X1 U907 ( .A1(n820), .A2(n819), .ZN(n823) );
  NAND2_X1 U908 ( .A1(G95), .A2(n915), .ZN(n821) );
  XNOR2_X1 U909 ( .A(KEYINPUT87), .B(n821), .ZN(n822) );
  NOR2_X1 U910 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U911 ( .A1(n912), .A2(G107), .ZN(n824) );
  NAND2_X1 U912 ( .A1(n825), .A2(n824), .ZN(n901) );
  NAND2_X1 U913 ( .A1(G1991), .A2(n901), .ZN(n826) );
  XNOR2_X1 U914 ( .A(n826), .B(KEYINPUT88), .ZN(n835) );
  NAND2_X1 U915 ( .A1(G129), .A2(n633), .ZN(n828) );
  NAND2_X1 U916 ( .A1(G141), .A2(n916), .ZN(n827) );
  NAND2_X1 U917 ( .A1(n828), .A2(n827), .ZN(n831) );
  NAND2_X1 U918 ( .A1(n915), .A2(G105), .ZN(n829) );
  XOR2_X1 U919 ( .A(KEYINPUT38), .B(n829), .Z(n830) );
  NOR2_X1 U920 ( .A1(n831), .A2(n830), .ZN(n833) );
  NAND2_X1 U921 ( .A1(n912), .A2(G117), .ZN(n832) );
  NAND2_X1 U922 ( .A1(n833), .A2(n832), .ZN(n903) );
  NAND2_X1 U923 ( .A1(G1996), .A2(n903), .ZN(n834) );
  NAND2_X1 U924 ( .A1(n835), .A2(n834), .ZN(n953) );
  XNOR2_X1 U925 ( .A(G1986), .B(G290), .ZN(n1005) );
  NAND2_X1 U926 ( .A1(n849), .A2(n1005), .ZN(n838) );
  NOR2_X1 U927 ( .A1(G1996), .A2(n903), .ZN(n839) );
  XOR2_X1 U928 ( .A(KEYINPUT103), .B(n839), .Z(n964) );
  NOR2_X1 U929 ( .A1(G1986), .A2(G290), .ZN(n840) );
  NOR2_X1 U930 ( .A1(G1991), .A2(n901), .ZN(n947) );
  NOR2_X1 U931 ( .A1(n840), .A2(n947), .ZN(n841) );
  NOR2_X1 U932 ( .A1(n953), .A2(n841), .ZN(n842) );
  NOR2_X1 U933 ( .A1(n964), .A2(n842), .ZN(n843) );
  XNOR2_X1 U934 ( .A(n843), .B(KEYINPUT39), .ZN(n844) );
  XNOR2_X1 U935 ( .A(n844), .B(KEYINPUT104), .ZN(n845) );
  NAND2_X1 U936 ( .A1(n846), .A2(n845), .ZN(n848) );
  NAND2_X1 U937 ( .A1(n847), .A2(n909), .ZN(n954) );
  NAND2_X1 U938 ( .A1(n848), .A2(n954), .ZN(n850) );
  NAND2_X1 U939 ( .A1(n850), .A2(n849), .ZN(n851) );
  XOR2_X1 U940 ( .A(KEYINPUT105), .B(n851), .Z(n852) );
  XNOR2_X1 U941 ( .A(n853), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U942 ( .A1(G2106), .A2(n854), .ZN(G217) );
  NAND2_X1 U943 ( .A1(G15), .A2(G2), .ZN(n856) );
  INV_X1 U944 ( .A(G661), .ZN(n855) );
  NOR2_X1 U945 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U946 ( .A(n857), .B(KEYINPUT107), .ZN(G259) );
  NAND2_X1 U947 ( .A1(G3), .A2(G1), .ZN(n858) );
  XNOR2_X1 U948 ( .A(KEYINPUT108), .B(n858), .ZN(n860) );
  NAND2_X1 U949 ( .A1(n860), .A2(n859), .ZN(G188) );
  INV_X1 U951 ( .A(G120), .ZN(G236) );
  INV_X1 U952 ( .A(G96), .ZN(G221) );
  INV_X1 U953 ( .A(G69), .ZN(G235) );
  NOR2_X1 U954 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U955 ( .A(n863), .B(KEYINPUT109), .ZN(G261) );
  INV_X1 U956 ( .A(G261), .ZN(G325) );
  INV_X1 U957 ( .A(n864), .ZN(G319) );
  XOR2_X1 U958 ( .A(G2096), .B(KEYINPUT43), .Z(n866) );
  XNOR2_X1 U959 ( .A(G2090), .B(G2678), .ZN(n865) );
  XNOR2_X1 U960 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U961 ( .A(n867), .B(KEYINPUT110), .Z(n869) );
  XNOR2_X1 U962 ( .A(G2067), .B(G2072), .ZN(n868) );
  XNOR2_X1 U963 ( .A(n869), .B(n868), .ZN(n873) );
  XOR2_X1 U964 ( .A(KEYINPUT42), .B(G2100), .Z(n871) );
  XNOR2_X1 U965 ( .A(G2078), .B(G2084), .ZN(n870) );
  XNOR2_X1 U966 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U967 ( .A(n873), .B(n872), .ZN(G227) );
  XOR2_X1 U968 ( .A(G1961), .B(G1956), .Z(n875) );
  XNOR2_X1 U969 ( .A(G1986), .B(G1966), .ZN(n874) );
  XNOR2_X1 U970 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U971 ( .A(n876), .B(G2474), .Z(n878) );
  XNOR2_X1 U972 ( .A(G1976), .B(G1971), .ZN(n877) );
  XNOR2_X1 U973 ( .A(n878), .B(n877), .ZN(n882) );
  XOR2_X1 U974 ( .A(KEYINPUT41), .B(G1981), .Z(n880) );
  XNOR2_X1 U975 ( .A(G1996), .B(G1991), .ZN(n879) );
  XNOR2_X1 U976 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U977 ( .A(n882), .B(n881), .ZN(G229) );
  NAND2_X1 U978 ( .A1(n912), .A2(G112), .ZN(n883) );
  XOR2_X1 U979 ( .A(KEYINPUT111), .B(n883), .Z(n885) );
  NAND2_X1 U980 ( .A1(n915), .A2(G100), .ZN(n884) );
  NAND2_X1 U981 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U982 ( .A(KEYINPUT112), .B(n886), .ZN(n891) );
  NAND2_X1 U983 ( .A1(n633), .A2(G124), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n887), .B(KEYINPUT44), .ZN(n889) );
  NAND2_X1 U985 ( .A1(G136), .A2(n916), .ZN(n888) );
  NAND2_X1 U986 ( .A1(n889), .A2(n888), .ZN(n890) );
  NOR2_X1 U987 ( .A1(n891), .A2(n890), .ZN(G162) );
  NAND2_X1 U988 ( .A1(G103), .A2(n915), .ZN(n893) );
  NAND2_X1 U989 ( .A1(G139), .A2(n916), .ZN(n892) );
  NAND2_X1 U990 ( .A1(n893), .A2(n892), .ZN(n899) );
  NAND2_X1 U991 ( .A1(G127), .A2(n633), .ZN(n895) );
  NAND2_X1 U992 ( .A1(G115), .A2(n912), .ZN(n894) );
  NAND2_X1 U993 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U994 ( .A(KEYINPUT113), .B(n896), .ZN(n897) );
  XNOR2_X1 U995 ( .A(KEYINPUT47), .B(n897), .ZN(n898) );
  NOR2_X1 U996 ( .A1(n899), .A2(n898), .ZN(n956) );
  XOR2_X1 U997 ( .A(G164), .B(n956), .Z(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n905) );
  XOR2_X1 U999 ( .A(G160), .B(G162), .Z(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n911) );
  XOR2_X1 U1002 ( .A(KEYINPUT46), .B(KEYINPUT114), .Z(n907) );
  XNOR2_X1 U1003 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(n911), .B(n910), .ZN(n924) );
  NAND2_X1 U1007 ( .A1(G130), .A2(n633), .ZN(n914) );
  NAND2_X1 U1008 ( .A1(G118), .A2(n912), .ZN(n913) );
  NAND2_X1 U1009 ( .A1(n914), .A2(n913), .ZN(n921) );
  NAND2_X1 U1010 ( .A1(G106), .A2(n915), .ZN(n918) );
  NAND2_X1 U1011 ( .A1(G142), .A2(n916), .ZN(n917) );
  NAND2_X1 U1012 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1013 ( .A(KEYINPUT45), .B(n919), .Z(n920) );
  NOR2_X1 U1014 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1015 ( .A(n948), .B(n922), .ZN(n923) );
  XNOR2_X1 U1016 ( .A(n924), .B(n923), .ZN(n925) );
  NOR2_X1 U1017 ( .A1(G37), .A2(n925), .ZN(G395) );
  XNOR2_X1 U1018 ( .A(G286), .B(G301), .ZN(n927) );
  XNOR2_X1 U1019 ( .A(n927), .B(n926), .ZN(n928) );
  XNOR2_X1 U1020 ( .A(n928), .B(n1009), .ZN(n929) );
  NOR2_X1 U1021 ( .A1(G37), .A2(n929), .ZN(G397) );
  XOR2_X1 U1022 ( .A(G2443), .B(G2427), .Z(n931) );
  XNOR2_X1 U1023 ( .A(G2438), .B(G2454), .ZN(n930) );
  XNOR2_X1 U1024 ( .A(n931), .B(n930), .ZN(n932) );
  XOR2_X1 U1025 ( .A(n932), .B(G2435), .Z(n934) );
  XNOR2_X1 U1026 ( .A(G1341), .B(G1348), .ZN(n933) );
  XNOR2_X1 U1027 ( .A(n934), .B(n933), .ZN(n938) );
  XOR2_X1 U1028 ( .A(G2430), .B(G2446), .Z(n936) );
  XNOR2_X1 U1029 ( .A(KEYINPUT106), .B(G2451), .ZN(n935) );
  XNOR2_X1 U1030 ( .A(n936), .B(n935), .ZN(n937) );
  XOR2_X1 U1031 ( .A(n938), .B(n937), .Z(n939) );
  NAND2_X1 U1032 ( .A1(G14), .A2(n939), .ZN(n945) );
  NAND2_X1 U1033 ( .A1(G319), .A2(n945), .ZN(n942) );
  NOR2_X1 U1034 ( .A1(G227), .A2(G229), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(KEYINPUT49), .B(n940), .ZN(n941) );
  NOR2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n944) );
  NOR2_X1 U1037 ( .A1(G395), .A2(G397), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(G225) );
  INV_X1 U1039 ( .A(G225), .ZN(G308) );
  INV_X1 U1040 ( .A(G108), .ZN(G238) );
  INV_X1 U1041 ( .A(n945), .ZN(G401) );
  XOR2_X1 U1042 ( .A(G2084), .B(G160), .Z(n946) );
  NOR2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n951) );
  NOR2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(KEYINPUT116), .B(n952), .ZN(n969) );
  INV_X1 U1047 ( .A(n953), .ZN(n955) );
  NAND2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n961) );
  XOR2_X1 U1049 ( .A(G2072), .B(n956), .Z(n958) );
  XOR2_X1 U1050 ( .A(G164), .B(G2078), .Z(n957) );
  NOR2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1052 ( .A(KEYINPUT50), .B(n959), .Z(n960) );
  NOR2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n967) );
  XNOR2_X1 U1054 ( .A(G2090), .B(G162), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(n962), .B(KEYINPUT117), .ZN(n963) );
  NOR2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1057 ( .A(KEYINPUT51), .B(n965), .Z(n966) );
  NAND2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1059 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1060 ( .A(KEYINPUT52), .B(n970), .ZN(n971) );
  INV_X1 U1061 ( .A(KEYINPUT55), .ZN(n990) );
  NAND2_X1 U1062 ( .A1(n971), .A2(n990), .ZN(n972) );
  NAND2_X1 U1063 ( .A1(n972), .A2(G29), .ZN(n1053) );
  XNOR2_X1 U1064 ( .A(G2090), .B(G35), .ZN(n985) );
  XNOR2_X1 U1065 ( .A(G2067), .B(G26), .ZN(n974) );
  XNOR2_X1 U1066 ( .A(G33), .B(G2072), .ZN(n973) );
  NOR2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n979) );
  XOR2_X1 U1068 ( .A(G1991), .B(G25), .Z(n975) );
  NAND2_X1 U1069 ( .A1(n975), .A2(G28), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(G32), .B(G1996), .ZN(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n982) );
  XOR2_X1 U1073 ( .A(G27), .B(n980), .Z(n981) );
  NOR2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(KEYINPUT53), .B(n983), .ZN(n984) );
  NOR2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n988) );
  XOR2_X1 U1077 ( .A(G2084), .B(KEYINPUT54), .Z(n986) );
  XNOR2_X1 U1078 ( .A(G34), .B(n986), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(n990), .B(n989), .ZN(n992) );
  INV_X1 U1081 ( .A(G29), .ZN(n991) );
  NAND2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1083 ( .A1(G11), .A2(n993), .ZN(n1051) );
  XNOR2_X1 U1084 ( .A(G16), .B(KEYINPUT56), .ZN(n1020) );
  XNOR2_X1 U1085 ( .A(G1966), .B(G168), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(n996), .B(KEYINPUT118), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(KEYINPUT57), .B(n997), .ZN(n1018) );
  XNOR2_X1 U1089 ( .A(n998), .B(G1341), .ZN(n1016) );
  XNOR2_X1 U1090 ( .A(G1956), .B(KEYINPUT120), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(n999), .B(G299), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(G1961), .B(G301), .ZN(n1000) );
  NOR2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(G1971), .A2(G303), .ZN(n1002) );
  NAND2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1013) );
  XOR2_X1 U1098 ( .A(G1348), .B(KEYINPUT119), .Z(n1008) );
  XNOR2_X1 U1099 ( .A(n1009), .B(n1008), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(KEYINPUT121), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1049) );
  XOR2_X1 U1106 ( .A(G16), .B(KEYINPUT122), .Z(n1047) );
  XOR2_X1 U1107 ( .A(G1986), .B(KEYINPUT126), .Z(n1021) );
  XNOR2_X1 U1108 ( .A(G24), .B(n1021), .ZN(n1025) );
  XNOR2_X1 U1109 ( .A(G1976), .B(G23), .ZN(n1023) );
  XNOR2_X1 U1110 ( .A(G1971), .B(G22), .ZN(n1022) );
  NOR2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1113 ( .A(n1026), .B(KEYINPUT127), .ZN(n1027) );
  XNOR2_X1 U1114 ( .A(KEYINPUT58), .B(n1027), .ZN(n1031) );
  XNOR2_X1 U1115 ( .A(G1966), .B(G21), .ZN(n1029) );
  XNOR2_X1 U1116 ( .A(G5), .B(G1961), .ZN(n1028) );
  NOR2_X1 U1117 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1044) );
  XOR2_X1 U1119 ( .A(KEYINPUT124), .B(G4), .Z(n1033) );
  XNOR2_X1 U1120 ( .A(G1348), .B(KEYINPUT59), .ZN(n1032) );
  XNOR2_X1 U1121 ( .A(n1033), .B(n1032), .ZN(n1040) );
  XOR2_X1 U1122 ( .A(G1341), .B(G19), .Z(n1037) );
  XNOR2_X1 U1123 ( .A(G1981), .B(G6), .ZN(n1035) );
  XNOR2_X1 U1124 ( .A(G20), .B(G1956), .ZN(n1034) );
  NOR2_X1 U1125 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1126 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XOR2_X1 U1127 ( .A(KEYINPUT123), .B(n1038), .Z(n1039) );
  NOR2_X1 U1128 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XNOR2_X1 U1129 ( .A(KEYINPUT125), .B(n1041), .ZN(n1042) );
  XNOR2_X1 U1130 ( .A(KEYINPUT60), .B(n1042), .ZN(n1043) );
  NOR2_X1 U1131 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  XNOR2_X1 U1132 ( .A(n1045), .B(KEYINPUT61), .ZN(n1046) );
  NAND2_X1 U1133 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  NAND2_X1 U1134 ( .A1(n1049), .A2(n1048), .ZN(n1050) );
  NOR2_X1 U1135 ( .A1(n1051), .A2(n1050), .ZN(n1052) );
  NAND2_X1 U1136 ( .A1(n1053), .A2(n1052), .ZN(n1054) );
  XOR2_X1 U1137 ( .A(KEYINPUT62), .B(n1054), .Z(G311) );
  INV_X1 U1138 ( .A(G311), .ZN(G150) );
endmodule

