//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1228, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT0), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G97), .A2(G257), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  OAI21_X1  g0010(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT66), .Z(new_n213));
  AOI211_X1 g0013(.A(new_n211), .B(new_n213), .C1(G77), .C2(G244), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AND2_X1   g0019(.A1(G107), .A2(G264), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n203), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT65), .ZN(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n207), .B(new_n222), .C1(new_n226), .C2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G264), .ZN(new_n235));
  INV_X1    g0035(.A(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n233), .B(new_n237), .Z(G358));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT67), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G97), .B(G107), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(KEYINPUT3), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G1698), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G222), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G223), .A2(G1698), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n251), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n255), .B(new_n256), .C1(G77), .C2(new_n251), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G226), .ZN(new_n263));
  INV_X1    g0063(.A(new_n256), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n259), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n257), .B(new_n262), .C1(new_n263), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G200), .ZN(new_n267));
  INV_X1    g0067(.A(G190), .ZN(new_n268));
  OAI21_X1  g0068(.A(KEYINPUT68), .B1(new_n203), .B2(new_n248), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT68), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n270), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n269), .A2(new_n223), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT8), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(new_n215), .B2(KEYINPUT69), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT69), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(KEYINPUT8), .A3(G58), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n224), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G150), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NOR3_X1   g0082(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n283));
  OAI22_X1  g0083(.A1(new_n280), .A2(new_n282), .B1(new_n283), .B2(new_n224), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n272), .B1(new_n279), .B2(new_n284), .ZN(new_n285));
  OR2_X1    g0085(.A1(new_n285), .A2(KEYINPUT70), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(KEYINPUT70), .ZN(new_n287));
  INV_X1    g0087(.A(G50), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n258), .A2(G13), .A3(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n286), .A2(new_n287), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n272), .B1(new_n258), .B2(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n291), .B1(new_n288), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT9), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n267), .B1(new_n268), .B2(new_n266), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n294), .A2(new_n295), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT10), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n266), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT71), .B1(new_n266), .B2(G179), .ZN(new_n303));
  OR3_X1    g0103(.A1(new_n266), .A2(KEYINPUT71), .A3(G179), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n294), .A2(new_n302), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  AND2_X1   g0105(.A1(KEYINPUT3), .A2(G33), .ZN(new_n306));
  NOR2_X1   g0106(.A1(KEYINPUT3), .A2(G33), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(new_n216), .B2(G1698), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n263), .A2(new_n252), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n309), .A2(new_n310), .B1(G33), .B2(G97), .ZN(new_n311));
  OAI221_X1 g0111(.A(new_n262), .B1(new_n210), .B2(new_n265), .C1(new_n311), .C2(new_n264), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n312), .A2(KEYINPUT13), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(KEYINPUT13), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT14), .B1(new_n315), .B2(new_n301), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(G179), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n312), .B(KEYINPUT13), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT14), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n318), .A2(new_n319), .A3(G169), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n316), .A2(new_n317), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n281), .A2(G50), .ZN(new_n322));
  INV_X1    g0122(.A(G77), .ZN(new_n323));
  OAI221_X1 g0123(.A(new_n322), .B1(new_n224), .B2(G68), .C1(new_n323), .C2(new_n278), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n324), .A2(new_n272), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n325), .A2(KEYINPUT11), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(KEYINPUT11), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n290), .A2(new_n209), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n328), .B(KEYINPUT12), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n292), .A2(G68), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n326), .A2(new_n327), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n321), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(G200), .B1(new_n313), .B2(new_n314), .ZN(new_n333));
  INV_X1    g0133(.A(new_n331), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n333), .B(new_n334), .C1(new_n268), .C2(new_n318), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT72), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n331), .B1(new_n315), .B2(G190), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT72), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(new_n338), .A3(new_n333), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n300), .A2(new_n305), .A3(new_n332), .A4(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT17), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT75), .ZN(new_n343));
  OAI211_X1 g0143(.A(G226), .B(G1698), .C1(new_n306), .C2(new_n307), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT74), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT74), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n251), .A2(new_n346), .A3(G226), .A4(G1698), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n251), .A2(G223), .A3(new_n252), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G33), .A2(G87), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n343), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(G1698), .B1(new_n249), .B2(new_n250), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(G223), .B1(G33), .B2(G87), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n354), .A2(KEYINPUT75), .A3(new_n345), .A4(new_n347), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n352), .A2(new_n256), .A3(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n265), .A2(new_n216), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(new_n261), .ZN(new_n358));
  AND3_X1   g0158(.A1(new_n356), .A2(new_n268), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(G200), .B1(new_n356), .B2(new_n358), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT77), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n356), .A2(new_n361), .A3(new_n268), .A4(new_n358), .ZN(new_n363));
  INV_X1    g0163(.A(new_n272), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n249), .A2(new_n224), .A3(new_n250), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT7), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n249), .A2(KEYINPUT7), .A3(new_n224), .A4(new_n250), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n209), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n215), .A2(new_n209), .ZN(new_n370));
  NOR2_X1   g0170(.A1(G58), .A2(G68), .ZN(new_n371));
  OAI21_X1  g0171(.A(G20), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n281), .A2(G159), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n364), .B1(new_n375), .B2(KEYINPUT16), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n367), .A2(KEYINPUT73), .A3(new_n368), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT73), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n365), .A2(new_n378), .A3(new_n366), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(G68), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n374), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n376), .B1(new_n382), .B2(KEYINPUT16), .ZN(new_n383));
  MUX2_X1   g0183(.A(new_n293), .B(new_n289), .S(new_n277), .Z(new_n384));
  NAND3_X1  g0184(.A1(new_n363), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n342), .B1(new_n362), .B2(new_n385), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n363), .A2(new_n383), .A3(new_n384), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n356), .A2(new_n358), .ZN(new_n388));
  INV_X1    g0188(.A(G200), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n356), .A2(new_n268), .A3(new_n358), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(KEYINPUT77), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n387), .A2(new_n392), .A3(KEYINPUT17), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n386), .A2(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n383), .A2(new_n384), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G179), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n356), .A2(new_n397), .A3(new_n358), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(G169), .B1(new_n356), .B2(new_n358), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n399), .A2(new_n400), .A3(KEYINPUT76), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT76), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n388), .A2(new_n301), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n402), .B1(new_n403), .B2(new_n398), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n396), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT18), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT76), .B1(new_n399), .B2(new_n400), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n403), .A2(new_n402), .A3(new_n398), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n395), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT18), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n394), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G238), .A2(G1698), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n251), .B(new_n413), .C1(new_n216), .C2(G1698), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n414), .B(new_n256), .C1(G107), .C2(new_n251), .ZN(new_n415));
  INV_X1    g0215(.A(G244), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n415), .B(new_n262), .C1(new_n416), .C2(new_n265), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G200), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n268), .B2(new_n417), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT8), .B(G58), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n421), .A2(new_n281), .B1(G20), .B2(G77), .ZN(new_n422));
  XOR2_X1   g0222(.A(KEYINPUT15), .B(G87), .Z(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n422), .B1(new_n278), .B2(new_n424), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n425), .A2(new_n272), .B1(G77), .B2(new_n292), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(G77), .B2(new_n289), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n419), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n417), .A2(new_n301), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n427), .B(new_n429), .C1(G179), .C2(new_n417), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n412), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n341), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n218), .B1(new_n249), .B2(new_n250), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT4), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n436), .A2(KEYINPUT79), .ZN(new_n437));
  OAI21_X1  g0237(.A(G1698), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G33), .A2(G283), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(G244), .B1(new_n306), .B2(new_n307), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n440), .B1(new_n441), .B2(new_n437), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(G244), .B(new_n252), .C1(new_n306), .C2(new_n307), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n436), .B1(new_n444), .B2(KEYINPUT79), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT80), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(KEYINPUT79), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT4), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT80), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n448), .A2(new_n449), .A3(new_n438), .A4(new_n442), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n446), .A2(new_n256), .A3(new_n450), .ZN(new_n451));
  XNOR2_X1  g0251(.A(KEYINPUT5), .B(G41), .ZN(new_n452));
  INV_X1    g0252(.A(G45), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(G1), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G274), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n455), .A2(new_n256), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n457), .B1(G257), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n451), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G200), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n377), .A2(G107), .A3(new_n379), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n282), .A2(new_n323), .ZN(new_n463));
  INV_X1    g0263(.A(G107), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(KEYINPUT6), .A3(G97), .ZN(new_n465));
  INV_X1    g0265(.A(G97), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(new_n464), .ZN(new_n467));
  NOR2_X1   g0267(.A1(G97), .A2(G107), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n465), .B1(new_n469), .B2(KEYINPUT6), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n463), .B1(new_n470), .B2(G20), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n462), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n272), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n289), .B1(G1), .B2(new_n248), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n272), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G97), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n290), .A2(new_n466), .ZN(new_n477));
  XNOR2_X1  g0277(.A(new_n477), .B(KEYINPUT78), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n473), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n451), .A2(G190), .A3(new_n459), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n461), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT81), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n461), .A2(new_n479), .A3(KEYINPUT81), .A4(new_n480), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n451), .A2(new_n397), .A3(new_n459), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n485), .B(KEYINPUT82), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n479), .B1(new_n301), .B2(new_n460), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n483), .A2(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT86), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n353), .A2(G257), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT85), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n251), .A2(G264), .A3(G1698), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n308), .A2(G303), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT85), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n353), .A2(new_n494), .A3(G257), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n491), .A2(new_n492), .A3(new_n493), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n256), .ZN(new_n497));
  NOR3_X1   g0297(.A1(new_n455), .A2(new_n236), .A3(new_n256), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n497), .A2(G179), .A3(new_n456), .A4(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n289), .A2(G116), .ZN(new_n501));
  INV_X1    g0301(.A(G116), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n272), .A2(new_n474), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(G20), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n439), .B(new_n224), .C1(G33), .C2(new_n466), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n272), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT20), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n272), .A2(KEYINPUT20), .A3(new_n504), .A4(new_n505), .ZN(new_n509));
  AOI211_X1 g0309(.A(new_n501), .B(new_n503), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n489), .B1(new_n500), .B2(new_n510), .ZN(new_n511));
  AOI211_X1 g0311(.A(new_n498), .B(new_n457), .C1(new_n496), .C2(new_n256), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n503), .B1(new_n508), .B2(new_n509), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(G116), .B2(new_n289), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n512), .A2(new_n514), .A3(KEYINPUT86), .A4(G179), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT21), .ZN(new_n517));
  INV_X1    g0317(.A(new_n512), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n510), .A2(new_n301), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR4_X1   g0320(.A1(new_n512), .A2(new_n510), .A3(KEYINPUT21), .A4(new_n301), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n516), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n251), .A2(G257), .A3(G1698), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n251), .A2(G250), .A3(new_n252), .ZN(new_n524));
  INV_X1    g0324(.A(G294), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n523), .B(new_n524), .C1(new_n248), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n256), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n458), .A2(G264), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(new_n456), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n301), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(G179), .B2(new_n529), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT24), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT87), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n224), .B(G87), .C1(new_n306), .C2(new_n307), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT22), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT22), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n251), .A2(new_n536), .A3(new_n224), .A4(G87), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n224), .A2(G107), .ZN(new_n539));
  XNOR2_X1  g0339(.A(new_n539), .B(KEYINPUT23), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n248), .A2(new_n502), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n224), .ZN(new_n542));
  AND4_X1   g0342(.A1(new_n533), .A2(new_n538), .A3(new_n540), .A4(new_n542), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n535), .A2(new_n537), .B1(new_n224), .B2(new_n541), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n533), .B1(new_n544), .B2(new_n540), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n532), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n538), .A2(new_n540), .A3(new_n542), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT87), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n544), .A2(new_n533), .A3(new_n540), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(KEYINPUT24), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n546), .A2(new_n272), .A3(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT25), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n289), .B2(G107), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n290), .A2(KEYINPUT25), .A3(new_n464), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n475), .A2(G107), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n531), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n522), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n514), .B1(new_n512), .B2(G190), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n389), .B2(new_n512), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n529), .A2(new_n389), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n527), .A2(new_n528), .A3(new_n268), .A4(new_n456), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(KEYINPUT88), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT88), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n529), .A2(new_n563), .A3(new_n389), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n551), .A2(new_n562), .A3(new_n555), .A4(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n218), .B1(new_n453), .B2(G1), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n454), .A2(new_n260), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n264), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n416), .A2(G1698), .ZN(new_n569));
  OAI221_X1 g0369(.A(new_n569), .B1(G238), .B2(G1698), .C1(new_n306), .C2(new_n307), .ZN(new_n570));
  INV_X1    g0370(.A(new_n541), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(G190), .B(new_n568), .C1(new_n572), .C2(new_n264), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n264), .B1(new_n570), .B2(new_n571), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n264), .A2(new_n566), .A3(new_n567), .ZN(new_n575));
  OAI21_X1  g0375(.A(G200), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n424), .A2(new_n290), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT84), .ZN(new_n579));
  AND2_X1   g0379(.A1(KEYINPUT83), .A2(G87), .ZN(new_n580));
  NOR2_X1   g0380(.A1(KEYINPUT83), .A2(G87), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n468), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n224), .B1(new_n248), .B2(new_n466), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n582), .A2(KEYINPUT19), .A3(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n224), .B(G68), .C1(new_n306), .C2(new_n307), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT19), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n278), .B2(new_n466), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n579), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n582), .A2(KEYINPUT19), .A3(new_n583), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n590), .A2(KEYINPUT84), .A3(new_n585), .A4(new_n587), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n591), .A3(new_n272), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n475), .A2(G87), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n577), .A2(new_n578), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n475), .A2(new_n423), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n592), .A2(new_n595), .A3(new_n578), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n574), .A2(new_n575), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n397), .ZN(new_n598));
  INV_X1    g0398(.A(new_n597), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n301), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n596), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n594), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n565), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n488), .A2(new_n557), .A3(new_n559), .A4(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n434), .A2(new_n604), .ZN(G372));
  NOR2_X1   g0405(.A1(new_n410), .A2(KEYINPUT18), .ZN(new_n606));
  AOI211_X1 g0406(.A(new_n406), .B(new_n395), .C1(new_n408), .C2(new_n409), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g0408(.A(new_n430), .B(KEYINPUT91), .Z(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n335), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n332), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n362), .A2(new_n342), .A3(new_n385), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT17), .B1(new_n387), .B2(new_n392), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n608), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n300), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n305), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n486), .A2(new_n487), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n619), .A2(KEYINPUT26), .A3(new_n602), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT26), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n486), .A2(new_n487), .ZN(new_n622));
  INV_X1    g0422(.A(new_n602), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n601), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT90), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n483), .A2(new_n484), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n629), .A2(new_n603), .A3(new_n622), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT89), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n522), .A2(new_n556), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT89), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n488), .A2(new_n633), .A3(new_n603), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n628), .A2(new_n631), .A3(new_n632), .A4(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n557), .B1(new_n630), .B2(KEYINPUT89), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n628), .B1(new_n636), .B2(new_n634), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n627), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n618), .B1(new_n639), .B2(new_n434), .ZN(G369));
  INV_X1    g0440(.A(G13), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n641), .A2(G20), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n258), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(G213), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(G343), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n514), .A2(new_n648), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n522), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n522), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(new_n559), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G330), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n648), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n522), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n556), .ZN(new_n658));
  INV_X1    g0458(.A(new_n565), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n655), .B1(new_n551), .B2(new_n555), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n556), .A2(new_n655), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n657), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n662), .ZN(G399));
  OR2_X1    g0466(.A1(new_n582), .A2(G116), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n204), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(G41), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n668), .A2(G1), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n227), .B2(new_n671), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT28), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT29), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n638), .A2(new_n675), .A3(new_n655), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT94), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n620), .A2(new_n677), .A3(new_n624), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n619), .A2(KEYINPUT94), .A3(KEYINPUT26), .A4(new_n602), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n632), .A2(new_n488), .A3(new_n603), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n678), .A2(new_n601), .A3(new_n679), .A4(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n655), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT29), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n676), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT30), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n512), .A2(G179), .A3(new_n459), .A4(new_n451), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n597), .A2(new_n527), .A3(new_n528), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT92), .ZN(new_n689));
  AOI21_X1  g0489(.A(G179), .B1(new_n451), .B2(new_n459), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n690), .A2(new_n518), .A3(new_n529), .A4(new_n599), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n460), .A2(new_n500), .ZN(new_n693));
  INV_X1    g0493(.A(new_n687), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(KEYINPUT30), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n689), .B1(new_n688), .B2(new_n691), .ZN(new_n697));
  OAI211_X1 g0497(.A(KEYINPUT31), .B(new_n648), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT31), .B1(new_n604), .B2(new_n648), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n688), .A2(new_n695), .A3(new_n691), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT93), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n688), .A2(new_n695), .A3(KEYINPUT93), .A4(new_n691), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(new_n648), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n699), .B1(new_n700), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n653), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n684), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n674), .B1(new_n708), .B2(G1), .ZN(G364));
  NAND2_X1  g0509(.A1(new_n642), .A2(G45), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n671), .A2(G1), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n652), .A2(new_n653), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n654), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(G13), .A2(G33), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G20), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n652), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n228), .A2(new_n453), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n669), .A2(new_n251), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n718), .B(new_n719), .C1(new_n242), .C2(new_n453), .ZN(new_n720));
  INV_X1    g0520(.A(G355), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n251), .A2(new_n204), .ZN(new_n722));
  OAI221_X1 g0522(.A(new_n720), .B1(G116), .B2(new_n204), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT95), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n223), .B1(G20), .B2(new_n301), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n716), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT96), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n711), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n224), .A2(new_n397), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(G190), .A3(G200), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G326), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G179), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G190), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G20), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n251), .B1(new_n736), .B2(G294), .ZN(new_n737));
  INV_X1    g0537(.A(G283), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n389), .A2(G179), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n224), .A2(G190), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n733), .B(new_n737), .C1(new_n738), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n730), .A2(G200), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G190), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  XOR2_X1   g0545(.A(KEYINPUT33), .B(G317), .Z(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n397), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n740), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G311), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n224), .A2(new_n268), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n752), .A2(new_n748), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G322), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR4_X1   g0556(.A1(new_n742), .A2(new_n747), .A3(new_n751), .A4(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G303), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n752), .A2(new_n739), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n759), .A2(KEYINPUT98), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(KEYINPUT98), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n757), .B1(new_n758), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n740), .A2(new_n734), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n763), .B1(G329), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT99), .ZN(new_n767));
  INV_X1    g0567(.A(new_n762), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n580), .A2(new_n581), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n308), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n770), .B1(new_n288), .B2(new_n731), .C1(new_n215), .C2(new_n754), .ZN(new_n771));
  INV_X1    g0571(.A(new_n749), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n772), .A2(G77), .B1(new_n736), .B2(G97), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n773), .B1(new_n464), .B2(new_n741), .C1(new_n745), .C2(new_n209), .ZN(new_n774));
  INV_X1    g0574(.A(G159), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n764), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT97), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT32), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n771), .A2(new_n774), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n725), .B1(new_n767), .B2(new_n779), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n717), .A2(new_n728), .A3(new_n729), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n713), .A2(new_n781), .ZN(G396));
  NAND3_X1  g0582(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(KEYINPUT90), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n636), .A2(new_n628), .A3(new_n634), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n648), .B1(new_n786), .B2(new_n627), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n427), .A2(new_n648), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n609), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n431), .A2(new_n789), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n788), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n638), .A2(new_n655), .A3(new_n793), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n795), .A2(new_n707), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n711), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT101), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n795), .A2(new_n796), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(new_n653), .B2(new_n706), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n797), .A2(KEYINPUT101), .A3(new_n711), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n800), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n793), .A2(new_n715), .ZN(new_n805));
  INV_X1    g0605(.A(new_n725), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n765), .A2(G132), .ZN(new_n807));
  INV_X1    g0607(.A(new_n736), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n744), .A2(G150), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n732), .A2(G137), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n772), .A2(G159), .ZN(new_n811));
  XOR2_X1   g0611(.A(KEYINPUT100), .B(G143), .Z(new_n812));
  NAND2_X1  g0612(.A1(new_n753), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n809), .A2(new_n810), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n807), .B1(new_n215), .B2(new_n808), .C1(new_n815), .C2(KEYINPUT34), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n308), .B(new_n816), .C1(KEYINPUT34), .C2(new_n815), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n817), .B1(new_n288), .B2(new_n762), .C1(new_n209), .C2(new_n741), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n762), .A2(new_n464), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n308), .B1(new_n731), .B2(new_n758), .C1(new_n808), .C2(new_n466), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n745), .A2(new_n738), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n754), .A2(new_n525), .B1(new_n764), .B2(new_n750), .ZN(new_n822));
  NOR4_X1   g0622(.A1(new_n819), .A2(new_n820), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n823), .B1(new_n217), .B2(new_n741), .C1(new_n502), .C2(new_n749), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n806), .B1(new_n818), .B2(new_n824), .ZN(new_n825));
  NOR3_X1   g0625(.A1(new_n725), .A2(G77), .A3(new_n714), .ZN(new_n826));
  NOR4_X1   g0626(.A1(new_n805), .A2(new_n711), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n804), .A2(new_n828), .ZN(G384));
  OAI21_X1  g0629(.A(new_n614), .B1(new_n606), .B2(new_n607), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n395), .A2(new_n646), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n387), .A2(new_n392), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n405), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(KEYINPUT37), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT37), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n405), .A2(new_n832), .A3(new_n836), .A4(new_n833), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n830), .A2(new_n831), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(KEYINPUT103), .B1(new_n838), .B2(KEYINPUT38), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n410), .A2(new_n831), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n836), .B1(new_n840), .B2(new_n833), .ZN(new_n841));
  INV_X1    g0641(.A(new_n837), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n412), .A2(new_n832), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT103), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT38), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n367), .A2(new_n368), .ZN(new_n847));
  OAI211_X1 g0647(.A(KEYINPUT16), .B(new_n381), .C1(new_n847), .C2(new_n209), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT16), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n369), .B2(new_n374), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n848), .A2(new_n272), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n384), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT102), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT102), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n384), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n408), .B2(new_n409), .ZN(new_n857));
  INV_X1    g0657(.A(new_n646), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n853), .A2(new_n858), .A3(new_n855), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n362), .B2(new_n385), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT37), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n837), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n862), .B(KEYINPUT38), .C1(new_n412), .C2(new_n859), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n839), .A2(new_n846), .A3(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT31), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n705), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n700), .B2(new_n705), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n331), .A2(new_n648), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n337), .B2(new_n333), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n332), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n868), .B1(new_n340), .B2(new_n332), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n793), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n864), .A2(KEYINPUT40), .A3(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT40), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n340), .A2(new_n332), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n869), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n794), .B1(new_n879), .B2(new_n871), .ZN(new_n880));
  INV_X1    g0680(.A(new_n705), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n629), .A2(new_n603), .A3(new_n622), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n882), .A2(new_n559), .A3(new_n557), .A4(new_n655), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n881), .B1(new_n883), .B2(KEYINPUT31), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n880), .B1(new_n884), .B2(new_n866), .ZN(new_n885));
  INV_X1    g0685(.A(new_n863), .ZN(new_n886));
  INV_X1    g0686(.A(new_n859), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n830), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT38), .B1(new_n888), .B2(new_n862), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n877), .B1(new_n885), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n876), .A2(new_n891), .A3(G330), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n700), .A2(new_n705), .ZN(new_n893));
  INV_X1    g0693(.A(new_n866), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n653), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n433), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n897), .B(KEYINPUT104), .Z(new_n898));
  INV_X1    g0698(.A(new_n867), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n876), .A2(new_n891), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n898), .B1(new_n434), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT39), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n886), .A2(new_n889), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n864), .B2(new_n902), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n332), .A2(new_n648), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n904), .A2(new_n905), .B1(new_n608), .B2(new_n646), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n430), .A2(new_n648), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n796), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n872), .A2(new_n873), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n909), .B(new_n911), .C1(new_n889), .C2(new_n886), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n906), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n617), .B1(new_n684), .B2(new_n433), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n913), .B(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n901), .B(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n258), .B2(new_n642), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n502), .B1(new_n470), .B2(KEYINPUT35), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n918), .B(new_n226), .C1(KEYINPUT35), .C2(new_n470), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT36), .ZN(new_n920));
  OAI21_X1  g0720(.A(G77), .B1(new_n215), .B2(new_n209), .ZN(new_n921));
  OAI22_X1  g0721(.A1(new_n921), .A2(new_n227), .B1(G50), .B2(new_n209), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(G1), .A3(new_n641), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n917), .A2(new_n920), .A3(new_n923), .ZN(G367));
  NOR2_X1   g0724(.A1(new_n741), .A2(new_n323), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n768), .A2(G58), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n772), .A2(G50), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n736), .A2(G68), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n732), .A2(new_n812), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n926), .A2(new_n927), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  AOI211_X1 g0730(.A(new_n925), .B(new_n930), .C1(G137), .C2(new_n765), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n308), .B1(new_n753), .B2(G150), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n931), .B(new_n932), .C1(new_n775), .C2(new_n745), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT106), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n741), .A2(new_n466), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n745), .A2(new_n525), .B1(new_n731), .B2(new_n750), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n754), .A2(new_n758), .B1(new_n749), .B2(new_n738), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n768), .A2(KEYINPUT46), .A3(G116), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT46), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n762), .B2(new_n502), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  AOI211_X1 g0742(.A(new_n935), .B(new_n942), .C1(G317), .C2(new_n765), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n943), .B(new_n308), .C1(new_n464), .C2(new_n808), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n934), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT47), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n725), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n592), .A2(new_n578), .A3(new_n593), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n648), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n602), .A2(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n601), .A2(new_n949), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n950), .A2(new_n716), .A3(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n719), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n726), .B1(new_n204), .B2(new_n424), .C1(new_n237), .C2(new_n953), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n947), .A2(new_n729), .A3(new_n952), .A4(new_n954), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT107), .Z(new_n956));
  NAND2_X1  g0756(.A1(new_n710), .A2(G1), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n708), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n662), .B1(new_n663), .B2(new_n656), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n488), .B1(new_n479), .B2(new_n655), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n619), .A2(new_n648), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OR3_X1    g0764(.A1(new_n961), .A2(KEYINPUT44), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(KEYINPUT44), .B1(new_n961), .B2(new_n964), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n654), .A2(new_n663), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT45), .ZN(new_n971));
  INV_X1    g0771(.A(new_n964), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n971), .B1(new_n972), .B2(new_n960), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n961), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AND3_X1   g0775(.A1(new_n968), .A2(new_n970), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n970), .B1(new_n968), .B2(new_n975), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n657), .B(new_n664), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n959), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n670), .B(KEYINPUT41), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n958), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n656), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n664), .A2(new_n632), .A3(new_n488), .A4(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT42), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n962), .A2(new_n658), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n648), .B1(new_n988), .B2(new_n622), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n950), .A2(new_n951), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n990), .B1(KEYINPUT43), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n969), .A2(new_n964), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT105), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n993), .B(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n992), .B(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n956), .B1(new_n984), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(G387));
  NAND2_X1  g0799(.A1(new_n959), .A2(new_n979), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n708), .A2(new_n980), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1000), .A2(new_n1001), .A3(new_n670), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n744), .A2(G311), .B1(G317), .B2(new_n753), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n758), .B2(new_n749), .C1(new_n755), .C2(new_n731), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT48), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n738), .B2(new_n808), .C1(new_n525), .C2(new_n762), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT49), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n251), .B1(new_n765), .B2(G326), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1007), .B(new_n1008), .C1(new_n502), .C2(new_n741), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n736), .A2(new_n423), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n775), .B2(new_n731), .C1(new_n762), .C2(new_n323), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n935), .B(new_n1011), .C1(G150), .C2(new_n765), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n753), .A2(G50), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n745), .A2(new_n277), .B1(new_n749), .B2(new_n209), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT110), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1012), .A2(new_n251), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n806), .B1(new_n1009), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n233), .A2(G45), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT108), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n420), .A2(G50), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1022), .A2(new_n668), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1019), .A2(new_n719), .A3(new_n1024), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(G107), .B2(new_n204), .C1(new_n668), .C2(new_n722), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1017), .B1(new_n727), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n663), .A2(new_n716), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1027), .A2(new_n729), .A3(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT111), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1002), .B(new_n1030), .C1(new_n958), .C2(new_n979), .ZN(G393));
  INV_X1    g0831(.A(new_n978), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n1001), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(KEYINPUT114), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n978), .A2(new_n708), .A3(new_n980), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT114), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1032), .A2(new_n1036), .A3(new_n1001), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1034), .A2(new_n670), .A3(new_n1035), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n978), .A2(new_n957), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n251), .B1(new_n772), .B2(G294), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n464), .B2(new_n741), .C1(new_n745), .C2(new_n758), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n732), .A2(G317), .B1(new_n753), .B2(G311), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT112), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT52), .Z(new_n1044));
  AOI211_X1 g0844(.A(new_n1041), .B(new_n1044), .C1(G322), .C2(new_n765), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n502), .B2(new_n808), .C1(new_n738), .C2(new_n762), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT113), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n808), .A2(new_n323), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n812), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n251), .B1(new_n1049), .B2(new_n764), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1048), .B(new_n1050), .C1(new_n421), .C2(new_n772), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n754), .A2(new_n775), .B1(new_n731), .B2(new_n280), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT51), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n768), .A2(G68), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n741), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n744), .A2(G50), .B1(new_n1055), .B2(G87), .ZN(new_n1056));
  AND4_X1   g0856(.A1(new_n1051), .A2(new_n1053), .A3(new_n1054), .A4(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n725), .B1(new_n1047), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n245), .A2(new_n719), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1059), .B(new_n726), .C1(new_n466), .C2(new_n204), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1058), .A2(new_n729), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n716), .B2(new_n972), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1038), .A2(new_n1039), .A3(new_n1063), .ZN(G390));
  INV_X1    g0864(.A(KEYINPUT118), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n681), .A2(new_n655), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n907), .B1(new_n1066), .B2(new_n793), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n893), .A2(new_n698), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1068), .A2(G330), .A3(new_n793), .A4(new_n911), .ZN(new_n1069));
  NOR3_X1   g0869(.A1(new_n867), .A2(new_n653), .A3(new_n794), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1067), .B(new_n1069), .C1(new_n911), .C2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1068), .A2(G330), .A3(new_n793), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n1072), .A2(new_n910), .B1(new_n880), .B2(new_n895), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n907), .B1(new_n787), .B2(new_n793), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1071), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1075), .A2(new_n896), .A3(new_n914), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n864), .A2(new_n902), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n903), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n910), .B1(new_n796), .B2(new_n908), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1079), .B1(new_n1080), .B2(new_n905), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n908), .B1(new_n682), .B2(new_n794), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n911), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n905), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1083), .A2(new_n864), .A3(new_n1084), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n1081), .A2(new_n1085), .A3(new_n1069), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n895), .A2(new_n880), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n1081), .B2(new_n1085), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1076), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n911), .B1(new_n895), .B2(new_n793), .ZN(new_n1090));
  NOR4_X1   g0890(.A1(new_n706), .A2(new_n910), .A3(new_n653), .A4(new_n794), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n706), .A2(new_n653), .A3(new_n794), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1087), .B1(new_n1093), .B2(new_n911), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1092), .A2(new_n1067), .B1(new_n1094), .B2(new_n909), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n683), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n787), .B2(new_n675), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n618), .B(new_n896), .C1(new_n1097), .C2(new_n434), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1081), .A2(new_n1085), .A3(new_n1069), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1085), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1084), .B1(new_n1074), .B2(new_n910), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1101), .B1(new_n1102), .B2(new_n1079), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1099), .B(new_n1100), .C1(new_n1103), .C2(new_n1087), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n1089), .A2(new_n1104), .A3(new_n670), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n957), .B(new_n1100), .C1(new_n1103), .C2(new_n1087), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1079), .A2(new_n714), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n725), .A2(new_n714), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n277), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n741), .A2(new_n209), .B1(new_n764), .B2(new_n525), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT117), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n731), .A2(new_n738), .B1(new_n749), .B2(new_n466), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G107), .B2(new_n744), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT116), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n308), .B1(new_n754), .B2(new_n502), .ZN(new_n1115));
  OR3_X1    g0915(.A1(new_n1114), .A2(new_n1048), .A3(new_n1115), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1111), .B(new_n1116), .C1(G87), .C2(new_n768), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n762), .A2(new_n280), .ZN(new_n1118));
  XOR2_X1   g0918(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n288), .B2(new_n741), .ZN(new_n1121));
  INV_X1    g0921(.A(G128), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n808), .A2(new_n775), .B1(new_n731), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(G137), .B2(new_n744), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n308), .B1(new_n753), .B2(G132), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1124), .B(new_n1125), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1126));
  XOR2_X1   g0926(.A(KEYINPUT54), .B(G143), .Z(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1128), .A2(new_n749), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n765), .A2(G125), .ZN(new_n1130));
  NOR4_X1   g0930(.A1(new_n1121), .A2(new_n1126), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n725), .B1(new_n1117), .B2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1107), .A2(new_n729), .A3(new_n1109), .A4(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1106), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1065), .B1(new_n1105), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1089), .A2(new_n1104), .A3(new_n670), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1136), .A2(KEYINPUT118), .A3(new_n1106), .A4(new_n1133), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1135), .A2(new_n1137), .ZN(G378));
  INV_X1    g0938(.A(KEYINPUT120), .ZN(new_n1139));
  XOR2_X1   g0939(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n300), .A2(new_n305), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1141), .B1(new_n300), .B2(new_n305), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n294), .A2(new_n858), .ZN(new_n1144));
  OR3_X1    g0944(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1144), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n892), .A2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1147), .A2(new_n876), .A3(new_n891), .A4(G330), .ZN(new_n1150));
  AND4_X1   g0950(.A1(new_n912), .A2(new_n1149), .A3(new_n906), .A4(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1149), .A2(new_n1150), .B1(new_n906), .B2(new_n912), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1139), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n913), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1149), .A2(new_n906), .A3(new_n912), .A4(new_n1150), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(KEYINPUT120), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1098), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1153), .A2(new_n1157), .B1(new_n1104), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(KEYINPUT121), .B1(new_n1159), .B2(KEYINPUT57), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1155), .A2(KEYINPUT120), .A3(new_n1156), .ZN(new_n1161));
  AOI21_X1  g0961(.A(KEYINPUT120), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(new_n1086), .A2(new_n1088), .A3(new_n1076), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n1161), .A2(new_n1162), .B1(new_n1163), .B2(new_n1098), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT121), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT57), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n1104), .B2(new_n1158), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n671), .B1(new_n1169), .B2(KEYINPUT57), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1160), .A2(new_n1167), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n711), .B1(new_n288), .B2(new_n1108), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n1148), .B2(new_n715), .ZN(new_n1173));
  INV_X1    g0973(.A(G41), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1174), .B1(new_n502), .B2(new_n731), .C1(new_n745), .C2(new_n466), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n928), .B1(new_n762), .B2(new_n323), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n741), .A2(new_n215), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n308), .B1(new_n764), .B2(new_n738), .ZN(new_n1178));
  NOR4_X1   g0978(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n464), .B2(new_n754), .C1(new_n424), .C2(new_n749), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT58), .ZN(new_n1181));
  AOI21_X1  g0981(.A(G50), .B1(new_n250), .B2(new_n1174), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT119), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n768), .A2(new_n1127), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n753), .A2(G128), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n772), .A2(G137), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n744), .A2(G132), .B1(G150), .B2(new_n736), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G125), .B2(new_n732), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT59), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(G33), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1192));
  AOI21_X1  g0992(.A(G41), .B1(new_n765), .B2(G124), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(new_n775), .C2(new_n741), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1181), .B(new_n1183), .C1(new_n1191), .C2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1173), .B1(new_n725), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1153), .A2(new_n1157), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1196), .B1(new_n1197), .B2(new_n957), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1171), .A2(new_n1198), .ZN(G375));
  NAND2_X1  g0999(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1200), .A2(new_n1076), .A3(new_n982), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n745), .A2(new_n502), .B1(new_n464), .B2(new_n749), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1202), .A2(KEYINPUT122), .B1(G283), .B2(new_n753), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1203), .B(new_n1010), .C1(KEYINPUT122), .C2(new_n1202), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n762), .A2(new_n466), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n308), .B1(new_n764), .B2(new_n758), .C1(new_n731), .C2(new_n525), .ZN(new_n1206));
  NOR4_X1   g1006(.A1(new_n1204), .A2(new_n925), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n732), .A2(G132), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT123), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n775), .B2(new_n762), .C1(new_n745), .C2(new_n1128), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n764), .A2(new_n1122), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n753), .A2(G137), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n308), .B1(new_n736), .B2(G50), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n215), .B2(new_n741), .C1(new_n280), .C2(new_n749), .ZN(new_n1214));
  NOR4_X1   g1014(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n725), .B1(new_n1207), .B2(new_n1215), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n729), .B(new_n1216), .C1(new_n911), .C2(new_n715), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n209), .B2(new_n1108), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1075), .B2(new_n957), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1201), .A2(new_n1219), .ZN(G381));
  NOR2_X1   g1020(.A1(new_n1105), .A2(new_n1134), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(G375), .A2(new_n1222), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n998), .A2(new_n1038), .A3(new_n1039), .A4(new_n1063), .ZN(new_n1224));
  OR3_X1    g1024(.A1(G393), .A2(G381), .A3(G396), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1224), .A2(G384), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1223), .A2(new_n1226), .ZN(G407));
  OAI21_X1  g1027(.A(new_n1223), .B1(new_n1226), .B2(new_n647), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(G213), .ZN(G409));
  INV_X1    g1029(.A(G213), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1230), .A2(G343), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1171), .A2(G378), .A3(new_n1198), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT124), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1168), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1155), .A2(KEYINPUT124), .A3(new_n1156), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(new_n957), .A3(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1164), .B2(new_n983), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1221), .B1(new_n1237), .B2(new_n1196), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1231), .B1(new_n1232), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT60), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n671), .B1(new_n1200), .B2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1095), .A2(new_n1098), .A3(KEYINPUT60), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1241), .A2(new_n1076), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1219), .ZN(new_n1244));
  INV_X1    g1044(.A(G384), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1243), .A2(G384), .A3(new_n1219), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1246), .A2(KEYINPUT125), .A3(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1231), .A2(G2897), .ZN(new_n1249));
  OR2_X1    g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT125), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1247), .ZN(new_n1252));
  AOI21_X1  g1052(.A(G384), .B1(new_n1243), .B2(new_n1219), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1251), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1254), .A2(new_n1249), .A3(new_n1248), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1250), .A2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(KEYINPUT63), .B1(new_n1239), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1239), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1257), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1239), .A2(KEYINPUT63), .A3(new_n1259), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT126), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(G390), .A2(G387), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1224), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(G393), .B(G396), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1264), .A2(new_n1224), .A3(new_n1266), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1270), .A2(KEYINPUT61), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n1231), .B(new_n1258), .C1(new_n1232), .C2(new_n1238), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT126), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(new_n1273), .A3(KEYINPUT63), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1261), .A2(new_n1263), .A3(new_n1271), .A4(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT62), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n1272), .A2(new_n1276), .B1(new_n1239), .B2(new_n1256), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1232), .A2(new_n1238), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1231), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1278), .A2(new_n1276), .A3(new_n1279), .A4(new_n1259), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT61), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1270), .B1(new_n1277), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1275), .A2(new_n1283), .ZN(G405));
  INV_X1    g1084(.A(new_n1232), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1222), .B1(new_n1171), .B2(new_n1198), .ZN(new_n1286));
  OR2_X1    g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1258), .A2(KEYINPUT127), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1268), .B(new_n1269), .C1(KEYINPUT127), .C2(new_n1258), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1258), .A2(KEYINPUT127), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1269), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1266), .B1(new_n1264), .B2(new_n1224), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1291), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1290), .A2(new_n1294), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1289), .B(new_n1295), .ZN(G402));
endmodule


