//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  AND2_X1   g001(.A1(new_n187), .A2(G952), .ZN(new_n188));
  NAND2_X1  g002(.A1(G234), .A2(G237), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(G902), .A3(G953), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT21), .B(G898), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n191), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(G214), .B1(G237), .B2(G902), .ZN(new_n197));
  OAI21_X1  g011(.A(G210), .B1(G237), .B2(G902), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT79), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(KEYINPUT3), .ZN(new_n200));
  INV_X1    g014(.A(G104), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G107), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(KEYINPUT3), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n200), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(G107), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT79), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G104), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n205), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(G101), .B1(new_n204), .B2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n208), .A2(G104), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n212), .B1(new_n200), .B2(new_n202), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n206), .A2(KEYINPUT79), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n207), .B1(new_n215), .B2(new_n209), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n213), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n211), .A2(KEYINPUT4), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n214), .B1(new_n213), .B2(new_n216), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT4), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT2), .ZN(new_n223));
  INV_X1    g037(.A(G113), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT69), .B1(KEYINPUT2), .B2(G113), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT2), .A2(G113), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(G116), .B(G119), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n227), .A2(new_n228), .A3(new_n230), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n218), .A2(new_n221), .A3(new_n234), .A4(KEYINPUT81), .ZN(new_n235));
  OAI21_X1  g049(.A(G101), .B1(new_n202), .B2(new_n212), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n217), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT5), .ZN(new_n238));
  INV_X1    g052(.A(G119), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(new_n239), .A3(G116), .ZN(new_n240));
  OAI211_X1 g054(.A(G113), .B(new_n240), .C1(new_n231), .C2(new_n238), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n237), .A2(new_n233), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n235), .A2(new_n242), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n220), .A2(new_n219), .B1(new_n232), .B2(new_n233), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT81), .B1(new_n244), .B2(new_n218), .ZN(new_n245));
  XNOR2_X1  g059(.A(G110), .B(G122), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NOR3_X1   g061(.A1(new_n243), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  XOR2_X1   g063(.A(new_n246), .B(KEYINPUT82), .Z(new_n250));
  AND2_X1   g064(.A1(new_n250), .A2(KEYINPUT83), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n251), .B1(new_n243), .B2(new_n245), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT6), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI211_X1 g068(.A(KEYINPUT6), .B(new_n251), .C1(new_n243), .C2(new_n245), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n249), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G128), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(KEYINPUT1), .ZN(new_n258));
  INV_X1    g072(.A(G146), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G143), .ZN(new_n260));
  INV_X1    g074(.A(G143), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G146), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n258), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n259), .A2(KEYINPUT64), .A3(G143), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT64), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n265), .B1(new_n261), .B2(G146), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n261), .A2(G146), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n264), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n269));
  OAI21_X1  g083(.A(G128), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n263), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G125), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT0), .B(G128), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT64), .B1(new_n259), .B2(G143), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n260), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n274), .B1(new_n276), .B2(new_n264), .ZN(new_n277));
  AND2_X1   g091(.A1(KEYINPUT0), .A2(G128), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n260), .A2(new_n262), .A3(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(G125), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(G224), .A3(new_n187), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n187), .A2(G224), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n273), .A2(new_n283), .A3(new_n280), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n256), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G902), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n246), .B(KEYINPUT8), .ZN(new_n288));
  AND4_X1   g102(.A1(new_n233), .A2(new_n241), .A3(new_n217), .A4(new_n236), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n241), .A2(new_n233), .B1(new_n217), .B2(new_n236), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n273), .A2(new_n280), .A3(KEYINPUT7), .A4(new_n283), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT7), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n281), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n291), .A2(new_n282), .A3(new_n292), .A4(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n287), .B1(new_n248), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n198), .B1(new_n286), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n198), .ZN(new_n299));
  AOI211_X1 g113(.A(new_n299), .B(new_n296), .C1(new_n256), .C2(new_n285), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n196), .B(new_n197), .C1(new_n298), .C2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G221), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT9), .B(G234), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n303), .B1(new_n305), .B2(new_n287), .ZN(new_n306));
  INV_X1    g120(.A(G469), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(new_n287), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT66), .B(G131), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT65), .ZN(new_n310));
  INV_X1    g124(.A(G134), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n310), .A2(KEYINPUT11), .B1(new_n311), .B2(G137), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT11), .ZN(new_n313));
  INV_X1    g127(.A(G137), .ZN(new_n314));
  AND4_X1   g128(.A1(KEYINPUT65), .A2(new_n313), .A3(new_n314), .A4(G134), .ZN(new_n315));
  AOI22_X1  g129(.A1(KEYINPUT65), .A2(new_n313), .B1(new_n314), .B2(G134), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n309), .B(new_n312), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G131), .ZN(new_n319));
  OAI22_X1  g133(.A1(new_n310), .A2(KEYINPUT11), .B1(new_n311), .B2(G137), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT65), .A4(G134), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n319), .B1(new_n322), .B2(new_n312), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n217), .A2(new_n236), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n271), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n258), .A2(new_n260), .A3(new_n262), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n260), .A2(new_n262), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n257), .B1(new_n260), .B2(KEYINPUT1), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n217), .A2(new_n330), .A3(new_n236), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n324), .B1(new_n326), .B2(new_n331), .ZN(new_n332));
  NOR3_X1   g146(.A1(new_n332), .A2(KEYINPUT80), .A3(KEYINPUT12), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n259), .A2(KEYINPUT64), .A3(G143), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n334), .B1(new_n260), .B2(new_n275), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n327), .B1(new_n335), .B2(new_n329), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n237), .A2(KEYINPUT10), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n274), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n279), .B1(new_n268), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n218), .A2(new_n339), .A3(new_n221), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT10), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n331), .A2(new_n341), .ZN(new_n342));
  AND4_X1   g156(.A1(new_n324), .A2(new_n337), .A3(new_n340), .A4(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n333), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(G110), .B(G140), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n187), .A2(G227), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT80), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n349), .B1(new_n332), .B2(KEYINPUT12), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n326), .A2(new_n331), .ZN(new_n351));
  OAI22_X1  g165(.A1(KEYINPUT65), .A2(new_n313), .B1(new_n314), .B2(G134), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(new_n320), .B2(new_n321), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n317), .B1(new_n353), .B2(new_n319), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT12), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n350), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n344), .A2(new_n348), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n337), .A2(new_n340), .A3(new_n342), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n354), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n337), .A2(new_n340), .A3(new_n324), .A4(new_n342), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n347), .ZN(new_n364));
  AOI21_X1  g178(.A(G902), .B1(new_n359), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n308), .B1(new_n365), .B2(new_n307), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n350), .A2(new_n357), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n355), .A2(new_n349), .A3(new_n356), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n362), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n347), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n363), .A2(new_n347), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(G469), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n306), .B1(new_n366), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G478), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(KEYINPUT15), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n257), .A2(G143), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n261), .A2(G128), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(new_n311), .ZN(new_n380));
  INV_X1    g194(.A(G122), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G116), .ZN(new_n382));
  INV_X1    g196(.A(G116), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G122), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT85), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(G116), .B(G122), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(KEYINPUT85), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n208), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n383), .A2(KEYINPUT14), .A3(G122), .ZN(new_n391));
  OAI211_X1 g205(.A(G107), .B(new_n391), .C1(new_n385), .C2(KEYINPUT14), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n380), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n379), .A2(new_n311), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n385), .A2(new_n386), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n388), .A2(KEYINPUT85), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n396), .A3(G107), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(G107), .B1(new_n395), .B2(new_n396), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n394), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT87), .ZN(new_n401));
  XOR2_X1   g215(.A(KEYINPUT86), .B(KEYINPUT13), .Z(new_n402));
  OAI21_X1  g216(.A(new_n401), .B1(new_n402), .B2(new_n377), .ZN(new_n403));
  XNOR2_X1  g217(.A(KEYINPUT86), .B(KEYINPUT13), .ZN(new_n404));
  INV_X1    g218(.A(new_n377), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n405), .A3(KEYINPUT87), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n378), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n408), .B1(new_n404), .B2(new_n405), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n311), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n393), .B1(new_n400), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G217), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n304), .A2(new_n413), .A3(G953), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n393), .B(new_n414), .C1(new_n400), .C2(new_n411), .ZN(new_n417));
  AOI21_X1  g231(.A(G902), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT88), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI211_X1 g234(.A(KEYINPUT88), .B(G902), .C1(new_n416), .C2(new_n417), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n376), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n417), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n390), .A2(new_n397), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n409), .B1(new_n403), .B2(new_n406), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n424), .B(new_n394), .C1(new_n311), .C2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n414), .B1(new_n426), .B2(new_n393), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n287), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n376), .B1(new_n428), .B2(KEYINPUT88), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n422), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G237), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(new_n187), .A3(G214), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n261), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n432), .A2(new_n187), .A3(G143), .A4(G214), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(KEYINPUT18), .A2(G131), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G140), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G125), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n272), .A2(G140), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G146), .ZN(new_n443));
  XNOR2_X1  g257(.A(G125), .B(G140), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n259), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n436), .A2(new_n438), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n446), .B1(new_n436), .B2(new_n438), .ZN(new_n447));
  INV_X1    g261(.A(new_n309), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n436), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n434), .A2(new_n309), .A3(new_n435), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n451), .A2(KEYINPUT17), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT16), .ZN(new_n453));
  OR3_X1    g267(.A1(new_n272), .A2(KEYINPUT16), .A3(G140), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n259), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n453), .A2(new_n454), .A3(G146), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT17), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n456), .B(new_n457), .C1(new_n449), .C2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n447), .B1(new_n452), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G113), .B(G122), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(new_n201), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n447), .B(new_n462), .C1(new_n452), .C2(new_n459), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n287), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G475), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n444), .A2(KEYINPUT19), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n444), .A2(KEYINPUT19), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n259), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n451), .A2(new_n457), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT84), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n447), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n463), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n473), .B1(new_n472), .B2(new_n447), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n465), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT20), .ZN(new_n478));
  NOR2_X1   g292(.A1(G475), .A2(G902), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n478), .B1(new_n477), .B2(new_n479), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n468), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n431), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n302), .A2(new_n374), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT68), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n314), .A2(G134), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n311), .A2(G137), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n319), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n317), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n486), .B1(new_n491), .B2(new_n271), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n489), .B1(new_n353), .B2(new_n309), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(new_n336), .A3(KEYINPUT68), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT67), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n354), .A2(new_n496), .A3(new_n339), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n339), .B1(new_n318), .B2(new_n323), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT67), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n495), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT71), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n501), .A3(new_n234), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n493), .A2(new_n336), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(new_n234), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n501), .B1(new_n500), .B2(new_n234), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT28), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n505), .A2(KEYINPUT28), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT26), .B(G101), .ZN(new_n513));
  INV_X1    g327(.A(G210), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n514), .A2(G237), .A3(G953), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n513), .B(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT30), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n500), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n504), .A2(new_n519), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n520), .A2(new_n234), .A3(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n518), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n506), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT31), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n521), .B1(new_n500), .B2(new_n519), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n505), .B1(new_n528), .B2(new_n234), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(KEYINPUT31), .A3(new_n524), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n512), .A2(new_n518), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(G472), .A2(G902), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT32), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n508), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(new_n506), .A3(new_n502), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n510), .B1(new_n536), .B2(KEYINPUT28), .ZN(new_n537));
  AND4_X1   g351(.A1(KEYINPUT31), .A2(new_n523), .A3(new_n506), .A4(new_n524), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT31), .B1(new_n529), .B2(new_n524), .ZN(new_n539));
  OAI22_X1  g353(.A1(new_n537), .A2(new_n524), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT32), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n541), .A3(new_n532), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT29), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n523), .A2(new_n506), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n518), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n543), .B(new_n545), .C1(new_n512), .C2(new_n518), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT72), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n504), .A2(new_n234), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n506), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n504), .A2(KEYINPUT72), .A3(new_n234), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(KEYINPUT28), .A3(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n551), .A2(KEYINPUT29), .A3(new_n511), .A4(new_n524), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n552), .A2(new_n287), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n546), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n534), .A2(new_n542), .B1(new_n554), .B2(G472), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n239), .A2(G128), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n257), .A2(G119), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT24), .B(G110), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT74), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT23), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT23), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT74), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n562), .A2(new_n557), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(KEYINPUT23), .A2(G119), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT73), .B1(new_n566), .B2(G128), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT73), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n568), .A2(new_n257), .A3(KEYINPUT23), .A4(G119), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n565), .A2(new_n567), .A3(new_n556), .A4(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n560), .B1(new_n570), .B2(G110), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(new_n457), .A3(new_n445), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT76), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n570), .A2(G110), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT75), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT75), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n570), .A2(new_n576), .A3(G110), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n558), .A2(new_n559), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n456), .B2(new_n457), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n573), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n570), .A2(new_n576), .A3(G110), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n576), .B1(new_n570), .B2(G110), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n580), .B(new_n573), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n572), .B1(new_n581), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT22), .B(G137), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n587), .B(new_n588), .Z(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n572), .B(new_n589), .C1(new_n581), .C2(new_n585), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n287), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT77), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT25), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n593), .A2(new_n594), .A3(KEYINPUT25), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n413), .B1(G234), .B2(new_n287), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n591), .A2(new_n592), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n599), .A2(G902), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT78), .B1(new_n555), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n554), .A2(G472), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n531), .A2(KEYINPUT32), .A3(new_n533), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n541), .B1(new_n540), .B2(new_n532), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT78), .ZN(new_n610));
  INV_X1    g424(.A(new_n604), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n485), .B1(new_n605), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(new_n214), .ZN(G3));
  OAI21_X1  g428(.A(G472), .B1(new_n531), .B2(G902), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n540), .A2(new_n532), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n611), .A2(new_n615), .A3(new_n616), .A4(new_n374), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT90), .ZN(new_n618));
  INV_X1    g432(.A(new_n482), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n619), .A2(new_n480), .B1(G475), .B2(new_n467), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT89), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(KEYINPUT89), .A2(KEYINPUT33), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n623), .B(new_n624), .C1(new_n423), .C2(new_n427), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n416), .A2(new_n621), .A3(new_n622), .A4(new_n417), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n375), .A2(G902), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n627), .A2(new_n628), .B1(new_n375), .B2(new_n428), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n620), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n618), .B1(new_n301), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n197), .ZN(new_n633));
  INV_X1    g447(.A(new_n285), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n248), .B1(new_n253), .B2(new_n252), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n634), .B1(new_n635), .B2(new_n255), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n299), .B1(new_n636), .B2(new_n296), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n286), .A2(new_n198), .A3(new_n297), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n633), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n639), .A2(KEYINPUT90), .A3(new_n196), .A4(new_n630), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n617), .B1(new_n632), .B2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT91), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT34), .B(G104), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  NAND2_X1  g458(.A1(new_n431), .A2(new_n620), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n617), .A2(new_n301), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT35), .B(G107), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  NOR2_X1   g462(.A1(new_n590), .A2(KEYINPUT36), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n586), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n602), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n600), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n615), .A2(new_n616), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n485), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n654), .B(KEYINPUT92), .Z(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT37), .B(G110), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  NAND2_X1  g471(.A1(new_n652), .A2(new_n374), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT93), .B(G900), .Z(new_n660));
  AOI21_X1  g474(.A(new_n191), .B1(new_n193), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n468), .B(new_n662), .C1(new_n481), .C2(new_n482), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(KEYINPUT94), .A3(new_n431), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT94), .ZN(new_n666));
  INV_X1    g480(.A(new_n376), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n428), .A2(KEYINPUT88), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n418), .A2(new_n419), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n429), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n666), .B1(new_n671), .B2(new_n663), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n665), .A2(new_n639), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n609), .A2(new_n659), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT95), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n534), .A2(new_n542), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n658), .B1(new_n678), .B2(new_n606), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(KEYINPUT95), .A3(new_n674), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G128), .ZN(G30));
  XOR2_X1   g496(.A(new_n661), .B(KEYINPUT39), .Z(new_n683));
  NAND2_X1  g497(.A1(new_n374), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT40), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n549), .A2(new_n550), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n287), .B1(new_n686), .B2(new_n524), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n529), .A2(new_n518), .ZN(new_n688));
  OAI21_X1  g502(.A(G472), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n678), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n637), .A2(new_n638), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n691), .B(KEYINPUT38), .Z(new_n692));
  INV_X1    g506(.A(new_n599), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n595), .B2(new_n596), .ZN(new_n694));
  AOI22_X1  g508(.A1(new_n694), .A2(new_n598), .B1(new_n602), .B2(new_n650), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n671), .A2(new_n620), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n695), .A2(new_n197), .A3(new_n696), .ZN(new_n697));
  NOR4_X1   g511(.A1(new_n685), .A2(new_n690), .A3(new_n692), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(new_n261), .ZN(G45));
  NAND2_X1  g513(.A1(new_n691), .A2(new_n197), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n630), .A2(new_n662), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n679), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT96), .B(G146), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G48));
  NAND2_X1  g519(.A1(new_n632), .A2(new_n640), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n365), .B(new_n307), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n306), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n706), .A2(new_n609), .A3(new_n611), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT41), .B(G113), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NOR2_X1   g525(.A1(new_n301), .A2(new_n645), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n609), .A2(new_n611), .A3(new_n712), .A4(new_n708), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G116), .ZN(G18));
  NOR3_X1   g528(.A1(new_n700), .A2(new_n306), .A3(new_n707), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n652), .A2(new_n196), .A3(new_n484), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n609), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G119), .ZN(G21));
  NAND2_X1  g532(.A1(new_n639), .A2(new_n696), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n527), .A2(new_n530), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n551), .A2(new_n511), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n518), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n533), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n538), .A2(new_n539), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n524), .B1(new_n509), .B2(new_n511), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n287), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n724), .B1(new_n727), .B2(G472), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n707), .A2(new_n306), .A3(new_n195), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n720), .A2(new_n728), .A3(new_n729), .A4(new_n611), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  INV_X1    g545(.A(new_n701), .ZN(new_n732));
  AOI21_X1  g546(.A(KEYINPUT97), .B1(new_n728), .B2(new_n652), .ZN(new_n733));
  INV_X1    g547(.A(G472), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n540), .B2(new_n287), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT97), .ZN(new_n736));
  NOR4_X1   g550(.A1(new_n735), .A2(new_n695), .A3(new_n736), .A4(new_n724), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n732), .B(new_n715), .C1(new_n733), .C2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  INV_X1    g553(.A(new_n306), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT99), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n344), .A2(new_n358), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT98), .B1(new_n742), .B2(new_n347), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n372), .A2(new_n370), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n743), .B1(new_n744), .B2(KEYINPUT98), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n741), .B1(new_n745), .B2(G469), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n348), .B1(new_n344), .B2(new_n358), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT98), .B1(new_n747), .B2(new_n371), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT98), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n370), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n748), .A2(new_n741), .A3(G469), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n366), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n740), .B1(new_n746), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT100), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT100), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n755), .B(new_n740), .C1(new_n746), .C2(new_n752), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n691), .A2(new_n633), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n754), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n555), .A2(new_n604), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT101), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT42), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n701), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n758), .A2(new_n759), .A3(new_n762), .A4(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n757), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n766), .B1(new_n753), .B2(KEYINPUT100), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n759), .A2(new_n767), .A3(new_n756), .A4(new_n762), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n763), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(KEYINPUT102), .B(G131), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n770), .B(new_n771), .ZN(G33));
  AND2_X1   g586(.A1(new_n665), .A2(new_n672), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n758), .A2(KEYINPUT103), .A3(new_n759), .A4(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n759), .A2(new_n767), .A3(new_n773), .A4(new_n756), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT103), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  XOR2_X1   g592(.A(KEYINPUT104), .B(G134), .Z(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(G36));
  NAND2_X1  g594(.A1(new_n745), .A2(KEYINPUT45), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n307), .B1(new_n744), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n308), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT46), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT105), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n365), .A2(new_n307), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n787), .B1(new_n784), .B2(KEYINPUT46), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n683), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n789), .A2(new_n306), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n615), .A2(new_n616), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n483), .A2(new_n629), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT43), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n794), .A3(new_n652), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT44), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n766), .B1(new_n795), .B2(new_n796), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n791), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G137), .ZN(G39));
  NAND4_X1  g614(.A1(new_n555), .A2(new_n604), .A3(new_n732), .A4(new_n757), .ZN(new_n801));
  XOR2_X1   g615(.A(new_n801), .B(KEYINPUT106), .Z(new_n802));
  INV_X1    g616(.A(KEYINPUT47), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(new_n789), .B2(new_n306), .ZN(new_n804));
  OAI211_X1 g618(.A(KEYINPUT47), .B(new_n740), .C1(new_n786), .C2(new_n788), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(new_n439), .ZN(G42));
  AOI21_X1  g621(.A(KEYINPUT95), .B1(new_n679), .B2(new_n674), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n555), .A2(new_n658), .A3(new_n673), .A4(new_n676), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n738), .B(new_n703), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n690), .A2(new_n719), .ZN(new_n811));
  INV_X1    g625(.A(new_n753), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n652), .A2(new_n661), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT110), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT52), .B1(new_n810), .B2(new_n815), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n677), .A2(new_n680), .B1(new_n679), .B2(new_n702), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n817), .A2(new_n818), .A3(new_n738), .A4(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n816), .A2(KEYINPUT53), .A3(new_n820), .ZN(new_n821));
  AND4_X1   g635(.A1(new_n709), .A2(new_n713), .A3(new_n717), .A4(new_n730), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n822), .A2(new_n769), .A3(new_n765), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT109), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n732), .B1(new_n733), .B2(new_n737), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n767), .A2(new_n756), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n724), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n615), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n736), .B1(new_n829), .B2(new_n695), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n728), .A2(KEYINPUT97), .A3(new_n652), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n701), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n758), .A3(KEYINPUT109), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n827), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(KEYINPUT107), .B1(new_n670), .B2(new_n429), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT107), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n422), .A2(new_n430), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n483), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n838), .A2(KEYINPUT108), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n631), .B1(new_n838), .B2(KEYINPUT108), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n302), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI22_X1  g655(.A1(new_n841), .A2(new_n617), .B1(new_n485), .B2(new_n653), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n757), .A2(new_n664), .A3(new_n835), .A4(new_n837), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n555), .A2(new_n843), .A3(new_n658), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n613), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n778), .A2(new_n834), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT112), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT112), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n834), .A2(new_n778), .A3(new_n845), .A4(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n821), .A2(new_n823), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n823), .A2(new_n816), .A3(new_n820), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n852), .B1(new_n853), .B2(new_n846), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n850), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n853), .A2(new_n852), .A3(new_n846), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT111), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n858), .A3(new_n854), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n823), .A2(new_n816), .A3(new_n820), .ZN(new_n860));
  INV_X1    g674(.A(new_n846), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT53), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n856), .B1(new_n862), .B2(KEYINPUT111), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n855), .B1(new_n864), .B2(new_n851), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n794), .A2(new_n191), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n866), .A2(new_n611), .A3(new_n728), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n692), .A2(new_n633), .A3(new_n708), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n867), .A2(KEYINPUT50), .A3(new_n868), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT117), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n867), .A2(new_n868), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n871), .A2(KEYINPUT114), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT116), .ZN(new_n873));
  XNOR2_X1  g687(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n874), .B1(new_n871), .B2(KEYINPUT114), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n873), .B1(new_n872), .B2(new_n875), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n870), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n604), .A2(new_n190), .ZN(new_n879));
  AND4_X1   g693(.A1(new_n690), .A2(new_n708), .A3(new_n757), .A4(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(new_n620), .A3(new_n629), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT118), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n830), .A2(new_n831), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n866), .A2(new_n708), .A3(new_n757), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n867), .A2(new_n757), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT113), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n804), .A2(new_n805), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n707), .A2(new_n740), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n878), .A2(new_n885), .A3(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT51), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n867), .A2(new_n715), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n188), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n884), .A2(new_n759), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT48), .Z(new_n898));
  AOI211_X1 g712(.A(new_n896), .B(new_n898), .C1(new_n630), .C2(new_n880), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n893), .A2(new_n894), .A3(new_n899), .ZN(new_n900));
  OAI22_X1  g714(.A1(new_n865), .A2(new_n900), .B1(G952), .B2(G953), .ZN(new_n901));
  AND4_X1   g715(.A1(new_n611), .A2(new_n740), .A3(new_n197), .A4(new_n793), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n707), .B(KEYINPUT49), .Z(new_n903));
  NAND4_X1  g717(.A1(new_n690), .A2(new_n902), .A3(new_n903), .A4(new_n692), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n901), .A2(new_n904), .ZN(G75));
  NOR2_X1   g719(.A1(new_n187), .A2(G952), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT119), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n850), .A2(new_n854), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(G902), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n909), .B1(new_n911), .B2(new_n514), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n256), .B(new_n285), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT55), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n912), .A2(new_n915), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n908), .B1(new_n916), .B2(new_n917), .ZN(G51));
  INV_X1    g732(.A(KEYINPUT120), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n781), .A2(new_n783), .ZN(new_n920));
  AOI211_X1 g734(.A(new_n287), .B(new_n920), .C1(new_n850), .C2(new_n854), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n308), .B(KEYINPUT57), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n850), .A2(new_n851), .A3(new_n854), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n851), .B1(new_n850), .B2(new_n854), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n359), .A2(new_n364), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n921), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n919), .B1(new_n927), .B2(new_n906), .ZN(new_n928));
  INV_X1    g742(.A(new_n906), .ZN(new_n929));
  INV_X1    g743(.A(new_n926), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n847), .A2(new_n849), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n823), .A2(new_n816), .A3(KEYINPUT53), .A4(new_n820), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT54), .B1(new_n933), .B2(new_n862), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n855), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n930), .B1(new_n935), .B2(new_n922), .ZN(new_n936));
  OAI211_X1 g750(.A(KEYINPUT120), .B(new_n929), .C1(new_n936), .C2(new_n921), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n928), .A2(new_n937), .ZN(G54));
  INV_X1    g752(.A(new_n477), .ZN(new_n939));
  NAND2_X1  g753(.A1(KEYINPUT58), .A2(G475), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n939), .B1(new_n911), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n929), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n911), .A2(new_n939), .A3(new_n940), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(G60));
  NAND2_X1  g758(.A1(G478), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT59), .Z(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n627), .B1(new_n865), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n935), .A2(new_n627), .A3(new_n947), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n907), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n948), .A2(new_n950), .ZN(G63));
  NAND2_X1  g765(.A1(G217), .A2(G902), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT121), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT60), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n910), .A2(new_n650), .A3(new_n954), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n955), .B(new_n907), .C1(KEYINPUT122), .C2(KEYINPUT61), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n910), .A2(new_n954), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n957), .A2(new_n601), .ZN(new_n958));
  NAND2_X1  g772(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n956), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n957), .A2(new_n601), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n907), .B1(KEYINPUT122), .B2(KEYINPUT61), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(new_n957), .B2(new_n650), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n959), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n961), .A2(new_n965), .ZN(G66));
  INV_X1    g780(.A(G224), .ZN(new_n967));
  OAI21_X1  g781(.A(G953), .B1(new_n194), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n613), .A2(new_n842), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n969), .A2(new_n822), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n968), .B1(new_n970), .B2(G953), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n635), .B(new_n255), .C1(G898), .C2(new_n187), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(G69));
  NAND2_X1  g787(.A1(new_n759), .A2(new_n720), .ZN(new_n974));
  NOR4_X1   g788(.A1(new_n789), .A2(new_n306), .A3(new_n790), .A4(new_n974), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n806), .A2(new_n770), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n778), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT123), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n799), .A2(new_n978), .A3(new_n738), .A4(new_n817), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n799), .A2(new_n738), .A3(new_n817), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(KEYINPUT123), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n977), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n469), .A2(new_n470), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n528), .B(new_n983), .Z(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n187), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n984), .B1(G900), .B2(new_n187), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n605), .A2(new_n612), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n766), .A2(new_n684), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n990), .B(new_n991), .C1(new_n839), .C2(new_n840), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n799), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n993), .A2(new_n806), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n810), .A2(new_n698), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n994), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n989), .B1(new_n999), .B2(new_n187), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT124), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n987), .A2(new_n1001), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1002), .ZN(new_n1005));
  OR2_X1    g819(.A1(new_n1003), .A2(new_n1002), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n1005), .B(new_n1006), .C1(new_n986), .C2(new_n1000), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n1004), .A2(new_n1007), .ZN(G72));
  NAND2_X1  g822(.A1(G472), .A2(G902), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT63), .Z(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(KEYINPUT125), .Z(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n999), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1012), .B1(new_n1013), .B2(new_n970), .ZN(new_n1014));
  INV_X1    g828(.A(new_n688), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n525), .A2(KEYINPUT127), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1016), .B(new_n545), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n1010), .ZN(new_n1018));
  OAI22_X1  g832(.A1(new_n1014), .A2(new_n1015), .B1(new_n864), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT126), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n529), .A2(new_n518), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n981), .A2(new_n979), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1022), .A2(new_n778), .A3(new_n970), .A4(new_n976), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1021), .B1(new_n1023), .B2(new_n1011), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1020), .B1(new_n1024), .B2(new_n906), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1012), .B1(new_n982), .B2(new_n970), .ZN(new_n1026));
  OAI211_X1 g840(.A(KEYINPUT126), .B(new_n929), .C1(new_n1026), .C2(new_n1021), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1019), .B1(new_n1025), .B2(new_n1027), .ZN(G57));
endmodule


