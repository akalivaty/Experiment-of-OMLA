//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 1 0 1 0 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n208), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n202), .A2(new_n203), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n213), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n210), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT64), .Z(new_n227));
  INV_X1    g0027(.A(KEYINPUT1), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n227), .A2(new_n228), .ZN(new_n230));
  AND3_X1   g0030(.A1(new_n219), .A2(new_n229), .A3(new_n230), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G68), .Z(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(KEYINPUT21), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n207), .A2(G45), .ZN(new_n248));
  OR2_X1    g0048(.A1(KEYINPUT5), .A2(G41), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT5), .A2(G41), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT65), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT65), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G33), .A3(G41), .ZN(new_n255));
  INV_X1    g0055(.A(new_n214), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n251), .A2(new_n257), .A3(G274), .ZN(new_n258));
  INV_X1    g0058(.A(G45), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G1), .ZN(new_n260));
  AND2_X1   g0060(.A1(KEYINPUT5), .A2(G41), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT5), .A2(G41), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n257), .A2(new_n263), .A3(G270), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G264), .A3(G1698), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(G257), .A3(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G303), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n272), .A2(new_n274), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n256), .A2(new_n252), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n266), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G169), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G116), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n214), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n291), .B(new_n285), .C1(G1), .C2(new_n268), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n288), .B1(new_n292), .B2(new_n287), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G283), .ZN(new_n294));
  INV_X1    g0094(.A(G97), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n294), .B(new_n208), .C1(G33), .C2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n287), .A2(G20), .ZN(new_n297));
  AND3_X1   g0097(.A1(new_n290), .A2(KEYINPUT84), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(KEYINPUT84), .B1(new_n290), .B2(new_n297), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n296), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(KEYINPUT20), .B(new_n296), .C1(new_n298), .C2(new_n299), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n293), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n247), .B1(new_n284), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n302), .A2(new_n303), .ZN(new_n306));
  INV_X1    g0106(.A(new_n293), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n308), .A2(KEYINPUT21), .A3(G169), .A4(new_n283), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n266), .A2(new_n282), .A3(G190), .ZN(new_n310));
  INV_X1    g0110(.A(new_n283), .ZN(new_n311));
  INV_X1    g0111(.A(G200), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n304), .B(new_n310), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n308), .A2(G179), .A3(new_n311), .ZN(new_n314));
  AND4_X1   g0114(.A1(new_n305), .A2(new_n309), .A3(new_n313), .A4(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G41), .ZN(new_n316));
  AOI21_X1  g0116(.A(G1), .B1(new_n316), .B2(new_n259), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n214), .B1(KEYINPUT65), .B2(new_n252), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(new_n255), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G238), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n257), .A2(G274), .A3(new_n317), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G226), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(G1698), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n275), .B2(new_n276), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT68), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(G33), .A2(G97), .ZN(new_n328));
  OAI211_X1 g0128(.A(G232), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n324), .B(KEYINPUT68), .C1(new_n276), .C2(new_n275), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n327), .A2(new_n328), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n281), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT69), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n331), .A2(KEYINPUT69), .A3(new_n281), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n322), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT13), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT71), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n322), .ZN(new_n339));
  AND3_X1   g0139(.A1(new_n331), .A2(KEYINPUT69), .A3(new_n281), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT69), .B1(new_n331), .B2(new_n281), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT71), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(new_n343), .A3(KEYINPUT13), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n337), .B(new_n339), .C1(new_n340), .C2(new_n341), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT70), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n346), .B(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n312), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n208), .A2(G33), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G77), .ZN(new_n352));
  NOR2_X1   g0152(.A1(G20), .A2(G33), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n291), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT11), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n356), .A2(KEYINPUT73), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(KEYINPUT73), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT12), .B1(new_n285), .B2(G68), .ZN(new_n359));
  OR3_X1    g0159(.A1(new_n285), .A2(KEYINPUT12), .A3(G68), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n286), .A2(new_n290), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n203), .B1(new_n207), .B2(G20), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n359), .A2(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n357), .A2(new_n358), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G190), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT72), .B1(new_n342), .B2(KEYINPUT13), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n346), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n336), .A2(KEYINPUT72), .A3(new_n337), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n365), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NOR3_X1   g0169(.A1(new_n349), .A2(new_n364), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G179), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n367), .B2(new_n368), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n346), .B(KEYINPUT70), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n338), .A2(new_n344), .ZN(new_n374));
  OAI21_X1  g0174(.A(G169), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n372), .B1(new_n375), .B2(KEYINPUT14), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n345), .A2(new_n348), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT14), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n377), .A2(KEYINPUT74), .A3(new_n378), .A4(G169), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n378), .B(G169), .C1(new_n373), .C2(new_n374), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT74), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n376), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n370), .B1(new_n383), .B2(new_n364), .ZN(new_n384));
  INV_X1    g0184(.A(new_n317), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n257), .A2(G232), .A3(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(G223), .A2(G1698), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n323), .B2(G1698), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n388), .A2(new_n271), .B1(G33), .B2(G87), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n321), .B(new_n386), .C1(new_n389), .C2(new_n280), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n390), .A2(new_n365), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(G200), .B2(new_n390), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT16), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n269), .A2(new_n208), .A3(new_n270), .ZN(new_n394));
  XNOR2_X1  g0194(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n277), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n203), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G58), .A2(G68), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT77), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT77), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n401), .A2(G58), .A3(G68), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n400), .A2(new_n402), .A3(new_n216), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G20), .ZN(new_n404));
  INV_X1    g0204(.A(G159), .ZN(new_n405));
  INV_X1    g0205(.A(new_n353), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n393), .B1(new_n398), .B2(new_n407), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n403), .A2(G20), .B1(G159), .B2(new_n353), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT76), .B1(new_n394), .B2(new_n395), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT7), .B1(new_n277), .B2(new_n208), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT7), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT75), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT75), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT7), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT76), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n417), .A2(new_n277), .A3(new_n418), .A4(new_n208), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G68), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n409), .B1(new_n412), .B2(new_n420), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n408), .B(new_n290), .C1(new_n421), .C2(new_n393), .ZN(new_n422));
  XNOR2_X1  g0222(.A(KEYINPUT8), .B(G58), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(new_n207), .B2(G20), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n424), .A2(new_n361), .B1(new_n286), .B2(new_n423), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n392), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT17), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n422), .A2(new_n425), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT78), .B1(new_n390), .B2(G179), .ZN(new_n430));
  INV_X1    g0230(.A(G169), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n390), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n323), .A2(G1698), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(G223), .B2(G1698), .ZN(new_n434));
  INV_X1    g0234(.A(G87), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n434), .A2(new_n277), .B1(new_n268), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(G274), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(new_n318), .B2(new_n255), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n436), .A2(new_n281), .B1(new_n438), .B2(new_n317), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT78), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n439), .A2(new_n440), .A3(new_n371), .A4(new_n386), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n430), .A2(new_n432), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n429), .A2(KEYINPUT18), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT79), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n429), .A2(new_n442), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT18), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n446), .A2(new_n444), .A3(new_n447), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n428), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n423), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n452), .A2(new_n351), .B1(G150), .B2(new_n353), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n204), .A2(G20), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n291), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n207), .A2(G20), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n361), .A2(G50), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(G50), .B2(new_n285), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT9), .ZN(new_n460));
  XNOR2_X1  g0260(.A(new_n459), .B(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n271), .A2(G222), .A3(new_n273), .ZN(new_n462));
  INV_X1    g0262(.A(G77), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n271), .A2(G1698), .ZN(new_n464));
  INV_X1    g0264(.A(G223), .ZN(new_n465));
  OAI221_X1 g0265(.A(new_n462), .B1(new_n463), .B2(new_n271), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n281), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n319), .A2(G226), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n467), .A2(new_n321), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G190), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n461), .B(new_n471), .C1(new_n312), .C2(new_n470), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n472), .B(KEYINPUT10), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n459), .B1(new_n469), .B2(new_n431), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n474), .A2(KEYINPUT66), .B1(new_n371), .B2(new_n470), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(KEYINPUT66), .B2(new_n474), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n271), .A2(G232), .A3(new_n273), .ZN(new_n477));
  INV_X1    g0277(.A(G107), .ZN(new_n478));
  INV_X1    g0278(.A(G238), .ZN(new_n479));
  OAI221_X1 g0279(.A(new_n477), .B1(new_n478), .B2(new_n271), .C1(new_n464), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n281), .ZN(new_n481));
  AOI22_X1  g0281(.A1(G244), .A2(new_n319), .B1(new_n438), .B2(new_n317), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G190), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n361), .A2(G77), .A3(new_n456), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(G77), .B2(new_n285), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n452), .A2(new_n353), .B1(G20), .B2(G77), .ZN(new_n488));
  XNOR2_X1  g0288(.A(KEYINPUT15), .B(G87), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n488), .B1(new_n489), .B2(new_n350), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n487), .B1(new_n490), .B2(new_n290), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n483), .A2(G200), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n485), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(G169), .B1(new_n481), .B2(new_n482), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT67), .B1(new_n495), .B2(new_n491), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n484), .A2(new_n371), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n495), .A2(KEYINPUT67), .A3(new_n491), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n494), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  AND4_X1   g0302(.A1(new_n451), .A2(new_n473), .A3(new_n476), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n384), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(G244), .B(new_n273), .C1(new_n275), .C2(new_n276), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT4), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n294), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G250), .A2(G1698), .ZN(new_n510));
  NAND2_X1  g0310(.A1(KEYINPUT4), .A2(G244), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n510), .B1(new_n511), .B2(G1698), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n509), .B1(new_n271), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n281), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n257), .A2(new_n263), .A3(G257), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n258), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(new_n517), .A3(G190), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT6), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n519), .A2(new_n295), .A3(G107), .ZN(new_n520));
  XNOR2_X1  g0320(.A(G97), .B(G107), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n520), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  OAI22_X1  g0322(.A1(new_n522), .A2(new_n208), .B1(new_n463), .B2(new_n406), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n478), .B1(new_n396), .B2(new_n397), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n290), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n285), .A2(G97), .ZN(new_n526));
  INV_X1    g0326(.A(new_n292), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n526), .B1(new_n527), .B2(G97), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n518), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT80), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n530), .B1(new_n514), .B2(new_n281), .ZN(new_n531));
  AOI211_X1 g0331(.A(KEYINPUT80), .B(new_n280), .C1(new_n508), .C2(new_n513), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n517), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n529), .B1(G200), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n515), .A2(KEYINPUT80), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n280), .B1(new_n508), .B2(new_n513), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n530), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT81), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n538), .A2(new_n539), .A3(new_n371), .A4(new_n517), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n371), .B(new_n517), .C1(new_n531), .C2(new_n532), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT81), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n524), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n521), .A2(new_n519), .ZN(new_n545));
  INV_X1    g0345(.A(new_n520), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(G20), .B1(G77), .B2(new_n353), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n291), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n528), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n258), .A2(new_n516), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n536), .A2(new_n551), .ZN(new_n552));
  OAI22_X1  g0352(.A1(new_n549), .A2(new_n550), .B1(G169), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n534), .B1(new_n543), .B2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(G257), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n556));
  OAI211_X1 g0356(.A(G250), .B(new_n273), .C1(new_n275), .C2(new_n276), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G294), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n281), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n257), .A2(new_n263), .A3(G264), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n562), .A2(new_n371), .A3(new_n258), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n560), .A2(new_n258), .A3(new_n561), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n431), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n208), .B(G87), .C1(new_n275), .C2(new_n276), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT22), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT22), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n271), .A2(new_n568), .A3(new_n208), .A4(G87), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G33), .A2(G116), .ZN(new_n571));
  OR3_X1    g0371(.A1(new_n571), .A2(KEYINPUT85), .A3(G20), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT23), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n208), .B2(G107), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n478), .A2(KEYINPUT23), .A3(G20), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(KEYINPUT85), .B1(new_n571), .B2(G20), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n572), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n570), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT24), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT24), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n570), .A2(new_n581), .A3(new_n578), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n291), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT25), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n285), .B2(G107), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n286), .A2(KEYINPUT25), .A3(new_n478), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n527), .A2(G107), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n563), .B(new_n565), .C1(new_n583), .C2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n564), .A2(new_n312), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n560), .A2(new_n365), .A3(new_n258), .A4(new_n561), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n570), .A2(new_n581), .A3(new_n578), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n581), .B1(new_n570), .B2(new_n578), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n290), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n592), .A2(new_n595), .A3(new_n587), .ZN(new_n596));
  AOI21_X1  g0396(.A(G250), .B1(new_n207), .B2(G45), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n437), .B2(new_n260), .ZN(new_n598));
  OAI211_X1 g0398(.A(G244), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n599));
  OAI211_X1 g0399(.A(G238), .B(new_n273), .C1(new_n275), .C2(new_n276), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n600), .A3(new_n571), .ZN(new_n601));
  AOI221_X4 g0401(.A(new_n365), .B1(new_n598), .B2(new_n257), .C1(new_n601), .C2(new_n281), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n281), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n598), .A2(new_n257), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n312), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n208), .B(G68), .C1(new_n275), .C2(new_n276), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT19), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n350), .B2(new_n295), .ZN(new_n609));
  NAND3_X1  g0409(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n610));
  NOR2_X1   g0410(.A1(G97), .A2(G107), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n208), .A2(new_n610), .B1(new_n611), .B2(new_n435), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT82), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n607), .B(new_n609), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n290), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n527), .A2(G87), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n489), .A2(new_n286), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n606), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n489), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n527), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n616), .A2(new_n622), .A3(new_n618), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(KEYINPUT83), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT83), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n616), .A2(new_n622), .A3(new_n625), .A4(new_n618), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n603), .A2(G179), .A3(new_n604), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n601), .A2(new_n281), .B1(new_n257), .B2(new_n598), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n627), .B1(new_n431), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n624), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  AND4_X1   g0430(.A1(new_n589), .A2(new_n596), .A3(new_n620), .A4(new_n630), .ZN(new_n631));
  AND4_X1   g0431(.A1(new_n315), .A2(new_n505), .A3(new_n555), .A4(new_n631), .ZN(G372));
  OR3_X1    g0432(.A1(new_n349), .A2(new_n364), .A3(new_n369), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n426), .B(KEYINPUT17), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n383), .A2(new_n364), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n499), .A2(new_n501), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n448), .A2(new_n443), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n473), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n551), .B1(new_n535), .B2(new_n537), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n539), .B1(new_n642), .B2(new_n371), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n541), .A2(KEYINPUT81), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n554), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n630), .A2(new_n620), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT26), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n629), .A2(new_n623), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n553), .B1(new_n540), .B2(new_n542), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n606), .A2(new_n619), .B1(new_n629), .B2(new_n623), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n647), .A2(new_n648), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n309), .A2(new_n305), .A3(new_n314), .ZN(new_n654));
  INV_X1    g0454(.A(new_n589), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n534), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n645), .A2(new_n657), .A3(new_n596), .A4(new_n651), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n656), .B1(new_n658), .B2(KEYINPUT86), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n651), .A2(new_n596), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n649), .A2(new_n660), .A3(new_n534), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT86), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n653), .B1(new_n659), .B2(new_n663), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n641), .B(new_n476), .C1(new_n504), .C2(new_n664), .ZN(G369));
  NAND3_X1  g0465(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n304), .A2(new_n672), .ZN(new_n673));
  MUX2_X1   g0473(.A(new_n315), .B(new_n654), .S(new_n673), .Z(new_n674));
  AND2_X1   g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n589), .A2(new_n596), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n672), .B1(new_n595), .B2(new_n587), .ZN(new_n677));
  OAI22_X1  g0477(.A1(new_n676), .A2(new_n677), .B1(new_n589), .B2(new_n672), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n654), .A2(new_n589), .A3(new_n596), .A4(new_n672), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n655), .A2(new_n672), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT87), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n680), .A2(KEYINPUT87), .A3(new_n681), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n679), .A2(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n211), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR4_X1   g0490(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G1), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n217), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n664), .A2(KEYINPUT29), .A3(new_n671), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT29), .ZN(new_n696));
  INV_X1    g0496(.A(new_n656), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n661), .ZN(new_n698));
  INV_X1    g0498(.A(new_n651), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT26), .B1(new_n645), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n646), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(new_n649), .A3(new_n650), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n648), .B(KEYINPUT91), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n698), .A2(new_n700), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n696), .B1(new_n704), .B2(new_n672), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n695), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n631), .A2(new_n555), .A3(new_n315), .A4(new_n672), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT90), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n552), .A2(G179), .A3(new_n282), .A4(new_n266), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT88), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n562), .A2(new_n711), .A3(new_n628), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n560), .A2(new_n561), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n603), .A2(new_n604), .ZN(new_n714));
  OAI21_X1  g0514(.A(KEYINPUT88), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n710), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT30), .B1(new_n716), .B2(KEYINPUT89), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT89), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n712), .A2(new_n715), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n718), .B(new_n719), .C1(new_n720), .C2(new_n710), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n311), .A2(G179), .A3(new_n628), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(new_n533), .A3(new_n564), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n717), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n671), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT31), .B1(new_n724), .B2(new_n671), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n709), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G330), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n706), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n694), .B1(new_n732), .B2(G1), .ZN(G364));
  INV_X1    g0533(.A(G13), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n207), .B1(new_n735), .B2(G45), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n689), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n675), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(G330), .B2(new_n674), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n214), .B1(G20), .B2(new_n431), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n365), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n208), .A2(new_n365), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n371), .A2(G200), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n745), .A2(new_n201), .B1(new_n748), .B2(new_n202), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n208), .A2(G190), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n747), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n751), .A2(KEYINPUT94), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(KEYINPUT94), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n749), .B1(new_n755), .B2(G77), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT95), .Z(new_n757));
  NAND3_X1  g0557(.A1(new_n746), .A2(new_n371), .A3(G200), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G87), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n750), .A2(new_n371), .A3(G200), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n760), .B(new_n271), .C1(new_n478), .C2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n743), .A2(G190), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G179), .A2(G200), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n208), .B1(new_n765), .B2(G190), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n764), .A2(new_n203), .B1(new_n766), .B2(new_n295), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n750), .A2(new_n765), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n405), .ZN(new_n769));
  XOR2_X1   g0569(.A(KEYINPUT96), .B(KEYINPUT32), .Z(new_n770));
  XNOR2_X1  g0570(.A(new_n769), .B(new_n770), .ZN(new_n771));
  OR4_X1    g0571(.A1(new_n757), .A2(new_n762), .A3(new_n767), .A4(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G322), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n277), .B1(new_n748), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n766), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n774), .B1(G294), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n751), .ZN(new_n777));
  INV_X1    g0577(.A(new_n768), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n777), .A2(G311), .B1(new_n778), .B2(G329), .ZN(new_n779));
  INV_X1    g0579(.A(new_n761), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G303), .A2(new_n759), .B1(new_n780), .B2(G283), .ZN(new_n781));
  XNOR2_X1  g0581(.A(KEYINPUT97), .B(G326), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT33), .B(G317), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n783), .A2(new_n744), .B1(new_n763), .B2(new_n784), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n776), .A2(new_n779), .A3(new_n781), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n742), .B1(new_n772), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n738), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n688), .A2(new_n277), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n789), .A2(G355), .B1(new_n287), .B2(new_n688), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n211), .A2(new_n277), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT92), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(G45), .B2(new_n217), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n245), .A2(new_n259), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n790), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G13), .A2(G33), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n741), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n788), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT93), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n787), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n800), .A2(new_n801), .ZN(new_n804));
  INV_X1    g0604(.A(new_n798), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n803), .B(new_n804), .C1(new_n674), .C2(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n740), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G396));
  NAND2_X1  g0608(.A1(new_n652), .A2(new_n648), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n650), .B1(new_n701), .B2(new_n649), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n697), .B1(new_n661), .B2(new_n662), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n658), .A2(KEYINPUT86), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n491), .A2(new_n672), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n493), .B(new_n815), .C1(new_n498), .C2(new_n500), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n637), .B2(new_n815), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n814), .A2(new_n672), .A3(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT100), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n814), .A2(KEYINPUT100), .A3(new_n672), .A4(new_n817), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n659), .A2(new_n663), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n671), .B1(new_n823), .B2(new_n811), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n822), .B1(new_n824), .B2(new_n817), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(new_n730), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n738), .B1(new_n825), .B2(new_n730), .ZN(new_n828));
  INV_X1    g0628(.A(new_n817), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n796), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n741), .A2(new_n796), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n738), .B1(G77), .B2(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n780), .A2(G87), .B1(new_n778), .B2(G311), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT98), .ZN(new_n835));
  INV_X1    g0635(.A(G294), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n277), .B1(new_n748), .B2(new_n836), .C1(new_n478), .C2(new_n758), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n755), .B2(G116), .ZN(new_n838));
  INV_X1    g0638(.A(G283), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n764), .A2(new_n839), .B1(new_n766), .B2(new_n295), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(G303), .B2(new_n744), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n835), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  AOI22_X1  g0642(.A1(G137), .A2(new_n744), .B1(new_n763), .B2(G150), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT99), .ZN(new_n844));
  INV_X1    g0644(.A(G143), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n844), .B1(new_n845), .B2(new_n748), .C1(new_n405), .C2(new_n754), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT34), .Z(new_n847));
  AOI22_X1  g0647(.A1(new_n780), .A2(G68), .B1(new_n778), .B2(G132), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n277), .B1(new_n759), .B2(G50), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n848), .B(new_n849), .C1(new_n202), .C2(new_n766), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n842), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n833), .B1(new_n851), .B2(new_n741), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n827), .A2(new_n828), .B1(new_n830), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(G384));
  OR2_X1    g0654(.A1(new_n547), .A2(KEYINPUT35), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n547), .A2(KEYINPUT35), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n855), .A2(G116), .A3(new_n215), .A4(new_n856), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT36), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n218), .A2(G77), .A3(new_n402), .A4(new_n400), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n859), .A2(KEYINPUT101), .B1(G50), .B2(new_n203), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(KEYINPUT101), .B2(new_n859), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n734), .A2(G1), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT40), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n707), .B(KEYINPUT90), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n724), .A2(new_n671), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT31), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n725), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n817), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n364), .A2(new_n671), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n636), .A2(new_n633), .A3(new_n870), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n364), .B(new_n671), .C1(new_n383), .C2(new_n370), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n425), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n421), .A2(KEYINPUT103), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT103), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n876), .B(new_n409), .C1(new_n412), .C2(new_n420), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n875), .A2(new_n393), .A3(new_n877), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n410), .A2(new_n411), .ZN(new_n879));
  INV_X1    g0679(.A(new_n420), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n407), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n291), .B1(new_n881), .B2(KEYINPUT16), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n874), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n442), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n426), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n883), .A2(new_n669), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT37), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n669), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n429), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n446), .A2(new_n889), .A3(new_n890), .A4(new_n426), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n290), .B1(new_n421), .B2(new_n393), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT16), .B1(new_n421), .B2(KEYINPUT103), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n893), .B1(new_n877), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n888), .B1(new_n895), .B2(new_n874), .ZN(new_n896));
  OAI211_X1 g0696(.A(KEYINPUT38), .B(new_n892), .C1(new_n451), .C2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT38), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n446), .A2(new_n889), .A3(new_n426), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(new_n890), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n889), .B1(new_n634), .B2(new_n639), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n863), .B1(new_n873), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n871), .A2(new_n872), .ZN(new_n905));
  INV_X1    g0705(.A(new_n869), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n449), .A2(new_n450), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n896), .B1(new_n907), .B2(new_n634), .ZN(new_n908));
  INV_X1    g0708(.A(new_n891), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n896), .B(new_n426), .C1(new_n884), .C2(new_n883), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n909), .B1(new_n910), .B2(KEYINPUT37), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n898), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT40), .B1(new_n912), .B2(new_n897), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n905), .A2(new_n906), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(G330), .B1(new_n904), .B2(new_n914), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n729), .A2(new_n384), .A3(G330), .A4(new_n503), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n917), .B(KEYINPUT104), .Z(new_n918));
  OAI211_X1 g0718(.A(new_n505), .B(new_n729), .C1(new_n904), .C2(new_n914), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n903), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n636), .A2(new_n671), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n912), .A2(KEYINPUT39), .A3(new_n897), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n640), .A2(new_n669), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n499), .A2(new_n501), .A3(new_n672), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n928), .B(KEYINPUT102), .Z(new_n929));
  AOI22_X1  g0729(.A1(new_n822), .A2(new_n929), .B1(new_n871), .B2(new_n872), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n912), .A2(new_n897), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n384), .B(new_n503), .C1(new_n695), .C2(new_n705), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n641), .A2(new_n476), .A3(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n932), .B(new_n934), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n920), .A2(new_n935), .B1(new_n207), .B2(new_n735), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n920), .A2(new_n935), .ZN(new_n937));
  OAI221_X1 g0737(.A(new_n858), .B1(new_n861), .B2(new_n862), .C1(new_n936), .C2(new_n937), .ZN(G367));
  NAND2_X1  g0738(.A1(new_n792), .A2(new_n238), .ZN(new_n939));
  INV_X1    g0739(.A(new_n799), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n688), .B2(new_n621), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n788), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n651), .B1(new_n619), .B2(new_n672), .ZN(new_n943));
  OR3_X1    g0743(.A1(new_n648), .A2(new_n619), .A3(new_n672), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(G150), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n271), .B1(new_n748), .B2(new_n946), .C1(new_n405), .C2(new_n764), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n780), .A2(G77), .ZN(new_n948));
  INV_X1    g0748(.A(G137), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n948), .B1(new_n202), .B2(new_n758), .C1(new_n949), .C2(new_n768), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n754), .A2(new_n201), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n775), .A2(G68), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n745), .B2(new_n845), .ZN(new_n953));
  OR4_X1    g0753(.A1(new_n947), .A2(new_n950), .A3(new_n951), .A4(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n758), .A2(new_n287), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n955), .A2(KEYINPUT46), .B1(new_n478), .B2(new_n766), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(G311), .B2(new_n744), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n755), .A2(G283), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n761), .A2(new_n295), .ZN(new_n959));
  INV_X1    g0759(.A(G303), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n277), .B1(new_n748), .B2(new_n960), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n959), .B(new_n961), .C1(G317), .C2(new_n778), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n955), .A2(KEYINPUT46), .B1(new_n763), .B2(G294), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n957), .A2(new_n958), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n954), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT109), .Z(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT47), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n942), .B1(new_n805), .B2(new_n945), .C1(new_n967), .C2(new_n742), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n679), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT105), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n645), .A2(new_n657), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n672), .B1(new_n525), .B2(new_n528), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n645), .A2(new_n672), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n971), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI221_X1 g0776(.A(KEYINPUT105), .B1(new_n645), .B2(new_n672), .C1(new_n972), .C2(new_n973), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n976), .A2(new_n684), .A3(new_n685), .A4(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT44), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n976), .A2(new_n977), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n686), .ZN(new_n981));
  XOR2_X1   g0781(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n980), .A2(new_n686), .A3(new_n982), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n970), .B1(new_n979), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT44), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n978), .B(new_n988), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n989), .A2(new_n679), .A3(new_n985), .A4(new_n984), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT107), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n654), .A2(new_n672), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n680), .B1(new_n678), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n675), .B(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n992), .B1(new_n731), .B2(new_n996), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n706), .A2(KEYINPUT107), .A3(new_n995), .A4(new_n730), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT108), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n991), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n997), .A2(KEYINPUT108), .A3(new_n998), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n731), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n689), .B(KEYINPUT41), .Z(new_n1004));
  OAI21_X1  g0804(.A(new_n736), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n680), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n980), .A2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT42), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n980), .A2(new_n655), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n671), .B1(new_n1010), .B2(new_n645), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1006), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n980), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n679), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1016), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n969), .B1(new_n1005), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(G387));
  OAI211_X1 g0823(.A(new_n999), .B(new_n689), .C1(new_n732), .C2(new_n995), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n748), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n1025), .A2(G317), .B1(G311), .B2(new_n763), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n773), .B2(new_n745), .C1(new_n754), .C2(new_n960), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT48), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n759), .A2(G294), .B1(new_n775), .B2(G283), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT49), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n277), .B1(new_n768), .B2(new_n782), .C1(new_n287), .C2(new_n761), .ZN(new_n1036));
  OR3_X1    g0836(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n758), .A2(new_n463), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n751), .A2(new_n203), .B1(new_n768), .B2(new_n946), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(G50), .C2(new_n1025), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n277), .B(new_n959), .C1(new_n452), .C2(new_n763), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n775), .A2(new_n621), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n744), .A2(G159), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n742), .B1(new_n1037), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n691), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n789), .A2(new_n1046), .B1(new_n478), .B2(new_n688), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n235), .A2(new_n259), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT110), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n691), .A2(KEYINPUT111), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n423), .A2(G50), .ZN(new_n1051));
  XOR2_X1   g0851(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1050), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n691), .A2(KEYINPUT111), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n259), .B1(new_n203), .B2(new_n463), .C1(new_n1053), .C2(new_n1051), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n792), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1047), .B1(new_n1049), .B2(new_n1058), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n788), .B(new_n1045), .C1(new_n799), .C2(new_n1059), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n678), .A2(new_n805), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1060), .A2(new_n1061), .B1(new_n995), .B2(new_n737), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1024), .A2(new_n1062), .ZN(G393));
  NAND2_X1  g0863(.A1(new_n999), .A2(new_n1000), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n991), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1064), .A2(new_n1002), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n690), .B1(new_n999), .B2(new_n991), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n991), .A2(KEYINPUT113), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n736), .B1(new_n991), .B2(KEYINPUT113), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1015), .A2(new_n798), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n792), .A2(new_n242), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n940), .B1(G97), .B2(new_n688), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n788), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT114), .Z(new_n1075));
  AOI22_X1  g0875(.A1(new_n1025), .A2(G311), .B1(G317), .B2(new_n744), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT52), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n758), .A2(new_n839), .B1(new_n768), .B2(new_n773), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT115), .Z(new_n1079));
  OAI221_X1 g0879(.A(new_n277), .B1(new_n751), .B2(new_n836), .C1(new_n478), .C2(new_n761), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n764), .A2(new_n960), .B1(new_n766), .B2(new_n287), .ZN(new_n1081));
  OR4_X1    g0881(.A1(new_n1077), .A2(new_n1079), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n758), .A2(new_n203), .B1(new_n768), .B2(new_n845), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n277), .B(new_n1083), .C1(G87), .C2(new_n780), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n745), .A2(new_n946), .B1(new_n748), .B2(new_n405), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT51), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n755), .A2(new_n452), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n775), .A2(G77), .B1(G50), .B2(new_n763), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1084), .A2(new_n1086), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n742), .B1(new_n1082), .B2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1075), .A2(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1069), .A2(new_n1070), .B1(new_n1071), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1068), .A2(new_n1092), .ZN(G390));
  INV_X1    g0893(.A(KEYINPUT118), .ZN(new_n1094));
  OAI211_X1 g0894(.A(G330), .B(new_n817), .C1(new_n864), .C2(new_n868), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n700), .A2(new_n702), .A3(new_n703), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n658), .A2(new_n656), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n672), .B(new_n817), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT116), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1099), .A2(new_n929), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1099), .A2(new_n929), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(KEYINPUT116), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n905), .A2(new_n1096), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1095), .A2(new_n871), .A3(new_n872), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT117), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1095), .A2(new_n871), .A3(KEYINPUT117), .A4(new_n872), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1104), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(KEYINPUT100), .B1(new_n824), .B2(new_n817), .ZN(new_n1110));
  NOR4_X1   g0910(.A1(new_n664), .A2(new_n819), .A3(new_n671), .A4(new_n829), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n929), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n1095), .A2(new_n871), .A3(new_n872), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1095), .B1(new_n871), .B2(new_n872), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1109), .A2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n641), .A2(new_n476), .A3(new_n933), .A4(new_n916), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1094), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  AOI211_X1 g0919(.A(KEYINPUT118), .B(new_n1117), .C1(new_n1109), .C2(new_n1115), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n923), .B1(new_n897), .B2(new_n902), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n905), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1103), .A2(new_n1101), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n923), .B1(new_n1112), .B2(new_n905), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n922), .A2(new_n924), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n1114), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1125), .B1(new_n1123), .B2(new_n1095), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1121), .A2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1129), .B(new_n1130), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(new_n1133), .A3(new_n689), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1127), .A2(new_n797), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n764), .A2(new_n949), .B1(new_n766), .B2(new_n405), .ZN(new_n1136));
  XOR2_X1   g0936(.A(KEYINPUT54), .B(G143), .Z(new_n1137));
  AOI21_X1  g0937(.A(new_n1136), .B1(new_n755), .B2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT119), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G132), .A2(new_n1025), .B1(new_n778), .B2(G125), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1140), .B(new_n271), .C1(new_n201), .C2(new_n761), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n758), .A2(KEYINPUT53), .A3(new_n946), .ZN(new_n1142));
  OAI21_X1  g0942(.A(KEYINPUT53), .B1(new_n758), .B2(new_n946), .ZN(new_n1143));
  INV_X1    g0943(.A(G128), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1143), .B1(new_n745), .B2(new_n1144), .ZN(new_n1145));
  NOR4_X1   g0945(.A1(new_n1139), .A2(new_n1141), .A3(new_n1142), .A4(new_n1145), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n780), .A2(G68), .B1(new_n778), .B2(G294), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1147), .B1(new_n287), .B2(new_n748), .C1(new_n754), .C2(new_n295), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n775), .A2(G77), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n760), .A2(new_n277), .A3(new_n1149), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n764), .A2(new_n478), .B1(new_n745), .B2(new_n839), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n1148), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n741), .B1(new_n1146), .B2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1153), .B(new_n738), .C1(new_n452), .C2(new_n832), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1135), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1131), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1155), .B1(new_n1156), .B2(new_n737), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1134), .A2(new_n1157), .ZN(G378));
  NAND2_X1  g0958(.A1(new_n473), .A2(new_n476), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n459), .A2(new_n669), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1159), .B(new_n1160), .Z(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n1161), .B(new_n1162), .Z(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(KEYINPUT122), .ZN(new_n1164));
  INV_X1    g0964(.A(G330), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n905), .A2(new_n903), .A3(new_n906), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(KEYINPUT40), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n873), .A2(new_n913), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1165), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1112), .A2(new_n931), .A3(new_n905), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1170), .A2(new_n925), .A3(new_n926), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n915), .A2(new_n932), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1164), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n915), .A2(new_n932), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1164), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n736), .B1(new_n1174), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1163), .A2(new_n796), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n738), .B1(G50), .B2(new_n832), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n1181), .B(KEYINPUT121), .Z(new_n1182));
  NAND2_X1  g0982(.A1(new_n277), .A2(new_n316), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1183), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1183), .B1(G283), .B2(new_n778), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1185), .B1(new_n478), .B2(new_n748), .C1(new_n489), .C2(new_n751), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1038), .B1(G58), .B2(new_n780), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G97), .A2(new_n763), .B1(new_n744), .B2(G116), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n952), .A3(new_n1188), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1186), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1184), .B1(new_n1190), .B2(KEYINPUT58), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT120), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n759), .A2(new_n1137), .B1(new_n1025), .B2(G128), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n777), .A2(G137), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n744), .A2(G125), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n775), .A2(G150), .B1(G132), .B2(new_n763), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1198));
  AOI211_X1 g0998(.A(G33), .B(G41), .C1(new_n778), .C2(G124), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n405), .B2(new_n761), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n1197), .B2(KEYINPUT59), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1198), .A2(new_n1201), .B1(new_n1190), .B2(KEYINPUT58), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1192), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1182), .B1(new_n1203), .B2(new_n741), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1180), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1179), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(KEYINPUT118), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1116), .A2(new_n1094), .A3(new_n1118), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1117), .B1(new_n1211), .B2(new_n1156), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1177), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1214));
  OAI21_X1  g1014(.A(KEYINPUT57), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n689), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1118), .B1(new_n1121), .B2(new_n1131), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1174), .A2(new_n1178), .ZN(new_n1218));
  AOI21_X1  g1018(.A(KEYINPUT57), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1207), .B1(new_n1216), .B2(new_n1219), .ZN(G375));
  INV_X1    g1020(.A(new_n1004), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1109), .A2(new_n1117), .A3(new_n1115), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1121), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1116), .A2(new_n737), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n738), .B1(G68), .B2(new_n832), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(G283), .A2(new_n1025), .B1(new_n778), .B2(G303), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1226), .B1(new_n295), .B2(new_n758), .C1(new_n754), .C2(new_n478), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(G116), .A2(new_n763), .B1(new_n744), .B2(G294), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n948), .A2(new_n1228), .A3(new_n1042), .A4(new_n277), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n759), .A2(G159), .B1(new_n778), .B2(G128), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1230), .B1(new_n949), .B2(new_n748), .C1(new_n946), .C2(new_n751), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n277), .B1(new_n780), .B2(G58), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1137), .A2(new_n763), .B1(G132), .B2(new_n744), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1232), .B(new_n1233), .C1(new_n201), .C2(new_n766), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n1227), .A2(new_n1229), .B1(new_n1231), .B2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1225), .B1(new_n1235), .B2(new_n741), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n905), .B2(new_n797), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1224), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1223), .A2(new_n1239), .ZN(G381));
  NOR4_X1   g1040(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1241), .A2(new_n1022), .A3(new_n1239), .A4(new_n1223), .ZN(new_n1242));
  OR3_X1    g1042(.A1(G375), .A2(new_n1242), .A3(G378), .ZN(G407));
  AND2_X1   g1043(.A1(new_n1134), .A2(new_n1157), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n670), .A2(G213), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G407), .B(G213), .C1(G375), .C2(new_n1247), .ZN(G409));
  INV_X1    g1048(.A(KEYINPUT124), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1022), .B2(G390), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(G393), .B(new_n807), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1016), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1018), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n997), .A2(KEYINPUT108), .A3(new_n998), .ZN(new_n1257));
  AOI21_X1  g1057(.A(KEYINPUT108), .B1(new_n997), .B2(new_n998), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1257), .A2(new_n1258), .A3(new_n991), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1221), .B1(new_n1259), .B2(new_n731), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1256), .B1(new_n1260), .B2(new_n736), .ZN(new_n1261));
  INV_X1    g1061(.A(G390), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1261), .A2(new_n969), .A3(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1004), .B1(new_n1066), .B2(new_n732), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1021), .B1(new_n1264), .B2(new_n737), .ZN(new_n1265));
  AOI21_X1  g1065(.A(G390), .B1(new_n1265), .B2(new_n968), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n1250), .A2(new_n1252), .B1(new_n1263), .B2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1262), .B1(new_n1261), .B2(new_n969), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1265), .A2(new_n968), .A3(G390), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1268), .A2(new_n1249), .A3(new_n1269), .A4(new_n1251), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1267), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT123), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1179), .B2(new_n1206), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1131), .B1(new_n1210), .B2(new_n1209), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1221), .B(new_n1218), .C1(new_n1274), .C2(new_n1117), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n737), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(KEYINPUT123), .A3(new_n1205), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1273), .A2(new_n1275), .A3(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1244), .ZN(new_n1279));
  OAI211_X1 g1079(.A(G378), .B(new_n1207), .C1(new_n1216), .C2(new_n1219), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1245), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1209), .A2(new_n1210), .A3(new_n1222), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1283), .A2(KEYINPUT60), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1222), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n689), .B1(new_n1285), .B2(KEYINPUT60), .ZN(new_n1286));
  OAI211_X1 g1086(.A(G384), .B(new_n1239), .C1(new_n1284), .C2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1286), .B1(new_n1283), .B2(KEYINPUT60), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n853), .B1(new_n1288), .B2(new_n1238), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1246), .A2(G2897), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1287), .A2(new_n1289), .A3(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1290), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT61), .B1(new_n1282), .B2(new_n1293), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1281), .A2(new_n1245), .A3(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(KEYINPUT62), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1294), .A2(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1296), .A2(KEYINPUT62), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1271), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT125), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1287), .A2(KEYINPUT63), .A3(new_n1289), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1281), .A2(new_n1245), .A3(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1270), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1269), .A2(KEYINPUT124), .ZN(new_n1305));
  AOI22_X1  g1105(.A1(new_n1305), .A2(new_n1251), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1303), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1246), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT63), .B1(new_n1309), .B2(new_n1295), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1301), .B1(new_n1311), .B2(new_n1294), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1271), .B1(new_n1309), .B2(new_n1302), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT63), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1296), .A2(new_n1314), .ZN(new_n1315));
  AND4_X1   g1115(.A1(new_n1301), .A2(new_n1294), .A3(new_n1313), .A4(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1300), .B1(new_n1312), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT126), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  OAI211_X1 g1119(.A(KEYINPUT126), .B(new_n1300), .C1(new_n1312), .C2(new_n1316), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(G405));
  XNOR2_X1  g1121(.A(G375), .B(G378), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1322), .B(new_n1295), .ZN(new_n1323));
  XNOR2_X1  g1123(.A(new_n1323), .B(new_n1307), .ZN(G402));
endmodule


