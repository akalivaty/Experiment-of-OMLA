//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1211, new_n1212, new_n1213,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n211), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n222), .B1(new_n202), .B2(new_n223), .C1(new_n203), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n213), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n216), .B(new_n221), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  NAND2_X1  g0047(.A1(G20), .A2(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT15), .B(G87), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n211), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  OAI221_X1 g0053(.A(new_n248), .B1(new_n249), .B2(new_n250), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n219), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n256), .B1(new_n210), .B2(G20), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G77), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n259), .B1(G77), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  OR2_X1    g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT66), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT66), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G1698), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  OAI221_X1 g0070(.A(new_n265), .B1(new_n224), .B2(new_n266), .C1(new_n270), .C2(new_n223), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n271), .B(new_n272), .C1(G107), .C2(new_n265), .ZN(new_n273));
  INV_X1    g0073(.A(G274), .ZN(new_n274));
  AND2_X1   g0074(.A1(G1), .A2(G13), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G45), .ZN(new_n279));
  AOI21_X1  g0079(.A(G1), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT65), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT65), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n277), .A2(new_n283), .A3(new_n280), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n272), .A2(new_n280), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G244), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n273), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G169), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n262), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n290), .A2(KEYINPUT68), .ZN(new_n291));
  AND2_X1   g0091(.A1(KEYINPUT67), .A2(G179), .ZN(new_n292));
  NOR2_X1   g0092(.A1(KEYINPUT67), .A2(G179), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n288), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n290), .A2(KEYINPUT68), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(G190), .ZN(new_n297));
  INV_X1    g0097(.A(new_n262), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(G200), .B2(new_n288), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n291), .A2(new_n296), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G223), .A2(G1698), .ZN(new_n301));
  INV_X1    g0101(.A(G222), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n265), .B(new_n301), .C1(new_n270), .C2(new_n302), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n303), .B(new_n272), .C1(G77), .C2(new_n265), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n286), .A2(G226), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(new_n285), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n289), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n260), .A2(G50), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(new_n258), .B2(G50), .ZN(new_n309));
  INV_X1    g0109(.A(G150), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n253), .A2(new_n250), .B1(new_n310), .B2(new_n252), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(G20), .B2(new_n204), .ZN(new_n312));
  INV_X1    g0112(.A(new_n256), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n309), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n294), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n307), .B(new_n314), .C1(new_n315), .C2(new_n306), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n306), .A2(G200), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT69), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT10), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT9), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n314), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n314), .A2(new_n321), .ZN(new_n323));
  INV_X1    g0123(.A(G190), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n306), .A2(new_n324), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n322), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n319), .A2(new_n320), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n320), .B1(new_n319), .B2(new_n326), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n300), .B(new_n316), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(KEYINPUT3), .A2(G33), .ZN(new_n330));
  NOR2_X1   g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT66), .B(G1698), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G226), .ZN(new_n334));
  NAND2_X1  g0134(.A1(G232), .A2(G1698), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n332), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(G33), .A2(G97), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n272), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n282), .A2(new_n284), .B1(G238), .B2(new_n286), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT13), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT13), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n339), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G200), .ZN(new_n346));
  INV_X1    g0146(.A(G77), .ZN(new_n347));
  OAI22_X1  g0147(.A1(new_n250), .A2(new_n347), .B1(new_n211), .B2(G68), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT70), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n348), .A2(new_n349), .B1(G50), .B2(new_n251), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n349), .B2(new_n348), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n256), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT11), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n351), .A2(KEYINPUT11), .A3(new_n256), .ZN(new_n355));
  INV_X1    g0155(.A(new_n260), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT12), .B1(new_n356), .B2(new_n203), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n356), .A2(KEYINPUT12), .A3(new_n203), .ZN(new_n358));
  AOI211_X1 g0158(.A(new_n357), .B(new_n358), .C1(G68), .C2(new_n258), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n354), .A2(new_n355), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n342), .A2(G190), .A3(new_n344), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n346), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT71), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n346), .A2(KEYINPUT71), .A3(new_n362), .A4(new_n361), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT14), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n345), .A2(new_n368), .A3(G169), .ZN(new_n369));
  INV_X1    g0169(.A(G179), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n369), .B1(new_n370), .B2(new_n345), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n368), .B1(new_n345), .B2(G169), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n360), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n367), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n329), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT74), .ZN(new_n376));
  AND2_X1   g0176(.A1(G226), .A2(G1698), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n265), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n377), .B1(new_n330), .B2(new_n331), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT74), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(G223), .B1(new_n330), .B2(new_n331), .ZN(new_n383));
  INV_X1    g0183(.A(G33), .ZN(new_n384));
  INV_X1    g0184(.A(G87), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n383), .A2(new_n270), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n272), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n282), .A2(new_n284), .B1(G232), .B2(new_n286), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n387), .A2(G190), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n275), .A2(new_n276), .ZN(new_n390));
  INV_X1    g0190(.A(new_n386), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(new_n391), .B2(new_n381), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n286), .A2(G232), .ZN(new_n393));
  INV_X1    g0193(.A(new_n284), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n283), .B1(new_n277), .B2(new_n280), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(G200), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n389), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT7), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(new_n265), .B2(G20), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT72), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n263), .A2(KEYINPUT7), .A3(new_n211), .A4(new_n264), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(G68), .B1(new_n403), .B2(new_n402), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n202), .A2(new_n203), .ZN(new_n408));
  NOR2_X1   g0208(.A1(G58), .A2(G68), .ZN(new_n409));
  OAI21_X1  g0209(.A(G20), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n251), .A2(G159), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n407), .A2(KEYINPUT16), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT73), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n401), .A2(new_n415), .A3(new_n403), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n332), .A2(new_n211), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(KEYINPUT73), .A3(new_n400), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(G68), .A3(new_n418), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n419), .A2(new_n413), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n256), .B(new_n414), .C1(new_n420), .C2(KEYINPUT16), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT17), .ZN(new_n422));
  INV_X1    g0222(.A(new_n253), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(new_n260), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n258), .B2(new_n423), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n399), .A2(new_n421), .A3(new_n422), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n414), .A2(new_n256), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT16), .B1(new_n419), .B2(new_n413), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n425), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT17), .B1(new_n429), .B2(new_n398), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(G169), .B1(new_n392), .B2(new_n396), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n386), .B1(new_n378), .B2(new_n380), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n388), .B(new_n315), .C1(new_n433), .C2(new_n390), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT75), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n435), .B1(new_n432), .B2(new_n434), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT18), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(new_n440), .A3(new_n429), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n432), .A2(new_n434), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT75), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(new_n429), .A3(new_n436), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT18), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n431), .A2(new_n441), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT76), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(new_n447), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n375), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n265), .A2(new_n211), .A3(G87), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n451), .B(KEYINPUT22), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n207), .A2(G20), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n453), .B(KEYINPUT23), .ZN(new_n454));
  OR2_X1    g0254(.A1(KEYINPUT83), .A2(G116), .ZN(new_n455));
  NAND2_X1  g0255(.A1(KEYINPUT83), .A2(G116), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(new_n384), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n454), .B1(new_n459), .B2(new_n211), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n452), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT24), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT24), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n452), .A2(new_n463), .A3(new_n460), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n313), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G257), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(new_n266), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n265), .A2(new_n467), .B1(G33), .B2(G294), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n265), .A2(new_n333), .A3(G250), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n390), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n210), .B(G45), .C1(new_n278), .C2(KEYINPUT5), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT5), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(G41), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n472), .A2(new_n277), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G264), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n390), .B1(new_n471), .B2(new_n474), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n470), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G190), .ZN(new_n481));
  INV_X1    g0281(.A(G200), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(new_n480), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n356), .A2(new_n207), .ZN(new_n484));
  OR2_X1    g0284(.A1(new_n484), .A2(KEYINPUT25), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(KEYINPUT25), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n210), .A2(G33), .ZN(new_n487));
  AND4_X1   g0287(.A1(new_n219), .A2(new_n260), .A3(new_n255), .A4(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n485), .B(new_n486), .C1(new_n207), .C2(new_n489), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n465), .A2(new_n483), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n480), .A2(G179), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n493), .B1(new_n289), .B2(new_n480), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(new_n465), .B2(new_n490), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  OAI221_X1 g0297(.A(new_n265), .B1(new_n477), .B2(new_n266), .C1(new_n270), .C2(new_n466), .ZN(new_n498));
  INV_X1    g0298(.A(G303), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n390), .B1(new_n332), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n478), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n498), .A2(new_n500), .B1(new_n501), .B2(G270), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n502), .A2(G179), .A3(new_n476), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n455), .A2(G20), .A3(new_n456), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G283), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n505), .B(new_n211), .C1(G33), .C2(new_n206), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n256), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT20), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n504), .A2(KEYINPUT20), .A3(new_n506), .A4(new_n256), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n488), .A2(G116), .B1(new_n458), .B2(new_n356), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n511), .A2(KEYINPUT86), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT86), .B1(new_n511), .B2(new_n512), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n503), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT87), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n503), .B(KEYINPUT87), .C1(new_n514), .C2(new_n513), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n513), .A2(new_n514), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n502), .A2(new_n476), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G200), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n520), .B(new_n522), .C1(new_n324), .C2(new_n521), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n289), .B1(new_n502), .B2(new_n476), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n513), .B2(new_n514), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT21), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT21), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n524), .B(new_n527), .C1(new_n513), .C2(new_n514), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n519), .A2(new_n523), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT88), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n517), .A2(new_n518), .B1(new_n526), .B2(new_n528), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(KEYINPUT88), .A3(new_n523), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n450), .A2(new_n497), .A3(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT81), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n260), .A2(G97), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n488), .B2(G97), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT77), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n541), .A2(KEYINPUT6), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G97), .A2(G107), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n542), .A2(new_n208), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT6), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT77), .ZN(new_n546));
  AND2_X1   g0346(.A1(G97), .A2(G107), .ZN(new_n547));
  NOR2_X1   g0347(.A1(G97), .A2(G107), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n206), .A2(KEYINPUT6), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n544), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT78), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n544), .A2(new_n549), .A3(KEYINPUT78), .A4(new_n550), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(G20), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n251), .A2(G77), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT79), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n416), .A2(G107), .A3(new_n418), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n555), .A2(KEYINPUT79), .A3(new_n556), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n540), .B1(new_n562), .B2(new_n256), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT80), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT4), .ZN(new_n565));
  OAI21_X1  g0365(.A(G244), .B1(new_n330), .B2(new_n331), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n565), .B1(new_n566), .B2(new_n270), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n265), .A2(new_n333), .A3(KEYINPUT4), .A4(G244), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n265), .A2(G250), .A3(G1698), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .A4(new_n505), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n272), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n390), .B(G257), .C1(new_n471), .C2(new_n474), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n476), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n564), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  AOI211_X1 g0375(.A(KEYINPUT80), .B(new_n573), .C1(new_n570), .C2(new_n272), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n289), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n573), .B1(new_n570), .B2(new_n272), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n294), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n563), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n561), .A2(new_n560), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT79), .B1(new_n555), .B2(new_n556), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n256), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n571), .A2(new_n574), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT80), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n578), .A2(new_n564), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(G190), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n585), .A2(G200), .ZN(new_n589));
  AND4_X1   g0389(.A1(new_n584), .A2(new_n588), .A3(new_n539), .A4(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n537), .B1(new_n581), .B2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n584), .A2(new_n588), .A3(new_n539), .A4(new_n589), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n592), .B(KEYINPUT81), .C1(new_n563), .C2(new_n580), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT85), .ZN(new_n595));
  INV_X1    g0395(.A(new_n249), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(new_n260), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n489), .A2(new_n385), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n265), .A2(new_n211), .A3(G68), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT19), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n250), .B2(new_n206), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n211), .B1(new_n337), .B2(new_n600), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n385), .A2(new_n206), .A3(new_n207), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT84), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT84), .B1(new_n602), .B2(new_n603), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n599), .B(new_n601), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  AOI211_X1 g0408(.A(new_n597), .B(new_n598), .C1(new_n608), .C2(new_n256), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n332), .A2(new_n224), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n610), .A2(new_n333), .B1(G33), .B2(new_n457), .ZN(new_n611));
  OAI21_X1  g0411(.A(KEYINPUT82), .B1(new_n566), .B2(new_n266), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT82), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n265), .A2(new_n613), .A3(G244), .A4(G1698), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n390), .B1(new_n611), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n210), .A2(G45), .ZN(new_n617));
  INV_X1    g0417(.A(G250), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n210), .A2(new_n274), .A3(G45), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n390), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(G200), .B1(new_n616), .B2(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n611), .A2(new_n615), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n621), .B1(new_n624), .B2(new_n390), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n609), .B(new_n623), .C1(new_n324), .C2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n597), .B1(new_n608), .B2(new_n256), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(new_n249), .B2(new_n489), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n294), .B(new_n621), .C1(new_n624), .C2(new_n390), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n289), .B1(new_n616), .B2(new_n622), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n594), .A2(new_n595), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n593), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n586), .A2(new_n587), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n636), .A2(new_n289), .B1(new_n294), .B2(new_n578), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n584), .A2(new_n539), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT81), .B1(new_n639), .B2(new_n592), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n633), .B1(new_n635), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT85), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n536), .B1(new_n634), .B2(new_n642), .ZN(G372));
  OR2_X1    g0443(.A1(new_n327), .A2(new_n328), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n291), .A2(new_n296), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n367), .A2(new_n645), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n646), .A2(new_n373), .B1(new_n430), .B2(new_n426), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n441), .A2(new_n445), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n644), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n316), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n491), .A2(new_n632), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n519), .A2(new_n529), .A3(new_n495), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n652), .A2(new_n653), .A3(new_n639), .A4(new_n592), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n581), .A2(KEYINPUT26), .A3(new_n633), .ZN(new_n655));
  AOI21_X1  g0455(.A(KEYINPUT26), .B1(new_n581), .B2(new_n633), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n654), .B(new_n631), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n450), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n651), .A2(new_n658), .ZN(G369));
  NAND3_X1  g0459(.A1(new_n210), .A2(new_n211), .A3(G13), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(new_n662), .A3(G213), .ZN(new_n663));
  INV_X1    g0463(.A(G343), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n535), .B1(new_n520), .B2(new_n666), .ZN(new_n667));
  OR3_X1    g0467(.A1(new_n533), .A2(new_n520), .A3(new_n666), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G330), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g0471(.A(new_n671), .B(KEYINPUT89), .Z(new_n672));
  INV_X1    g0472(.A(new_n465), .ZN(new_n673));
  INV_X1    g0473(.A(new_n490), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n666), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OAI22_X1  g0475(.A1(new_n496), .A2(new_n675), .B1(new_n495), .B2(new_n666), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n533), .A2(new_n665), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n497), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n495), .B2(new_n665), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n677), .A2(new_n681), .ZN(G399));
  INV_X1    g0482(.A(new_n214), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(G41), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G1), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n603), .A2(G116), .ZN(new_n687));
  OAI22_X1  g0487(.A1(new_n686), .A2(new_n687), .B1(new_n217), .B2(new_n685), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  AOI211_X1 g0489(.A(new_n665), .B(new_n496), .C1(new_n532), .C2(new_n534), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n595), .B1(new_n594), .B2(new_n633), .ZN(new_n691));
  AOI211_X1 g0491(.A(KEYINPUT85), .B(new_n632), .C1(new_n591), .C2(new_n593), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n480), .A2(G179), .A3(new_n502), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n625), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n695), .A2(new_n586), .A3(new_n587), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n480), .A2(new_n315), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n625), .A2(new_n699), .A3(new_n521), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n698), .B1(new_n578), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n696), .A2(new_n697), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n665), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT31), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n670), .B1(new_n693), .B2(new_n704), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n657), .A2(KEYINPUT29), .A3(new_n666), .ZN(new_n706));
  AOI21_X1  g0506(.A(KEYINPUT29), .B1(new_n657), .B2(new_n666), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n689), .B1(new_n709), .B2(G1), .ZN(G364));
  INV_X1    g0510(.A(G13), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G20), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n686), .B1(G45), .B2(new_n712), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n713), .A2(KEYINPUT90), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(KEYINPUT90), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n683), .A2(new_n332), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G355), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(G116), .B2(new_n214), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n683), .A2(new_n265), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n722), .B1(new_n279), .B2(new_n218), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n243), .A2(G45), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n720), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(G13), .A2(G33), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G20), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n219), .B1(G20), .B2(new_n289), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n717), .B1(new_n725), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(G311), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n294), .A2(new_n211), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G190), .A2(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n324), .A2(G200), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G322), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n733), .A2(new_n736), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n211), .A2(G179), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n735), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n265), .B1(new_n743), .B2(G329), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n741), .A2(G190), .A3(G200), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n744), .B1(new_n499), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n737), .A2(new_n370), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G294), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n741), .A2(new_n324), .A3(G200), .ZN(new_n751));
  INV_X1    g0551(.A(G283), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n749), .A2(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n740), .A2(new_n746), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n734), .A2(G200), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n324), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G326), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n755), .A2(G190), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  XOR2_X1   g0559(.A(KEYINPUT33), .B(G317), .Z(new_n760));
  OAI211_X1 g0560(.A(new_n754), .B(new_n757), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n202), .A2(new_n738), .B1(new_n736), .B2(new_n347), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(G50), .B2(new_n756), .ZN(new_n763));
  XOR2_X1   g0563(.A(new_n763), .B(KEYINPUT91), .Z(new_n764));
  NAND2_X1  g0564(.A1(new_n758), .A2(G68), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n265), .B1(new_n745), .B2(new_n385), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT92), .ZN(new_n767));
  INV_X1    g0567(.A(G159), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n742), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT32), .ZN(new_n770));
  INV_X1    g0570(.A(new_n751), .ZN(new_n771));
  AOI22_X1  g0571(.A1(G107), .A2(new_n771), .B1(new_n748), .B2(G97), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n765), .A2(new_n767), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n761), .B1(new_n764), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n732), .B1(new_n774), .B2(new_n729), .ZN(new_n775));
  INV_X1    g0575(.A(new_n669), .ZN(new_n776));
  INV_X1    g0576(.A(new_n728), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT93), .ZN(new_n779));
  INV_X1    g0579(.A(new_n672), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n717), .B1(new_n669), .B2(new_n670), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(G396));
  INV_X1    g0583(.A(new_n705), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n300), .B1(new_n262), .B2(new_n666), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n645), .A2(new_n298), .A3(new_n665), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n657), .A2(new_n666), .A3(new_n787), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n787), .B(KEYINPUT98), .Z(new_n789));
  AND2_X1   g0589(.A1(new_n657), .A2(new_n666), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n784), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n717), .B1(new_n784), .B2(new_n791), .ZN(new_n794));
  INV_X1    g0594(.A(new_n787), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n726), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n729), .A2(new_n726), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n717), .B1(G77), .B2(new_n797), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT94), .Z(new_n799));
  INV_X1    g0599(.A(new_n736), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n756), .A2(G303), .B1(new_n800), .B2(new_n457), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(new_n752), .B2(new_n759), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT95), .Z(new_n803));
  OAI22_X1  g0603(.A1(new_n385), .A2(new_n751), .B1(new_n745), .B2(new_n207), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n332), .B1(new_n742), .B2(new_n733), .C1(new_n749), .C2(new_n206), .ZN(new_n805));
  INV_X1    g0605(.A(new_n738), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n804), .B(new_n805), .C1(G294), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n808), .A2(KEYINPUT96), .ZN(new_n809));
  INV_X1    g0609(.A(G132), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n265), .B1(new_n742), .B2(new_n810), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n749), .A2(new_n202), .B1(new_n751), .B2(new_n203), .ZN(new_n812));
  INV_X1    g0612(.A(new_n745), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n811), .B(new_n812), .C1(G50), .C2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT97), .ZN(new_n815));
  AOI22_X1  g0615(.A1(G159), .A2(new_n800), .B1(new_n806), .B2(G143), .ZN(new_n816));
  INV_X1    g0616(.A(new_n756), .ZN(new_n817));
  INV_X1    g0617(.A(G137), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n816), .B1(new_n817), .B2(new_n818), .C1(new_n310), .C2(new_n759), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT34), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n815), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n808), .A2(KEYINPUT96), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n809), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n799), .B1(new_n825), .B2(new_n729), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n793), .A2(new_n794), .B1(new_n796), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G384));
  NOR2_X1   g0628(.A1(new_n712), .A2(new_n210), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n693), .A2(new_n704), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n450), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT101), .Z(new_n832));
  INV_X1    g0632(.A(KEYINPUT38), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT99), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n412), .B1(new_n404), .B2(new_n406), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n834), .B(new_n256), .C1(new_n835), .C2(KEYINPUT16), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n414), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT16), .ZN(new_n838));
  AOI21_X1  g0638(.A(KEYINPUT72), .B1(new_n417), .B2(new_n400), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n405), .B1(new_n839), .B2(new_n403), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n838), .B1(new_n840), .B2(new_n412), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n834), .B1(new_n841), .B2(new_n256), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n425), .B1(new_n837), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n663), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n446), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n399), .A2(new_n421), .A3(new_n425), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n429), .A2(new_n844), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n444), .A2(new_n849), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n439), .A2(new_n843), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n854), .A2(new_n845), .A3(new_n849), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n853), .B1(KEYINPUT37), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n833), .B1(new_n848), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n852), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n859), .A2(KEYINPUT38), .A3(new_n847), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n360), .A2(new_n665), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n374), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n862), .B1(new_n367), .B2(new_n373), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n795), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n535), .A2(new_n497), .A3(new_n666), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n642), .B2(new_n634), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT31), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n703), .B(new_n871), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n861), .B(new_n868), .C1(new_n870), .C2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT40), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n446), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n444), .A2(new_n849), .A3(new_n851), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n877), .A2(KEYINPUT37), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n876), .A2(new_n851), .B1(new_n878), .B2(new_n853), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n833), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n860), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n830), .A2(KEYINPUT40), .A3(new_n881), .A4(new_n868), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n875), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(G330), .B1(new_n832), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n884), .A2(KEYINPUT102), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n884), .A2(KEYINPUT102), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n885), .B(new_n886), .C1(new_n832), .C2(new_n883), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n864), .A2(new_n866), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n645), .A2(new_n666), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n889), .B1(new_n788), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n861), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n648), .A2(new_n663), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n373), .A2(new_n665), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n848), .A2(new_n856), .A3(new_n833), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT38), .B1(new_n859), .B2(new_n847), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT39), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT39), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n880), .A2(new_n899), .A3(new_n860), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n895), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT100), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n894), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n895), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n880), .A2(new_n899), .A3(new_n860), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n899), .B1(new_n857), .B2(new_n860), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n891), .A2(new_n861), .B1(new_n648), .B2(new_n663), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT100), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n903), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n707), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n657), .A2(KEYINPUT29), .A3(new_n666), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n911), .A2(new_n450), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n651), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n910), .B(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n829), .B1(new_n888), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n915), .B2(new_n888), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n553), .A2(new_n554), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT35), .ZN(new_n919));
  OAI211_X1 g0719(.A(G116), .B(new_n220), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n919), .B2(new_n918), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT36), .Z(new_n922));
  NOR3_X1   g0722(.A1(new_n408), .A2(new_n217), .A3(new_n347), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n203), .A2(G50), .ZN(new_n924));
  OAI211_X1 g0724(.A(G1), .B(new_n711), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n917), .A2(new_n922), .A3(new_n925), .ZN(G367));
  OAI211_X1 g0726(.A(new_n639), .B(new_n592), .C1(new_n563), .C2(new_n666), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n581), .A2(new_n665), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n930), .A2(new_n679), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n932), .A2(KEYINPUT42), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT103), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n609), .A2(new_n666), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n935), .A2(new_n628), .A3(new_n629), .A4(new_n630), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n632), .B2(new_n935), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n927), .A2(new_n495), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n665), .B1(new_n939), .B2(new_n639), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n932), .B2(KEYINPUT42), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n934), .A2(new_n938), .A3(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT104), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n942), .B(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n677), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n934), .A2(new_n941), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n937), .B(KEYINPUT43), .Z(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n944), .A2(new_n945), .A3(new_n929), .A4(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT105), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n944), .A2(new_n948), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n677), .B2(new_n930), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n684), .B(KEYINPUT41), .Z(new_n953));
  OAI21_X1  g0753(.A(new_n679), .B1(new_n676), .B2(new_n678), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n672), .B(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n709), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  OR3_X1    g0757(.A1(new_n681), .A2(KEYINPUT44), .A3(new_n929), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT44), .B1(new_n681), .B2(new_n929), .ZN(new_n959));
  AND3_X1   g0759(.A1(new_n681), .A2(KEYINPUT45), .A3(new_n929), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT45), .B1(new_n681), .B2(new_n929), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n958), .B(new_n959), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n677), .B(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n957), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n953), .B1(new_n964), .B2(new_n709), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n712), .A2(G45), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(G1), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT106), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n950), .B(new_n952), .C1(new_n965), .C2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n721), .A2(new_n239), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n971), .B(new_n730), .C1(new_n214), .C2(new_n249), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n716), .B1(new_n972), .B2(KEYINPUT107), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(KEYINPUT107), .B2(new_n972), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n265), .B1(new_n742), .B2(new_n818), .C1(new_n347), .C2(new_n751), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n749), .A2(new_n203), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n975), .B(new_n976), .C1(G58), .C2(new_n813), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n977), .B1(new_n201), .B2(new_n736), .C1(new_n310), .C2(new_n738), .ZN(new_n978));
  INV_X1    g0778(.A(G143), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n979), .A2(new_n817), .B1(new_n759), .B2(new_n768), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT46), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n458), .B2(new_n745), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n982), .B1(new_n738), .B2(new_n499), .C1(new_n752), .C2(new_n736), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n749), .A2(new_n207), .B1(new_n751), .B2(new_n206), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n265), .B1(new_n743), .B2(G317), .ZN(new_n985));
  NAND2_X1  g0785(.A1(KEYINPUT46), .A2(G116), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n985), .B1(new_n745), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(KEYINPUT108), .B(G311), .Z(new_n989));
  NAND2_X1  g0789(.A1(new_n756), .A2(new_n989), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n988), .B(new_n990), .C1(new_n750), .C2(new_n759), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n978), .A2(new_n980), .B1(new_n983), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT47), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n974), .B1(new_n993), .B2(new_n729), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n777), .B2(new_n937), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n970), .A2(new_n995), .ZN(G387));
  AOI22_X1  g0796(.A1(new_n718), .A2(new_n687), .B1(new_n207), .B2(new_n683), .ZN(new_n997));
  AOI211_X1 g0797(.A(G45), .B(new_n687), .C1(G68), .C2(G77), .ZN(new_n998));
  XNOR2_X1  g0798(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n423), .A2(new_n999), .A3(new_n201), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n999), .B1(new_n423), .B2(new_n201), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n721), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n236), .A2(new_n279), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n997), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n730), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n717), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n676), .A2(new_n777), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n332), .B1(new_n743), .B2(G150), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n347), .B2(new_n745), .C1(new_n206), .C2(new_n751), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT110), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n800), .A2(G68), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n806), .A2(G50), .B1(new_n596), .B2(new_n748), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G159), .A2(new_n756), .B1(new_n758), .B2(new_n423), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n265), .B1(new_n743), .B2(G326), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n749), .A2(new_n752), .B1(new_n745), .B2(new_n750), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G303), .A2(new_n800), .B1(new_n806), .B2(G317), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n758), .A2(new_n989), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(new_n739), .C2(new_n817), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT48), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1017), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n1021), .B2(new_n1020), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT49), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1016), .B1(new_n458), .B2(new_n751), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1015), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1007), .B(new_n1008), .C1(new_n729), .C2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n955), .B2(new_n969), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n956), .A2(new_n684), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n955), .A2(new_n709), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(G393));
  INV_X1    g0832(.A(new_n963), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n956), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n964), .A2(new_n1034), .A3(new_n684), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(KEYINPUT112), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT112), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1034), .A2(new_n964), .A3(new_n1037), .A4(new_n684), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n930), .A2(new_n728), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n730), .B1(new_n206), .B2(new_n214), .C1(new_n722), .C2(new_n246), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n717), .A2(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n756), .A2(G317), .B1(new_n806), .B2(G311), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT52), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n332), .B1(new_n742), .B2(new_n739), .C1(new_n207), .C2(new_n751), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n749), .A2(new_n458), .B1(new_n745), .B2(new_n752), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(G294), .C2(new_n800), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n499), .B2(new_n759), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n265), .B1(new_n742), .B2(new_n979), .C1(new_n385), .C2(new_n751), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n749), .A2(new_n347), .B1(new_n745), .B2(new_n203), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(new_n423), .C2(new_n800), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n201), .B2(new_n759), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n756), .A2(G150), .B1(new_n806), .B2(G159), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT51), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n1044), .A2(new_n1048), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT111), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1042), .B1(new_n1056), .B2(new_n729), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n963), .A2(new_n969), .B1(new_n1040), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1039), .A2(new_n1058), .ZN(G390));
  AOI21_X1  g0859(.A(new_n650), .B1(new_n708), .B2(new_n450), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n705), .A2(new_n450), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT113), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n705), .A2(new_n450), .ZN(new_n1064));
  OAI21_X1  g0864(.A(KEYINPUT113), .B1(new_n1064), .B2(new_n914), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n788), .A2(new_n890), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  OAI211_X1 g0867(.A(G330), .B(new_n787), .C1(new_n870), .C2(new_n872), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1067), .B1(new_n1068), .B2(new_n889), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n889), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n705), .B2(new_n789), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1068), .A2(new_n889), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n830), .A2(G330), .A3(new_n787), .A4(new_n1070), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1067), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1063), .B(new_n1065), .C1(new_n1072), .C2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n895), .B(new_n881), .C1(new_n1067), .C2(new_n889), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n898), .B(new_n900), .C1(new_n891), .C2(new_n904), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n1078), .A2(new_n1079), .A3(new_n1074), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1074), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n684), .B1(new_n1077), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT114), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1074), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1078), .A2(new_n1079), .A3(new_n1074), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1084), .B1(new_n1076), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n1066), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n705), .A2(new_n789), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n889), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1094), .A2(new_n1067), .A3(new_n1074), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1062), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1082), .A2(new_n1096), .A3(new_n1099), .A4(KEYINPUT114), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1083), .B1(new_n1090), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n898), .A2(new_n726), .A3(new_n900), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n717), .B1(new_n423), .B2(new_n797), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n332), .B1(new_n743), .B2(G125), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1104), .B1(new_n201), .B2(new_n751), .C1(new_n768), .C2(new_n749), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(G137), .B2(new_n758), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(KEYINPUT54), .B(G143), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT115), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n800), .A2(new_n1108), .B1(new_n806), .B2(G132), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n745), .A2(new_n310), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT53), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n756), .A2(G128), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1106), .A2(new_n1109), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n756), .A2(G283), .B1(new_n800), .B2(G97), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n207), .B2(new_n759), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT116), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n332), .B1(new_n742), .B2(new_n750), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(G87), .B2(new_n813), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(G68), .A2(new_n771), .B1(new_n748), .B2(G77), .ZN(new_n1119));
  INV_X1    g0919(.A(G116), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1118), .B(new_n1119), .C1(new_n1120), .C2(new_n738), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1113), .B1(new_n1116), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1103), .B1(new_n1122), .B2(new_n729), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1082), .A2(new_n969), .B1(new_n1102), .B2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT117), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1101), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(G378));
  NAND2_X1  g0927(.A1(new_n644), .A2(new_n316), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1128), .B(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n314), .A2(new_n844), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1130), .B(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1132), .A2(KEYINPUT119), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n902), .B1(new_n894), .B2(new_n901), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n875), .A2(G330), .A3(new_n882), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n907), .A2(new_n908), .A3(KEYINPUT100), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1136), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1134), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n883), .B(G330), .C1(new_n903), .C2(new_n909), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(new_n1133), .A3(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1140), .A2(new_n1143), .A3(new_n969), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n717), .B1(G50), .B2(new_n797), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n201), .B1(G33), .B2(G41), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n332), .B2(new_n278), .ZN(new_n1147));
  AOI211_X1 g0947(.A(G41), .B(new_n265), .C1(new_n743), .C2(G283), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n1148), .B1(new_n202), .B2(new_n751), .C1(new_n347), .C2(new_n745), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT118), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n800), .A2(new_n596), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n976), .B1(G107), .B2(new_n806), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G97), .A2(new_n758), .B1(new_n756), .B2(G116), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT58), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1147), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G125), .A2(new_n756), .B1(new_n758), .B2(G132), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n806), .A2(G128), .B1(G150), .B2(new_n748), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n800), .A2(G137), .B1(new_n1108), .B2(new_n813), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1160), .A2(KEYINPUT59), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(KEYINPUT59), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n771), .A2(G159), .ZN(new_n1163));
  AOI211_X1 g0963(.A(G33), .B(G41), .C1(new_n743), .C2(G124), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1156), .B1(new_n1155), .B2(new_n1154), .C1(new_n1161), .C2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1145), .B1(new_n1166), .B2(new_n729), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1132), .B2(new_n727), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1144), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT57), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT120), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1065), .A2(KEYINPUT120), .A3(new_n1063), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n1090), .B2(new_n1100), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1171), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1176), .A2(new_n1171), .A3(new_n1177), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n684), .B(new_n1178), .C1(new_n1179), .C2(KEYINPUT121), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT121), .ZN(new_n1181));
  NOR4_X1   g0981(.A1(new_n1176), .A2(new_n1177), .A3(new_n1181), .A4(new_n1171), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1170), .B1(new_n1180), .B2(new_n1182), .ZN(G375));
  OAI211_X1 g0983(.A(new_n1092), .B(new_n1095), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n953), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1184), .A2(new_n1076), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n889), .A2(new_n726), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT122), .Z(new_n1188));
  OAI21_X1  g0988(.A(new_n717), .B1(G68), .B2(new_n797), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n749), .A2(new_n249), .B1(new_n206), .B2(new_n745), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n332), .B1(new_n742), .B2(new_n499), .C1(new_n347), .C2(new_n751), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n207), .B2(new_n736), .C1(new_n752), .C2(new_n738), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n750), .A2(new_n817), .B1(new_n759), .B2(new_n458), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(G150), .A2(new_n800), .B1(new_n806), .B2(G137), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n751), .A2(new_n202), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n332), .B(new_n1196), .C1(G128), .C2(new_n743), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(G159), .A2(new_n813), .B1(new_n748), .B2(G50), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n758), .A2(new_n1108), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n817), .B2(new_n810), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n1193), .A2(new_n1194), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1189), .B1(new_n729), .B2(new_n1202), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1096), .A2(new_n969), .B1(new_n1188), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1186), .A2(new_n1204), .ZN(G381));
  NOR2_X1   g1005(.A1(G375), .A2(G378), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n970), .A2(new_n1039), .A3(new_n995), .A4(new_n1058), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NOR4_X1   g1008(.A1(G393), .A2(G396), .A3(G384), .A4(G381), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1206), .A2(new_n1208), .A3(new_n1209), .ZN(G407));
  NAND3_X1  g1010(.A1(new_n1206), .A2(G213), .A3(new_n664), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(G407), .A2(new_n1211), .A3(G213), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT123), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1212), .B(new_n1213), .ZN(G409));
  NAND2_X1  g1014(.A1(G387), .A2(G390), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n1207), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(G393), .B(new_n782), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1217), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1215), .A2(new_n1207), .A3(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(G378), .B(new_n1170), .C1(new_n1180), .C2(new_n1182), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1176), .A2(new_n953), .A3(new_n1177), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1126), .B1(new_n1223), .B2(new_n1169), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT62), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n664), .A2(G213), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT60), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1184), .A2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1184), .B1(new_n1077), .B2(new_n1228), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT124), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n684), .B(new_n1229), .C1(new_n1230), .C2(new_n1231), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1204), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n827), .ZN(new_n1235));
  OAI211_X1 g1035(.A(G384), .B(new_n1204), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .A4(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT61), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1222), .A2(new_n1224), .B1(G213), .B2(new_n664), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1237), .A2(G213), .A3(new_n664), .A4(G2897), .ZN(new_n1242));
  INV_X1    g1042(.A(G2897), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1235), .B(new_n1236), .C1(new_n1243), .C2(new_n1227), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1239), .B(new_n1240), .C1(new_n1241), .C2(new_n1245), .ZN(new_n1246));
  XOR2_X1   g1046(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n1241), .B2(new_n1238), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1221), .B1(new_n1246), .B2(new_n1248), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT61), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1215), .A2(new_n1207), .A3(new_n1219), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1219), .B1(new_n1215), .B2(new_n1207), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT63), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n1251), .B2(new_n1237), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1241), .A2(KEYINPUT63), .A3(new_n1238), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1252), .A2(new_n1255), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1249), .A2(new_n1259), .ZN(G405));
  INV_X1    g1060(.A(KEYINPUT126), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1218), .A2(KEYINPUT126), .A3(new_n1220), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(G375), .A2(new_n1126), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1264), .A2(new_n1237), .A3(new_n1222), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1237), .B1(new_n1264), .B2(new_n1222), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1262), .B(new_n1263), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1268), .A2(new_n1255), .A3(KEYINPUT126), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(G402));
endmodule


