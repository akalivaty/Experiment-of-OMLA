//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n495, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n579, new_n580,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n633, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1233, new_n1234;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT65), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT66), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT71), .ZN(new_n462));
  NAND2_X1  g037(.A1(G101), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  AND3_X1   g040(.A1(new_n465), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n466));
  AOI21_X1  g041(.A(KEYINPUT68), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT69), .A2(KEYINPUT3), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT69), .A2(KEYINPUT3), .ZN(new_n470));
  OAI21_X1  g045(.A(G2104), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g048(.A(KEYINPUT70), .B(G2104), .C1(new_n469), .C2(new_n470), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n468), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n464), .B1(new_n475), .B2(G137), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n462), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n468), .ZN(new_n478));
  XNOR2_X1  g053(.A(KEYINPUT69), .B(KEYINPUT3), .ZN(new_n479));
  AOI21_X1  g054(.A(KEYINPUT70), .B1(new_n479), .B2(G2104), .ZN(new_n480));
  INV_X1    g055(.A(new_n474), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n478), .B(G137), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(new_n463), .ZN(new_n483));
  INV_X1    g058(.A(G2105), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n483), .A2(KEYINPUT71), .A3(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(KEYINPUT3), .B(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G125), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n487), .B(new_n488), .ZN(new_n489));
  AND2_X1   g064(.A1(G113), .A2(G2104), .ZN(new_n490));
  OAI21_X1  g065(.A(G2105), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n477), .A2(new_n485), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT72), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n477), .A2(new_n485), .A3(KEYINPUT72), .A4(new_n491), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(G160));
  NAND2_X1  g071(.A1(new_n475), .A2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(KEYINPUT73), .A3(G124), .ZN(new_n499));
  INV_X1    g074(.A(new_n475), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G136), .ZN(new_n502));
  OR2_X1    g077(.A1(G100), .A2(G2105), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n503), .B(G2104), .C1(G112), .C2(new_n484), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n505));
  INV_X1    g080(.A(G124), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n497), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n499), .A2(new_n502), .A3(new_n504), .A4(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G162));
  NAND2_X1  g084(.A1(new_n473), .A2(new_n474), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(G126), .A3(new_n478), .ZN(new_n511));
  NAND2_X1  g086(.A1(G114), .A2(G2104), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n484), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT4), .A2(G138), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n510), .A2(new_n484), .A3(new_n478), .A4(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n486), .A2(G138), .A3(new_n484), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT4), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n465), .A2(G2105), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n516), .A2(new_n517), .B1(G102), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n513), .A2(new_n520), .ZN(G164));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n523), .B2(KEYINPUT74), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT74), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n525), .A2(KEYINPUT6), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n527), .A2(G50), .ZN(new_n528));
  AND2_X1   g103(.A1(G75), .A2(G651), .ZN(new_n529));
  OAI21_X1  g104(.A(G543), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G543), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT5), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT5), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n523), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G62), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT75), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n524), .A2(new_n526), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n539), .B2(new_n535), .ZN(new_n540));
  INV_X1    g115(.A(new_n535), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n541), .A2(new_n527), .A3(KEYINPUT75), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G88), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n530), .B(new_n537), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(G166));
  NAND3_X1  g121(.A1(new_n540), .A2(G89), .A3(new_n542), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n536), .A2(G63), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n539), .A2(new_n531), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G51), .ZN(new_n550));
  NAND3_X1  g125(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT7), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n547), .A2(new_n548), .A3(new_n550), .A4(new_n552), .ZN(G286));
  INV_X1    g128(.A(G286), .ZN(G168));
  NAND2_X1  g129(.A1(G77), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G64), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n535), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  XOR2_X1   g133(.A(KEYINPUT76), .B(G52), .Z(new_n559));
  NAND2_X1  g134(.A1(new_n549), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g135(.A(KEYINPUT77), .B(G90), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n558), .B(new_n560), .C1(new_n543), .C2(new_n562), .ZN(G301));
  INV_X1    g138(.A(G301), .ZN(G171));
  AND2_X1   g139(.A1(new_n540), .A2(new_n542), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n565), .A2(G81), .B1(G43), .B2(new_n549), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT78), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n541), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(new_n523), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n549), .A2(G43), .ZN(new_n571));
  INV_X1    g146(.A(G81), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n569), .B(new_n571), .C1(new_n543), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(KEYINPUT78), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G860), .ZN(G153));
  AND3_X1   g151(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G36), .ZN(G176));
  NAND2_X1  g153(.A1(G1), .A2(G3), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT8), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(new_n580), .ZN(G188));
  AND3_X1   g156(.A1(new_n540), .A2(G91), .A3(new_n542), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n527), .A2(G53), .A3(G543), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT9), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n583), .B(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(G65), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(G65), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n541), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(G78), .A2(G543), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n523), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR3_X1   g167(.A1(new_n582), .A2(new_n586), .A3(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G299));
  XNOR2_X1  g169(.A(new_n545), .B(KEYINPUT81), .ZN(G303));
  OAI21_X1  g170(.A(G651), .B1(new_n541), .B2(G74), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n549), .A2(G49), .ZN(new_n597));
  INV_X1    g172(.A(G87), .ZN(new_n598));
  OAI211_X1 g173(.A(new_n596), .B(new_n597), .C1(new_n543), .C2(new_n598), .ZN(G288));
  NAND2_X1  g174(.A1(G73), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G61), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n535), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G651), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n565), .A2(G86), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n549), .A2(G48), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(G305));
  NAND2_X1  g183(.A1(new_n565), .A2(G85), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n541), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n610), .A2(new_n523), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n549), .A2(G47), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n609), .A2(new_n611), .A3(new_n612), .ZN(G290));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  OR3_X1    g189(.A1(G171), .A2(KEYINPUT83), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(KEYINPUT83), .B1(G171), .B2(new_n614), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n565), .A2(new_n617), .A3(G92), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT84), .ZN(new_n620));
  INV_X1    g195(.A(G66), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n535), .ZN(new_n622));
  AOI22_X1  g197(.A1(G54), .A2(new_n549), .B1(new_n622), .B2(G651), .ZN(new_n623));
  INV_X1    g198(.A(G92), .ZN(new_n624));
  OAI21_X1  g199(.A(KEYINPUT10), .B1(new_n543), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n618), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n615), .B(new_n616), .C1(G868), .C2(new_n627), .ZN(G284));
  OAI211_X1 g203(.A(new_n615), .B(new_n616), .C1(G868), .C2(new_n627), .ZN(G321));
  NAND2_X1  g204(.A1(G286), .A2(G868), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n593), .B2(G868), .ZN(G297));
  OAI21_X1  g206(.A(new_n630), .B1(new_n593), .B2(G868), .ZN(G280));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n627), .B1(new_n633), .B2(G860), .ZN(G148));
  NAND2_X1  g209(.A1(new_n627), .A2(new_n633), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G868), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(G868), .B2(new_n575), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g213(.A1(new_n501), .A2(G135), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n498), .A2(G123), .ZN(new_n640));
  OR2_X1    g215(.A1(G99), .A2(G2105), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n641), .B(G2104), .C1(G111), .C2(new_n484), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n486), .A2(new_n518), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT85), .B(KEYINPUT12), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT13), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2100), .Z(new_n649));
  NAND2_X1  g224(.A1(new_n644), .A2(new_n649), .ZN(G156));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2430), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2435), .ZN(new_n652));
  XOR2_X1   g227(.A(G2427), .B(G2438), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(KEYINPUT14), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2451), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n661), .B(new_n662), .Z(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(G14), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G401));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2072), .B(G2078), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT18), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n667), .B(KEYINPUT87), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT17), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n666), .B2(new_n668), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n667), .A2(new_n668), .ZN(new_n674));
  MUX2_X1   g249(.A(new_n674), .B(new_n668), .S(new_n666), .Z(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n670), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT88), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2096), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n679), .A2(G2100), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(G2100), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1956), .B(G2474), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT89), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1961), .B(G1966), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT90), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n686), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT20), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n685), .A2(new_n688), .A3(new_n690), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(new_n688), .B2(new_n690), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n686), .A2(KEYINPUT91), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n692), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1981), .B(G1986), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n698), .A2(new_n700), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n683), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n703), .ZN(new_n705));
  INV_X1    g280(.A(new_n683), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n705), .A2(new_n706), .A3(new_n701), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(G1991), .B(G1996), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT92), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n708), .B(new_n710), .ZN(G229));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G25), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n510), .A2(G119), .A3(G2105), .A4(new_n478), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT93), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n475), .A2(G131), .A3(new_n484), .ZN(new_n717));
  OR2_X1    g292(.A1(G95), .A2(G2105), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n718), .B(G2104), .C1(G107), .C2(new_n484), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n475), .A2(KEYINPUT93), .A3(G119), .A4(G2105), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n716), .A2(new_n717), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n713), .B1(new_n722), .B2(new_n712), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT35), .B(G1991), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT94), .Z(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n723), .B(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(G16), .A2(G24), .ZN(new_n728));
  INV_X1    g303(.A(G290), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(G16), .ZN(new_n730));
  INV_X1    g305(.A(G1986), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G16), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G6), .ZN(new_n734));
  AND3_X1   g309(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n733), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT32), .B(G1981), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT95), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n736), .B(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  MUX2_X1   g315(.A(G23), .B(G288), .S(G16), .Z(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT33), .B(G1976), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n733), .A2(G22), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G166), .B2(new_n733), .ZN(new_n745));
  INV_X1    g320(.A(G1971), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  OR3_X1    g323(.A1(new_n740), .A2(KEYINPUT96), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(KEYINPUT96), .B1(new_n740), .B2(new_n748), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n751), .A2(KEYINPUT34), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT34), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n749), .B2(new_n750), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n727), .B(new_n732), .C1(new_n752), .C2(new_n754), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n755), .A2(KEYINPUT36), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n755), .A2(KEYINPUT36), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(G16), .A2(G19), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n575), .B2(G16), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(G1341), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n486), .A2(G127), .ZN(new_n762));
  INV_X1    g337(.A(G115), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(new_n465), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G2105), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n510), .A2(G139), .A3(new_n484), .A4(new_n478), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n518), .A2(G103), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT25), .Z(new_n768));
  AND3_X1   g343(.A1(new_n766), .A2(KEYINPUT99), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(KEYINPUT99), .B1(new_n766), .B2(new_n768), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n765), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G29), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT98), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G29), .B2(G33), .ZN(new_n775));
  OR3_X1    g350(.A1(new_n774), .A2(G29), .A3(G33), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n773), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(KEYINPUT100), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT100), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n773), .A2(new_n779), .A3(new_n775), .A4(new_n776), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G2072), .ZN(new_n782));
  NOR2_X1   g357(.A1(G27), .A2(G29), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G164), .B2(G29), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(G2078), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n475), .A2(G141), .A3(new_n484), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n510), .A2(G129), .A3(G2105), .A4(new_n478), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n518), .A2(G105), .ZN(new_n788));
  NAND3_X1  g363(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT26), .Z(new_n790));
  NAND4_X1  g365(.A1(new_n786), .A2(new_n787), .A3(new_n788), .A4(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G29), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G29), .B2(G32), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT27), .B(G1996), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AND4_X1   g371(.A1(new_n761), .A2(new_n782), .A3(new_n785), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(G286), .A2(G16), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n733), .A2(G21), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(KEYINPUT102), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT102), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n798), .A2(new_n802), .A3(new_n799), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT30), .B(G28), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n804), .A2(G1966), .B1(new_n712), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT31), .B(G11), .ZN(new_n807));
  NAND2_X1  g382(.A1(G171), .A2(G16), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G5), .B2(G16), .ZN(new_n809));
  INV_X1    g384(.A(G1961), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AND3_X1   g386(.A1(new_n806), .A2(new_n807), .A3(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(G1966), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n801), .A2(new_n813), .A3(new_n803), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT103), .Z(new_n815));
  INV_X1    g390(.A(KEYINPUT104), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n643), .A2(new_n712), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n812), .A2(new_n815), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n806), .A2(new_n818), .A3(new_n807), .A4(new_n811), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n814), .B(KEYINPUT103), .ZN(new_n821));
  OAI21_X1  g396(.A(KEYINPUT104), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n712), .A2(G26), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n510), .A2(G128), .A3(G2105), .A4(new_n478), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(KEYINPUT97), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n475), .A2(G140), .A3(new_n484), .ZN(new_n827));
  OR2_X1    g402(.A1(G104), .A2(G2105), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n828), .B(G2104), .C1(G116), .C2(new_n484), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT97), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n475), .A2(new_n830), .A3(G128), .A4(G2105), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n826), .A2(new_n827), .A3(new_n829), .A4(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n824), .B1(new_n833), .B2(new_n712), .ZN(new_n834));
  MUX2_X1   g409(.A(new_n824), .B(new_n834), .S(KEYINPUT28), .Z(new_n835));
  INV_X1    g410(.A(G2067), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n712), .A2(G35), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(G162), .B2(new_n712), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT29), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n840), .A2(G2090), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n797), .A2(new_n823), .A3(new_n837), .A4(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n781), .A2(G2072), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT101), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n840), .A2(G2090), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n809), .A2(new_n810), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n733), .A2(G4), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n627), .B2(new_n733), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(G1348), .Z(new_n849));
  NAND3_X1  g424(.A1(new_n733), .A2(KEYINPUT23), .A3(G20), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT23), .ZN(new_n851));
  INV_X1    g426(.A(G20), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n851), .B1(new_n852), .B2(G16), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n850), .B(new_n853), .C1(new_n593), .C2(new_n733), .ZN(new_n854));
  INV_X1    g429(.A(G1956), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n845), .A2(new_n846), .A3(new_n849), .A4(new_n856), .ZN(new_n857));
  OAI22_X1  g432(.A1(new_n794), .A2(new_n795), .B1(G2078), .B2(new_n784), .ZN(new_n858));
  NOR4_X1   g433(.A1(new_n842), .A2(new_n844), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT24), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n860), .A2(G34), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(G34), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n861), .A2(new_n862), .A3(new_n712), .ZN(new_n863));
  INV_X1    g438(.A(G160), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n864), .B2(new_n712), .ZN(new_n865));
  INV_X1    g440(.A(G2084), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n859), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT105), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n859), .A2(KEYINPUT105), .A3(new_n868), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n758), .B1(new_n871), .B2(new_n872), .ZN(G311));
  AND3_X1   g448(.A1(new_n859), .A2(KEYINPUT105), .A3(new_n868), .ZN(new_n874));
  AOI21_X1  g449(.A(KEYINPUT105), .B1(new_n859), .B2(new_n868), .ZN(new_n875));
  OAI22_X1  g450(.A1(new_n874), .A2(new_n875), .B1(new_n756), .B2(new_n757), .ZN(G150));
  NAND2_X1  g451(.A1(new_n565), .A2(G93), .ZN(new_n877));
  AOI22_X1  g452(.A1(new_n541), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(new_n523), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n549), .A2(G55), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n877), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(G860), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(KEYINPUT37), .Z(new_n883));
  NAND2_X1  g458(.A1(new_n575), .A2(new_n881), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n881), .B1(new_n569), .B2(new_n566), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT39), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n627), .A2(G559), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT38), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n888), .B(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n883), .B1(new_n891), .B2(G860), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT106), .ZN(G145));
  INV_X1    g468(.A(G37), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT107), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n511), .A2(new_n512), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(G2105), .ZN(new_n897));
  INV_X1    g472(.A(new_n520), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n513), .A2(new_n520), .A3(KEYINPUT107), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n792), .A2(new_n832), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n827), .A2(new_n829), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n904), .A2(new_n791), .A3(new_n826), .A4(new_n831), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n903), .A2(new_n771), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n771), .B1(new_n903), .B2(new_n905), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n902), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n903), .A2(new_n905), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n772), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n903), .A2(new_n905), .A3(new_n771), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n901), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n647), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n475), .A2(G130), .A3(G2105), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n475), .A2(G142), .A3(new_n484), .ZN(new_n916));
  OR2_X1    g491(.A1(G106), .A2(G2105), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n917), .B(G2104), .C1(G118), .C2(new_n484), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n721), .A2(new_n919), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n717), .A2(new_n719), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n921), .A2(new_n922), .A3(new_n716), .A4(new_n720), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n920), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n924), .B1(new_n920), .B2(new_n923), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n914), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n920), .A2(new_n923), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT108), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n920), .A2(new_n923), .A3(new_n924), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(new_n647), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n913), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT109), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n908), .A2(new_n912), .A3(new_n927), .A4(new_n931), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n494), .A2(new_n495), .A3(new_n508), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n508), .B1(new_n494), .B2(new_n495), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n643), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(G160), .A2(G162), .ZN(new_n940));
  INV_X1    g515(.A(new_n643), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n494), .A2(new_n495), .A3(new_n508), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n913), .A2(new_n932), .A3(KEYINPUT109), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n936), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AOI22_X1  g521(.A1(new_n912), .A2(new_n908), .B1(new_n927), .B2(new_n931), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n947), .A2(new_n944), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT110), .B1(new_n948), .B2(new_n935), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n939), .A2(new_n943), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n950), .A2(new_n933), .A3(KEYINPUT110), .A4(new_n935), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n894), .B(new_n946), .C1(new_n949), .C2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT111), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n950), .A2(new_n933), .A3(new_n935), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(G37), .B1(new_n957), .B2(new_n951), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT111), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n959), .A3(new_n946), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n954), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT40), .ZN(G395));
  AOI22_X1  g537(.A1(new_n565), .A2(G87), .B1(G49), .B2(new_n549), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n963), .A2(new_n545), .A3(new_n596), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n545), .B1(new_n963), .B2(new_n596), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n729), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n966), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n968), .A2(new_n964), .A3(G290), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(G305), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n967), .A2(new_n969), .A3(new_n735), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n887), .B(new_n635), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n626), .B(new_n593), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT113), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n627), .A2(new_n593), .ZN(new_n979));
  NAND2_X1  g554(.A1(G299), .A2(new_n626), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT41), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(KEYINPUT112), .B(KEYINPUT41), .Z(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n982), .B1(new_n976), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n975), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n978), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n975), .A2(KEYINPUT113), .A3(new_n985), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n988), .B1(new_n987), .B2(new_n989), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n974), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n987), .A2(new_n989), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT42), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n994), .A2(new_n973), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(G868), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n877), .A2(new_n879), .A3(new_n880), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(G868), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n998), .A2(new_n1001), .ZN(G295));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n998), .A2(new_n1003), .A3(new_n1001), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n614), .B1(new_n992), .B2(new_n996), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT114), .B1(new_n1005), .B2(new_n1000), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(G331));
  XNOR2_X1  g582(.A(G301), .B(G286), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n884), .A2(new_n886), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1008), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n999), .B1(new_n574), .B2(new_n570), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(new_n885), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n985), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1009), .A2(new_n1012), .A3(new_n976), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n973), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n894), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n973), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT43), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT41), .B1(new_n979), .B2(new_n980), .ZN(new_n1020));
  AOI221_X4 g595(.A(new_n1020), .B1(new_n976), .B2(new_n983), .C1(new_n1009), .C2(new_n1012), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1015), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n974), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT43), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1023), .A2(new_n1024), .A3(new_n894), .A4(new_n1016), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1019), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1017), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1027), .A2(KEYINPUT43), .A3(new_n1023), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1024), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  MUX2_X1   g605(.A(new_n1026), .B(new_n1030), .S(KEYINPUT44), .Z(G397));
  INV_X1    g606(.A(KEYINPUT45), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(new_n901), .B2(G1384), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n477), .A2(new_n485), .A3(G40), .A4(new_n491), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n832), .B(new_n836), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1036), .B1(new_n792), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1996), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1035), .A2(KEYINPUT46), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT46), .B1(new_n1035), .B2(new_n1039), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1038), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n1042), .B(KEYINPUT47), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n791), .B(new_n1039), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1037), .A2(new_n726), .A3(new_n722), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n833), .A2(new_n836), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1036), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1035), .A2(new_n731), .A3(new_n729), .ZN(new_n1048));
  XOR2_X1   g623(.A(new_n1048), .B(KEYINPUT48), .Z(new_n1049));
  XNOR2_X1  g624(.A(new_n721), .B(new_n726), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1050), .B(KEYINPUT115), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1037), .A2(new_n1044), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1049), .B1(new_n1035), .B2(new_n1054), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1043), .A2(new_n1047), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G8), .ZN(new_n1057));
  INV_X1    g632(.A(G1384), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n513), .B2(new_n520), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(KEYINPUT50), .B(new_n1058), .C1(new_n513), .C2(new_n520), .ZN(new_n1062));
  AOI211_X1 g637(.A(G2090), .B(new_n1034), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g638(.A(KEYINPUT45), .B(new_n1058), .C1(new_n899), .C2(new_n900), .ZN(new_n1064));
  INV_X1    g639(.A(new_n512), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(new_n475), .B2(G126), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n519), .B(new_n515), .C1(new_n1066), .C2(new_n484), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT45), .B1(new_n1067), .B2(new_n1058), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1068), .A2(new_n1034), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1064), .A2(new_n1069), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1063), .A2(KEYINPUT116), .B1(new_n1070), .B2(new_n746), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1072));
  INV_X1    g647(.A(G2090), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1034), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1057), .B1(new_n1071), .B2(new_n1077), .ZN(new_n1078));
  AND2_X1   g653(.A1(KEYINPUT117), .A2(KEYINPUT55), .ZN(new_n1079));
  NOR2_X1   g654(.A1(KEYINPUT117), .A2(KEYINPUT55), .ZN(new_n1080));
  AOI211_X1 g655(.A(new_n1079), .B(new_n1080), .C1(G303), .C2(G8), .ZN(new_n1081));
  AND2_X1   g656(.A1(G303), .A2(G8), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1082), .B2(new_n1080), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1078), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1070), .A2(new_n746), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1057), .B1(new_n1085), .B2(new_n1075), .ZN(new_n1086));
  OR2_X1    g661(.A1(new_n1086), .A2(new_n1083), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT49), .ZN(new_n1088));
  NAND2_X1  g663(.A1(G305), .A2(G1981), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(G305), .A2(G1981), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1088), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OR2_X1    g667(.A1(G305), .A2(G1981), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1093), .A2(KEYINPUT49), .A3(new_n1089), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1059), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1074), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1092), .A2(new_n1094), .A3(G8), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G1976), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT52), .B1(G288), .B2(new_n1099), .ZN(new_n1100));
  XOR2_X1   g675(.A(new_n1100), .B(KEYINPUT119), .Z(new_n1101));
  OAI221_X1 g676(.A(G8), .B1(new_n1099), .B2(G288), .C1(new_n1034), .C2(new_n1059), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT52), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OR3_X1    g680(.A1(new_n1101), .A2(new_n1102), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1103), .A2(KEYINPUT52), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1102), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1098), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1059), .A2(new_n1032), .ZN(new_n1110));
  OAI211_X1 g685(.A(KEYINPUT45), .B(new_n1058), .C1(new_n513), .C2(new_n520), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1074), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1034), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1112), .A2(new_n813), .B1(new_n1113), .B2(new_n866), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1114), .A2(new_n1057), .A3(G286), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1084), .A2(new_n1087), .A3(new_n1109), .A4(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT63), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1109), .B(new_n1119), .C1(new_n1078), .C2(new_n1083), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1113), .A2(KEYINPUT116), .A3(new_n1073), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1085), .A2(new_n1077), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1083), .B1(new_n1122), .B2(G8), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1101), .A2(new_n1102), .A3(new_n1105), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1108), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1097), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT120), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1120), .A2(new_n1127), .A3(KEYINPUT63), .A4(new_n1084), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1115), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1118), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1084), .A2(new_n1126), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1096), .A2(G8), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1097), .A2(new_n1099), .A3(new_n596), .A4(new_n963), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1132), .B1(new_n1133), .B2(new_n1093), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1130), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(G286), .A2(G8), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT51), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1137), .B(new_n1140), .C1(new_n1114), .C2(new_n1057), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT50), .B1(new_n1067), .B2(new_n1058), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1062), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1074), .B(new_n866), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1111), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1145), .A2(new_n1068), .A3(new_n1034), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1144), .B1(new_n1146), .B2(G1966), .ZN(new_n1147));
  OAI211_X1 g722(.A(G8), .B(new_n1139), .C1(new_n1147), .C2(G286), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1147), .A2(G8), .A3(G286), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1141), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1141), .A2(new_n1148), .A3(KEYINPUT126), .A4(new_n1149), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT62), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n1070), .A2(G2078), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT53), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1156), .A2(new_n1157), .B1(new_n810), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1157), .A2(G2078), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1146), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1152), .A2(new_n1163), .A3(new_n1153), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1155), .A2(G171), .A3(new_n1162), .A4(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n593), .B(KEYINPUT57), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1158), .A2(new_n855), .ZN(new_n1167));
  XOR2_X1   g742(.A(KEYINPUT121), .B(G2072), .Z(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT56), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1064), .A2(new_n1069), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1167), .A2(KEYINPUT122), .A3(new_n1170), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1166), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1167), .A2(new_n1166), .A3(new_n1170), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1074), .A2(new_n836), .A3(new_n1095), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1177), .B1(new_n1113), .B2(G1348), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1175), .B1(new_n627), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1064), .A2(new_n1069), .A3(new_n1039), .ZN(new_n1181));
  XOR2_X1   g756(.A(KEYINPUT58), .B(G1341), .Z(new_n1182));
  NAND2_X1  g757(.A1(new_n1096), .A2(new_n1182), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1181), .A2(new_n1183), .A3(KEYINPUT123), .ZN(new_n1184));
  AOI21_X1  g759(.A(KEYINPUT123), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n575), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT59), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT60), .ZN(new_n1189));
  AOI21_X1  g764(.A(G1348), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n1034), .A2(G2067), .A3(new_n1059), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1189), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  OAI211_X1 g767(.A(new_n1177), .B(KEYINPUT60), .C1(new_n1113), .C2(G1348), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1192), .A2(new_n627), .A3(new_n1193), .ZN(new_n1194));
  OR2_X1    g769(.A1(new_n1193), .A2(new_n627), .ZN(new_n1195));
  AND2_X1   g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OAI211_X1 g771(.A(KEYINPUT59), .B(new_n575), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1188), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  OR2_X1    g773(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1176), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT61), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1167), .A2(new_n1201), .A3(new_n1170), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1166), .A2(new_n1201), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1200), .A2(new_n1204), .ZN(new_n1205));
  NAND4_X1  g780(.A1(new_n1176), .A2(new_n1202), .A3(new_n1203), .A4(new_n1199), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1180), .B1(new_n1198), .B2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(G301), .B(KEYINPUT54), .ZN(new_n1209));
  AOI22_X1  g784(.A1(new_n1152), .A2(new_n1153), .B1(new_n1209), .B2(new_n1162), .ZN(new_n1210));
  INV_X1    g785(.A(new_n1209), .ZN(new_n1211));
  NAND4_X1  g786(.A1(new_n1033), .A2(new_n1160), .A3(new_n1074), .A4(new_n1064), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1159), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1208), .A2(new_n1210), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1165), .A2(new_n1214), .ZN(new_n1215));
  AND3_X1   g790(.A1(new_n1084), .A2(new_n1087), .A3(new_n1109), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1136), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g792(.A(G290), .B(new_n731), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1036), .B1(new_n1053), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1056), .B1(new_n1217), .B2(new_n1219), .ZN(G329));
  assign    G231 = 1'b0;
  AOI211_X1 g795(.A(new_n460), .B(G229), .C1(new_n1019), .C2(new_n1025), .ZN(new_n1222));
  NAND3_X1  g796(.A1(new_n664), .A2(new_n681), .A3(new_n680), .ZN(new_n1223));
  INV_X1    g797(.A(new_n1223), .ZN(new_n1224));
  NOR2_X1   g798(.A1(new_n953), .A2(KEYINPUT111), .ZN(new_n1225));
  AOI21_X1  g799(.A(new_n959), .B1(new_n958), .B2(new_n946), .ZN(new_n1226));
  OAI211_X1 g800(.A(new_n1222), .B(new_n1224), .C1(new_n1225), .C2(new_n1226), .ZN(new_n1227));
  INV_X1    g801(.A(KEYINPUT127), .ZN(new_n1228));
  NOR2_X1   g802(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g803(.A(new_n1223), .B1(new_n954), .B2(new_n960), .ZN(new_n1230));
  AOI21_X1  g804(.A(KEYINPUT127), .B1(new_n1230), .B2(new_n1222), .ZN(new_n1231));
  NOR2_X1   g805(.A1(new_n1229), .A2(new_n1231), .ZN(G308));
  NAND2_X1  g806(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1233));
  NAND3_X1  g807(.A1(new_n1230), .A2(KEYINPUT127), .A3(new_n1222), .ZN(new_n1234));
  NAND2_X1  g808(.A1(new_n1233), .A2(new_n1234), .ZN(G225));
endmodule


