

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U322 ( .A(KEYINPUT78), .B(n550), .ZN(n467) );
  XNOR2_X1 U323 ( .A(n328), .B(n327), .ZN(n550) );
  XOR2_X1 U324 ( .A(n326), .B(n325), .Z(n327) );
  XNOR2_X1 U325 ( .A(n408), .B(KEYINPUT118), .ZN(n409) );
  NOR2_X2 U326 ( .A1(n447), .A2(n527), .ZN(n558) );
  INV_X1 U327 ( .A(KEYINPUT32), .ZN(n357) );
  XNOR2_X1 U328 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U329 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U330 ( .A(n360), .B(n359), .ZN(n362) );
  XNOR2_X1 U331 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U332 ( .A(n451), .B(n450), .ZN(G1351GAT) );
  XOR2_X1 U333 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n291) );
  XNOR2_X1 U334 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n290) );
  XNOR2_X1 U335 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U336 ( .A(G141GAT), .B(n292), .Z(n417) );
  XNOR2_X1 U337 ( .A(G134GAT), .B(G120GAT), .ZN(n293) );
  XNOR2_X1 U338 ( .A(n293), .B(KEYINPUT0), .ZN(n432) );
  XOR2_X1 U339 ( .A(G162GAT), .B(n432), .Z(n295) );
  XOR2_X1 U340 ( .A(G113GAT), .B(G1GAT), .Z(n368) );
  XNOR2_X1 U341 ( .A(G29GAT), .B(n368), .ZN(n294) );
  XNOR2_X1 U342 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U343 ( .A(n417), .B(n296), .ZN(n309) );
  XOR2_X1 U344 ( .A(G85GAT), .B(G155GAT), .Z(n298) );
  XNOR2_X1 U345 ( .A(G127GAT), .B(G148GAT), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U347 ( .A(KEYINPUT1), .B(G57GAT), .Z(n300) );
  XNOR2_X1 U348 ( .A(KEYINPUT94), .B(KEYINPUT6), .ZN(n299) );
  XNOR2_X1 U349 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U350 ( .A(n302), .B(n301), .Z(n307) );
  XOR2_X1 U351 ( .A(KEYINPUT93), .B(KEYINPUT4), .Z(n304) );
  NAND2_X1 U352 ( .A1(G225GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U354 ( .A(KEYINPUT5), .B(n305), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n513) );
  XOR2_X1 U357 ( .A(KEYINPUT76), .B(KEYINPUT74), .Z(n311) );
  XNOR2_X1 U358 ( .A(G134GAT), .B(KEYINPUT65), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n328) );
  XOR2_X1 U360 ( .A(G50GAT), .B(G162GAT), .Z(n413) );
  XOR2_X1 U361 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n313) );
  XNOR2_X1 U362 ( .A(KEYINPUT11), .B(KEYINPUT75), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n413), .B(n314), .ZN(n316) );
  AND2_X1 U365 ( .A1(G232GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U367 ( .A(KEYINPUT71), .B(G92GAT), .Z(n318) );
  XNOR2_X1 U368 ( .A(G99GAT), .B(G85GAT), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U370 ( .A(G106GAT), .B(n319), .ZN(n361) );
  XNOR2_X1 U371 ( .A(n320), .B(n361), .ZN(n326) );
  XOR2_X1 U372 ( .A(G29GAT), .B(G43GAT), .Z(n322) );
  XNOR2_X1 U373 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n367) );
  XOR2_X1 U375 ( .A(KEYINPUT77), .B(G218GAT), .Z(n324) );
  XNOR2_X1 U376 ( .A(G36GAT), .B(G190GAT), .ZN(n323) );
  XNOR2_X1 U377 ( .A(n324), .B(n323), .ZN(n399) );
  XNOR2_X1 U378 ( .A(n367), .B(n399), .ZN(n325) );
  XNOR2_X1 U379 ( .A(KEYINPUT36), .B(n467), .ZN(n483) );
  XOR2_X1 U380 ( .A(KEYINPUT81), .B(KEYINPUT83), .Z(n330) );
  XNOR2_X1 U381 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n329) );
  XNOR2_X1 U382 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U383 ( .A(G22GAT), .B(G155GAT), .Z(n421) );
  XOR2_X1 U384 ( .A(n421), .B(G78GAT), .Z(n332) );
  XOR2_X1 U385 ( .A(G15GAT), .B(G127GAT), .Z(n433) );
  XNOR2_X1 U386 ( .A(G1GAT), .B(n433), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U388 ( .A(n334), .B(n333), .Z(n336) );
  NAND2_X1 U389 ( .A1(G231GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U390 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U391 ( .A(KEYINPUT80), .B(KEYINPUT15), .Z(n338) );
  XNOR2_X1 U392 ( .A(G64GAT), .B(KEYINPUT82), .ZN(n337) );
  XNOR2_X1 U393 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U394 ( .A(n340), .B(n339), .Z(n346) );
  XOR2_X1 U395 ( .A(KEYINPUT79), .B(G211GAT), .Z(n342) );
  XNOR2_X1 U396 ( .A(G8GAT), .B(G183GAT), .ZN(n341) );
  XNOR2_X1 U397 ( .A(n342), .B(n341), .ZN(n391) );
  XOR2_X1 U398 ( .A(KEYINPUT69), .B(KEYINPUT13), .Z(n344) );
  XNOR2_X1 U399 ( .A(G71GAT), .B(G57GAT), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n344), .B(n343), .ZN(n354) );
  XNOR2_X1 U401 ( .A(n391), .B(n354), .ZN(n345) );
  XOR2_X1 U402 ( .A(n346), .B(n345), .Z(n468) );
  INV_X1 U403 ( .A(n468), .ZN(n576) );
  NAND2_X1 U404 ( .A1(n483), .A2(n576), .ZN(n347) );
  XNOR2_X1 U405 ( .A(n347), .B(KEYINPUT45), .ZN(n348) );
  XNOR2_X1 U406 ( .A(n348), .B(KEYINPUT64), .ZN(n363) );
  XOR2_X1 U407 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n350) );
  NAND2_X1 U408 ( .A1(G230GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U409 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U410 ( .A(n351), .B(KEYINPUT31), .Z(n356) );
  XOR2_X1 U411 ( .A(G78GAT), .B(G148GAT), .Z(n353) );
  XNOR2_X1 U412 ( .A(KEYINPUT70), .B(G204GAT), .ZN(n352) );
  XNOR2_X1 U413 ( .A(n353), .B(n352), .ZN(n425) );
  XNOR2_X1 U414 ( .A(n425), .B(n354), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U416 ( .A(G176GAT), .B(G64GAT), .Z(n390) );
  XNOR2_X1 U417 ( .A(G120GAT), .B(n390), .ZN(n358) );
  XOR2_X1 U418 ( .A(n362), .B(n361), .Z(n571) );
  NOR2_X1 U419 ( .A1(n363), .A2(n571), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n364), .B(KEYINPUT112), .ZN(n382) );
  XOR2_X1 U421 ( .A(G22GAT), .B(G141GAT), .Z(n366) );
  XNOR2_X1 U422 ( .A(G169GAT), .B(G15GAT), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n381) );
  XOR2_X1 U424 ( .A(n368), .B(n367), .Z(n370) );
  XNOR2_X1 U425 ( .A(G50GAT), .B(G36GAT), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U427 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n372) );
  NAND2_X1 U428 ( .A1(G229GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U429 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U430 ( .A(n374), .B(n373), .Z(n379) );
  XOR2_X1 U431 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n376) );
  XNOR2_X1 U432 ( .A(G197GAT), .B(G8GAT), .ZN(n375) );
  XNOR2_X1 U433 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n377), .B(KEYINPUT66), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U436 ( .A(n381), .B(n380), .ZN(n499) );
  NAND2_X1 U437 ( .A1(n382), .A2(n499), .ZN(n388) );
  INV_X1 U438 ( .A(n499), .ZN(n568) );
  XOR2_X1 U439 ( .A(n571), .B(KEYINPUT41), .Z(n544) );
  NAND2_X1 U440 ( .A1(n568), .A2(n544), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n383), .B(KEYINPUT46), .ZN(n384) );
  XOR2_X1 U442 ( .A(n468), .B(KEYINPUT111), .Z(n560) );
  NAND2_X1 U443 ( .A1(n384), .A2(n560), .ZN(n385) );
  NOR2_X1 U444 ( .A1(n550), .A2(n385), .ZN(n386) );
  XNOR2_X1 U445 ( .A(KEYINPUT47), .B(n386), .ZN(n387) );
  NAND2_X1 U446 ( .A1(n388), .A2(n387), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n389), .B(KEYINPUT48), .ZN(n524) );
  XOR2_X1 U448 ( .A(n391), .B(n390), .Z(n393) );
  XNOR2_X1 U449 ( .A(G204GAT), .B(G92GAT), .ZN(n392) );
  XNOR2_X1 U450 ( .A(n393), .B(n392), .ZN(n403) );
  XOR2_X1 U451 ( .A(KEYINPUT95), .B(KEYINPUT97), .Z(n395) );
  NAND2_X1 U452 ( .A1(G226GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U453 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U454 ( .A(n396), .B(KEYINPUT96), .Z(n401) );
  XOR2_X1 U455 ( .A(KEYINPUT88), .B(KEYINPUT21), .Z(n398) );
  XNOR2_X1 U456 ( .A(G197GAT), .B(KEYINPUT87), .ZN(n397) );
  XNOR2_X1 U457 ( .A(n398), .B(n397), .ZN(n412) );
  XNOR2_X1 U458 ( .A(n412), .B(n399), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U460 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U461 ( .A(KEYINPUT85), .B(KEYINPUT17), .Z(n405) );
  XNOR2_X1 U462 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U464 ( .A(G169GAT), .B(n406), .Z(n446) );
  XOR2_X1 U465 ( .A(n407), .B(n446), .Z(n516) );
  AND2_X1 U466 ( .A1(n524), .A2(n516), .ZN(n410) );
  XNOR2_X1 U467 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n408) );
  NOR2_X1 U468 ( .A1(n513), .A2(n411), .ZN(n565) );
  XOR2_X1 U469 ( .A(n413), .B(n412), .Z(n415) );
  NAND2_X1 U470 ( .A1(G228GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n417), .B(n416), .ZN(n429) );
  XOR2_X1 U473 ( .A(G211GAT), .B(KEYINPUT23), .Z(n419) );
  XNOR2_X1 U474 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U476 ( .A(n420), .B(G106GAT), .Z(n423) );
  XNOR2_X1 U477 ( .A(n421), .B(G218GAT), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U479 ( .A(n424), .B(KEYINPUT91), .Z(n427) );
  XNOR2_X1 U480 ( .A(n425), .B(KEYINPUT92), .ZN(n426) );
  XNOR2_X1 U481 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n429), .B(n428), .ZN(n462) );
  NAND2_X1 U483 ( .A1(n565), .A2(n462), .ZN(n431) );
  XOR2_X1 U484 ( .A(KEYINPUT120), .B(KEYINPUT55), .Z(n430) );
  XNOR2_X1 U485 ( .A(n431), .B(n430), .ZN(n447) );
  XOR2_X1 U486 ( .A(n433), .B(n432), .Z(n435) );
  XNOR2_X1 U487 ( .A(G43GAT), .B(G190GAT), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U489 ( .A(KEYINPUT86), .B(G183GAT), .Z(n437) );
  NAND2_X1 U490 ( .A1(G227GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U492 ( .A(n439), .B(n438), .Z(n444) );
  XOR2_X1 U493 ( .A(KEYINPUT20), .B(G71GAT), .Z(n441) );
  XNOR2_X1 U494 ( .A(G99GAT), .B(G176GAT), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U496 ( .A(G113GAT), .B(n442), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U498 ( .A(n446), .B(n445), .ZN(n527) );
  NAND2_X1 U499 ( .A1(n558), .A2(n467), .ZN(n451) );
  XOR2_X1 U500 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n449) );
  INV_X1 U501 ( .A(G190GAT), .ZN(n448) );
  INV_X1 U502 ( .A(KEYINPUT100), .ZN(n458) );
  INV_X1 U503 ( .A(n527), .ZN(n518) );
  NAND2_X1 U504 ( .A1(n518), .A2(n516), .ZN(n452) );
  NAND2_X1 U505 ( .A1(n462), .A2(n452), .ZN(n453) );
  XOR2_X1 U506 ( .A(KEYINPUT25), .B(n453), .Z(n456) );
  XNOR2_X1 U507 ( .A(KEYINPUT27), .B(n516), .ZN(n460) );
  NOR2_X1 U508 ( .A1(n462), .A2(n518), .ZN(n454) );
  XNOR2_X1 U509 ( .A(n454), .B(KEYINPUT26), .ZN(n566) );
  NAND2_X1 U510 ( .A1(n460), .A2(n566), .ZN(n455) );
  NAND2_X1 U511 ( .A1(n456), .A2(n455), .ZN(n457) );
  XNOR2_X1 U512 ( .A(n458), .B(n457), .ZN(n459) );
  NOR2_X1 U513 ( .A1(n513), .A2(n459), .ZN(n465) );
  NAND2_X1 U514 ( .A1(n460), .A2(n513), .ZN(n461) );
  XNOR2_X1 U515 ( .A(n461), .B(KEYINPUT98), .ZN(n541) );
  XOR2_X1 U516 ( .A(n462), .B(KEYINPUT28), .Z(n520) );
  NOR2_X1 U517 ( .A1(n541), .A2(n520), .ZN(n525) );
  XNOR2_X1 U518 ( .A(KEYINPUT99), .B(n525), .ZN(n463) );
  NOR2_X1 U519 ( .A1(n518), .A2(n463), .ZN(n464) );
  NOR2_X1 U520 ( .A1(n465), .A2(n464), .ZN(n466) );
  XOR2_X1 U521 ( .A(KEYINPUT101), .B(n466), .Z(n484) );
  XOR2_X1 U522 ( .A(KEYINPUT84), .B(KEYINPUT16), .Z(n470) );
  NOR2_X1 U523 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U524 ( .A(n470), .B(n469), .ZN(n471) );
  NOR2_X1 U525 ( .A1(n484), .A2(n471), .ZN(n498) );
  OR2_X1 U526 ( .A1(n571), .A2(n499), .ZN(n472) );
  XNOR2_X1 U527 ( .A(n472), .B(KEYINPUT73), .ZN(n487) );
  NAND2_X1 U528 ( .A1(n498), .A2(n487), .ZN(n473) );
  XOR2_X1 U529 ( .A(KEYINPUT102), .B(n473), .Z(n481) );
  NAND2_X1 U530 ( .A1(n481), .A2(n513), .ZN(n474) );
  XNOR2_X1 U531 ( .A(n474), .B(KEYINPUT34), .ZN(n475) );
  XNOR2_X1 U532 ( .A(G1GAT), .B(n475), .ZN(G1324GAT) );
  XOR2_X1 U533 ( .A(G8GAT), .B(KEYINPUT103), .Z(n477) );
  NAND2_X1 U534 ( .A1(n481), .A2(n516), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n477), .B(n476), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n479) );
  NAND2_X1 U537 ( .A1(n518), .A2(n481), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U539 ( .A(G15GAT), .B(n480), .ZN(G1326GAT) );
  NAND2_X1 U540 ( .A1(n481), .A2(n520), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT106), .B(KEYINPUT39), .Z(n491) );
  XOR2_X1 U543 ( .A(KEYINPUT38), .B(KEYINPUT105), .Z(n489) );
  NOR2_X1 U544 ( .A1(n576), .A2(n484), .ZN(n485) );
  NAND2_X1 U545 ( .A1(n483), .A2(n485), .ZN(n486) );
  XNOR2_X1 U546 ( .A(KEYINPUT37), .B(n486), .ZN(n510) );
  NAND2_X1 U547 ( .A1(n487), .A2(n510), .ZN(n488) );
  XOR2_X1 U548 ( .A(n489), .B(n488), .Z(n496) );
  NAND2_X1 U549 ( .A1(n513), .A2(n496), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U551 ( .A(G29GAT), .B(n492), .ZN(G1328GAT) );
  NAND2_X1 U552 ( .A1(n496), .A2(n516), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n493), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U554 ( .A1(n496), .A2(n518), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n494), .B(KEYINPUT40), .ZN(n495) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  NAND2_X1 U557 ( .A1(n496), .A2(n520), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n497), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U559 ( .A(n498), .ZN(n500) );
  XOR2_X1 U560 ( .A(KEYINPUT107), .B(n544), .Z(n554) );
  NAND2_X1 U561 ( .A1(n499), .A2(n554), .ZN(n511) );
  NOR2_X1 U562 ( .A1(n500), .A2(n511), .ZN(n506) );
  NAND2_X1 U563 ( .A1(n513), .A2(n506), .ZN(n501) );
  XNOR2_X1 U564 ( .A(KEYINPUT42), .B(n501), .ZN(n502) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(n502), .ZN(G1332GAT) );
  NAND2_X1 U566 ( .A1(n516), .A2(n506), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n503), .B(KEYINPUT108), .ZN(n504) );
  XNOR2_X1 U568 ( .A(G64GAT), .B(n504), .ZN(G1333GAT) );
  NAND2_X1 U569 ( .A1(n506), .A2(n518), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n505), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n508) );
  NAND2_X1 U572 ( .A1(n506), .A2(n520), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U574 ( .A(G78GAT), .B(n509), .Z(G1335GAT) );
  XNOR2_X1 U575 ( .A(G85GAT), .B(KEYINPUT110), .ZN(n515) );
  INV_X1 U576 ( .A(n510), .ZN(n512) );
  NOR2_X1 U577 ( .A1(n512), .A2(n511), .ZN(n521) );
  NAND2_X1 U578 ( .A1(n513), .A2(n521), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(G1336GAT) );
  NAND2_X1 U580 ( .A1(n516), .A2(n521), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n517), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U582 ( .A1(n521), .A2(n518), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n519), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U584 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U585 ( .A(n522), .B(KEYINPUT44), .ZN(n523) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  XOR2_X1 U587 ( .A(G113GAT), .B(KEYINPUT113), .Z(n529) );
  NAND2_X1 U588 ( .A1(n524), .A2(n525), .ZN(n526) );
  NOR2_X1 U589 ( .A1(n527), .A2(n526), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n536), .A2(n568), .ZN(n528) );
  XNOR2_X1 U591 ( .A(n529), .B(n528), .ZN(G1340GAT) );
  XOR2_X1 U592 ( .A(G120GAT), .B(KEYINPUT49), .Z(n531) );
  NAND2_X1 U593 ( .A1(n536), .A2(n554), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  INV_X1 U595 ( .A(n536), .ZN(n532) );
  NOR2_X1 U596 ( .A1(n560), .A2(n532), .ZN(n534) );
  XNOR2_X1 U597 ( .A(KEYINPUT50), .B(KEYINPUT114), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U599 ( .A(G127GAT), .B(n535), .Z(G1342GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT51), .B(KEYINPUT115), .Z(n538) );
  NAND2_X1 U601 ( .A1(n536), .A2(n467), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U603 ( .A(G134GAT), .B(n539), .Z(G1343GAT) );
  NAND2_X1 U604 ( .A1(n524), .A2(n566), .ZN(n540) );
  NOR2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n551), .A2(n568), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n542), .B(KEYINPUT116), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(n543), .ZN(G1344GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT117), .B(KEYINPUT53), .Z(n546) );
  NAND2_X1 U610 ( .A1(n551), .A2(n544), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT52), .Z(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NAND2_X1 U614 ( .A1(n551), .A2(n576), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n549), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n552), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U618 ( .A1(n558), .A2(n568), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U620 ( .A1(n558), .A2(n554), .ZN(n556) );
  XOR2_X1 U621 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(G176GAT), .ZN(G1349GAT) );
  INV_X1 U624 ( .A(n558), .ZN(n559) );
  NOR2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n562) );
  XNOR2_X1 U626 ( .A(G183GAT), .B(KEYINPUT121), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1350GAT) );
  XNOR2_X1 U628 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT124), .ZN(n564) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(n564), .Z(n570) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n567), .B(KEYINPUT123), .ZN(n578) );
  NAND2_X1 U633 ( .A1(n578), .A2(n568), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n573) );
  NAND2_X1 U636 ( .A1(n578), .A2(n571), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n573), .B(n572), .ZN(n575) );
  XOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT125), .Z(n574) );
  XNOR2_X1 U639 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  NAND2_X1 U640 ( .A1(n578), .A2(n576), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n580) );
  NAND2_X1 U643 ( .A1(n578), .A2(n483), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

