//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n816, new_n817, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934;
  INV_X1    g000(.A(KEYINPUT14), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  AOI22_X1  g005(.A1(new_n205), .A2(new_n206), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(G43gat), .B(G50gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(KEYINPUT15), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT17), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(KEYINPUT91), .ZN(new_n213));
  XNOR2_X1  g012(.A(G15gat), .B(G22gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT16), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n214), .B1(new_n215), .B2(G1gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT90), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n216), .B(new_n217), .C1(G1gat), .C2(new_n214), .ZN(new_n218));
  INV_X1    g017(.A(G8gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT89), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(new_n211), .B2(KEYINPUT17), .ZN(new_n222));
  OR3_X1    g021(.A1(new_n211), .A2(new_n221), .A3(KEYINPUT17), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n213), .A2(new_n220), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G229gat), .A2(G233gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n220), .A2(new_n211), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT92), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n224), .A2(KEYINPUT18), .A3(new_n225), .A4(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n220), .A2(new_n211), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n225), .B(KEYINPUT13), .Z(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G113gat), .B(G141gat), .ZN(new_n235));
  INV_X1    g034(.A(G197gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT11), .B(G169gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT12), .Z(new_n240));
  NOR2_X1   g039(.A1(new_n234), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n224), .A2(new_n225), .A3(new_n228), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT93), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT18), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n242), .A2(new_n244), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT93), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n241), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n246), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n240), .B1(new_n249), .B2(new_n234), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT21), .ZN(new_n252));
  XNOR2_X1  g051(.A(G57gat), .B(G64gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT9), .ZN(new_n254));
  INV_X1    g053(.A(G71gat), .ZN(new_n255));
  INV_X1    g054(.A(G78gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n253), .B1(KEYINPUT94), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G71gat), .B(G78gat), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n258), .B(new_n259), .C1(KEYINPUT94), .C2(new_n257), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n253), .A2(new_n254), .ZN(new_n261));
  OR2_X1    g060(.A1(new_n261), .A2(new_n259), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n220), .B1(new_n252), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G183gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n266), .B(new_n267), .Z(new_n268));
  NAND2_X1  g067(.A1(new_n263), .A2(new_n252), .ZN(new_n269));
  INV_X1    g068(.A(G211gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n266), .B(new_n267), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(new_n271), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G127gat), .B(G155gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(G231gat), .A2(G233gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n273), .A2(new_n275), .A3(new_n279), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G134gat), .B(G162gat), .ZN(new_n284));
  XOR2_X1   g083(.A(G190gat), .B(G218gat), .Z(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT96), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n288));
  XOR2_X1   g087(.A(new_n287), .B(new_n288), .Z(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G99gat), .A2(G106gat), .ZN(new_n291));
  INV_X1    g090(.A(G85gat), .ZN(new_n292));
  INV_X1    g091(.A(G92gat), .ZN(new_n293));
  AOI22_X1  g092(.A1(KEYINPUT8), .A2(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(KEYINPUT95), .A2(G85gat), .A3(G92gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT7), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g096(.A1(KEYINPUT95), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n294), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  XOR2_X1   g098(.A(G99gat), .B(G106gat), .Z(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n213), .A2(new_n222), .A3(new_n223), .A4(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n211), .A2(new_n301), .ZN(new_n303));
  AND3_X1   g102(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n286), .A2(KEYINPUT96), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n290), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n306), .A2(new_n308), .A3(new_n290), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n284), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n311), .ZN(new_n313));
  INV_X1    g112(.A(new_n284), .ZN(new_n314));
  NOR3_X1   g113(.A1(new_n313), .A2(new_n314), .A3(new_n309), .ZN(new_n315));
  OR2_X1    g114(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n263), .A2(new_n301), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n263), .A2(new_n301), .ZN(new_n318));
  OR3_X1    g117(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT10), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(KEYINPUT10), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G230gat), .A2(G233gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n322), .B(KEYINPUT97), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n323), .B1(new_n317), .B2(new_n318), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT98), .B(G120gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(G148gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(G176gat), .B(G204gat), .ZN(new_n330));
  XOR2_X1   g129(.A(new_n329), .B(new_n330), .Z(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n325), .A2(new_n326), .A3(new_n331), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n283), .A2(new_n316), .A3(new_n336), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n337), .A2(KEYINPUT99), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(KEYINPUT99), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT85), .ZN(new_n341));
  XNOR2_X1  g140(.A(G211gat), .B(G218gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT22), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT74), .B(G211gat), .ZN(new_n345));
  INV_X1    g144(.A(G218gat), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n348));
  XNOR2_X1  g147(.A(G197gat), .B(G204gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n348), .B1(new_n347), .B2(new_n349), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n343), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n352), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(new_n350), .A3(new_n342), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n358));
  NAND2_X1  g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359));
  INV_X1    g158(.A(G155gat), .ZN(new_n360));
  INV_X1    g159(.A(G162gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G141gat), .B(G148gat), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n359), .B(new_n362), .C1(new_n363), .C2(KEYINPUT2), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT80), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n359), .B1(new_n362), .B2(KEYINPUT2), .ZN(new_n367));
  INV_X1    g166(.A(G141gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(G148gat), .ZN(new_n369));
  INV_X1    g168(.A(G148gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n370), .A2(G141gat), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n367), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT2), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(new_n369), .B2(new_n371), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n374), .A2(KEYINPUT80), .A3(new_n359), .A4(new_n362), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n366), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n357), .A2(new_n358), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(KEYINPUT3), .ZN(new_n378));
  NAND2_X1  g177(.A1(G228gat), .A2(G233gat), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n358), .B1(new_n376), .B2(KEYINPUT3), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n356), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n377), .A2(new_n378), .A3(new_n379), .A4(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n353), .A2(new_n355), .A3(new_n358), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT84), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT3), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n353), .A2(new_n355), .A3(KEYINPUT84), .A4(new_n358), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n388), .A2(new_n376), .B1(new_n380), .B2(new_n356), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n382), .B1(new_n389), .B2(new_n379), .ZN(new_n390));
  XNOR2_X1  g189(.A(G78gat), .B(G106gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(G22gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT31), .B(G50gat), .ZN(new_n394));
  INV_X1    g193(.A(new_n392), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n382), .B(new_n395), .C1(new_n389), .C2(new_n379), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n393), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n394), .B1(new_n393), .B2(new_n396), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G1gat), .B(G29gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(new_n292), .ZN(new_n401));
  XNOR2_X1  g200(.A(KEYINPUT0), .B(G57gat), .ZN(new_n402));
  XOR2_X1   g201(.A(new_n401), .B(new_n402), .Z(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G113gat), .B(G120gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(KEYINPUT1), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT69), .B(G134gat), .ZN(new_n409));
  INV_X1    g208(.A(G127gat), .ZN(new_n410));
  OR2_X1    g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(G134gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n412), .A2(G127gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n408), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  AND2_X1   g214(.A1(KEYINPUT70), .A2(G120gat), .ZN(new_n416));
  NOR2_X1   g215(.A1(KEYINPUT70), .A2(G120gat), .ZN(new_n417));
  OAI21_X1  g216(.A(G113gat), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT71), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT72), .ZN(new_n421));
  INV_X1    g220(.A(G113gat), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(G120gat), .ZN(new_n423));
  INV_X1    g222(.A(G120gat), .ZN(new_n424));
  NOR3_X1   g223(.A1(new_n424), .A2(KEYINPUT72), .A3(G113gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g225(.A(KEYINPUT71), .B(G113gat), .C1(new_n416), .C2(new_n417), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n420), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n410), .A2(G134gat), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n413), .A2(new_n429), .A3(KEYINPUT1), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT73), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n428), .A2(KEYINPUT73), .A3(new_n430), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n415), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n376), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI211_X1 g236(.A(new_n415), .B(new_n376), .C1(new_n433), .C2(new_n434), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n406), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT81), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(new_n440), .A3(KEYINPUT5), .ZN(new_n441));
  INV_X1    g240(.A(new_n415), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n428), .A2(KEYINPUT73), .A3(new_n430), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT73), .B1(new_n428), .B2(new_n430), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n376), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n436), .B(new_n442), .C1(new_n443), .C2(new_n444), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n405), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT5), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT81), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n447), .A2(KEYINPUT4), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT4), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n435), .A2(new_n452), .A3(new_n436), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n376), .A2(KEYINPUT3), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n435), .A2(new_n454), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n451), .A2(new_n453), .B1(new_n455), .B2(new_n378), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n441), .A2(new_n450), .B1(new_n405), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n451), .A2(new_n453), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n455), .A2(new_n378), .ZN(new_n459));
  AND4_X1   g258(.A1(KEYINPUT5), .A2(new_n458), .A3(new_n459), .A4(new_n405), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n404), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n456), .A2(new_n405), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n440), .B1(new_n439), .B2(KEYINPUT5), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n448), .A2(KEYINPUT81), .A3(new_n449), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n460), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n466), .A3(new_n403), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT6), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n461), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n465), .A2(KEYINPUT6), .A3(new_n466), .A4(new_n403), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT82), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n441), .A2(new_n450), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n460), .B1(new_n473), .B2(new_n462), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n474), .A2(KEYINPUT82), .A3(KEYINPUT6), .A4(new_n403), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n469), .A2(new_n472), .A3(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT77), .B(G64gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(G92gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(G8gat), .B(G36gat), .ZN(new_n479));
  XOR2_X1   g278(.A(new_n478), .B(new_n479), .Z(new_n480));
  AOI21_X1  g279(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n481), .B1(G169gat), .B2(G176gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(G183gat), .A2(G190gat), .ZN(new_n483));
  NOR2_X1   g282(.A1(G169gat), .A2(G176gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT26), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT68), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n482), .A2(KEYINPUT68), .A3(new_n483), .A4(new_n485), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT67), .ZN(new_n491));
  XOR2_X1   g290(.A(KEYINPUT27), .B(G183gat), .Z(new_n492));
  OAI211_X1 g291(.A(new_n491), .B(KEYINPUT28), .C1(new_n492), .C2(G190gat), .ZN(new_n493));
  INV_X1    g292(.A(new_n492), .ZN(new_n494));
  INV_X1    g293(.A(G190gat), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n491), .A2(KEYINPUT28), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n491), .A2(KEYINPUT28), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n494), .A2(new_n495), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n490), .A2(new_n493), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT25), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT24), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n265), .A2(new_n495), .A3(KEYINPUT64), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT64), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(G183gat), .B2(G190gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n506));
  AND4_X1   g305(.A1(new_n502), .A2(new_n503), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n484), .A2(KEYINPUT23), .ZN(new_n508));
  NAND2_X1  g307(.A1(G169gat), .A2(G176gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT23), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n510), .B1(G169gat), .B2(G176gat), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n500), .B1(new_n507), .B2(new_n512), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n501), .B1(new_n483), .B2(KEYINPUT65), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT65), .ZN(new_n516));
  OAI22_X1  g315(.A1(new_n502), .A2(new_n516), .B1(G183gat), .B2(G190gat), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n514), .B(KEYINPUT25), .C1(new_n515), .C2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(KEYINPUT66), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT66), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n521), .B1(new_n513), .B2(new_n518), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n499), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(G226gat), .A2(G233gat), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n524), .B(KEYINPUT76), .Z(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n523), .A2(new_n358), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n499), .A2(new_n519), .A3(new_n525), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n357), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n523), .A2(new_n525), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n499), .A2(new_n519), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(new_n358), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n526), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n356), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(KEYINPUT30), .B(new_n480), .C1(new_n529), .C2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n529), .A2(new_n534), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n480), .B(KEYINPUT78), .Z(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n480), .B1(new_n529), .B2(new_n534), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT79), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT79), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n542), .B(new_n480), .C1(new_n529), .C2(new_n534), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n545));
  AOI211_X1 g344(.A(new_n536), .B(new_n539), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n476), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT83), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT83), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n476), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n399), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT36), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n523), .A2(new_n445), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n435), .B(new_n499), .C1(new_n522), .C2(new_n520), .ZN(new_n554));
  NAND2_X1  g353(.A1(G227gat), .A2(G233gat), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT34), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT34), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n553), .A2(new_n554), .A3(new_n558), .A4(new_n555), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n555), .B1(new_n553), .B2(new_n554), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT32), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G15gat), .B(G43gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(G71gat), .B(G99gat), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n565), .B(new_n566), .Z(new_n567));
  OAI21_X1  g366(.A(new_n567), .B1(new_n561), .B2(KEYINPUT33), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n557), .B(new_n559), .C1(new_n562), .C2(new_n561), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n564), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n569), .B1(new_n564), .B2(new_n570), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n552), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n564), .A2(new_n570), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n568), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n576), .A2(KEYINPUT36), .A3(new_n571), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n341), .B1(new_n551), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n539), .B1(new_n544), .B2(new_n545), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n535), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n458), .A2(new_n459), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(new_n406), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT86), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n446), .A2(new_n405), .A3(new_n447), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n587), .B1(new_n583), .B2(new_n406), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT39), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n586), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n584), .A2(new_n585), .A3(KEYINPUT39), .A4(new_n587), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n590), .A2(new_n404), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT40), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n590), .A2(KEYINPUT40), .A3(new_n404), .A4(new_n591), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n582), .A2(new_n467), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n527), .A2(new_n528), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n357), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT87), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT87), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n597), .A2(new_n600), .A3(new_n357), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n530), .A2(new_n533), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n599), .B(new_n601), .C1(new_n357), .C2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT38), .B1(new_n603), .B2(KEYINPUT37), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT37), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n538), .B1(new_n537), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n607), .A2(new_n475), .A3(new_n472), .A4(new_n469), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n537), .A2(new_n605), .ZN(new_n609));
  INV_X1    g408(.A(new_n480), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n537), .A2(new_n605), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT38), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n544), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n596), .B(new_n399), .C1(new_n608), .C2(new_n614), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n397), .A2(new_n398), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n476), .A2(new_n546), .A3(new_n549), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n549), .B1(new_n476), .B2(new_n546), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n619), .A2(KEYINPUT85), .A3(new_n578), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n580), .A2(new_n615), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n576), .A2(new_n571), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n616), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n548), .A2(new_n623), .A3(new_n550), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT35), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT35), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT88), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n572), .A2(new_n573), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT88), .B1(new_n576), .B2(new_n571), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n399), .B(new_n626), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n630), .A2(new_n547), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n625), .A2(new_n632), .ZN(new_n633));
  AOI211_X1 g432(.A(new_n251), .B(new_n340), .C1(new_n621), .C2(new_n633), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n476), .A2(KEYINPUT100), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n476), .A2(KEYINPUT100), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g438(.A1(new_n634), .A2(new_n582), .ZN(new_n640));
  XOR2_X1   g439(.A(KEYINPUT16), .B(G8gat), .Z(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT42), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n640), .A2(KEYINPUT42), .A3(new_n641), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n644), .B(new_n645), .C1(new_n219), .C2(new_n640), .ZN(G1325gat));
  NOR2_X1   g445(.A1(new_n628), .A2(new_n629), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n634), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(G15gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n651), .A2(KEYINPUT101), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(KEYINPUT101), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n574), .A2(new_n577), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n654), .B1(new_n574), .B2(new_n577), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n657), .B(KEYINPUT103), .Z(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n659), .A2(new_n650), .ZN(new_n660));
  AOI22_X1  g459(.A1(new_n652), .A2(new_n653), .B1(new_n634), .B2(new_n660), .ZN(G1326gat));
  NAND2_X1  g460(.A1(new_n634), .A2(new_n616), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT43), .B(G22gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1327gat));
  AOI21_X1  g463(.A(new_n316), .B1(new_n621), .B2(new_n633), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n283), .A2(new_n251), .A3(new_n335), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n667), .A2(new_n203), .A3(new_n637), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT45), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n619), .A2(new_n615), .A3(new_n657), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n633), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n312), .A2(new_n315), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(new_n665), .B2(new_n672), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n666), .B(KEYINPUT104), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n637), .ZN(new_n679));
  OAI21_X1  g478(.A(G29gat), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n669), .A2(new_n680), .ZN(G1328gat));
  NAND3_X1  g480(.A1(new_n667), .A2(new_n204), .A3(new_n582), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT46), .Z(new_n683));
  OAI21_X1  g482(.A(G36gat), .B1(new_n678), .B2(new_n546), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(G1329gat));
  INV_X1    g484(.A(G43gat), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n665), .A2(new_n686), .A3(new_n648), .A4(new_n666), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT47), .ZN(new_n688));
  INV_X1    g487(.A(new_n657), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n675), .A2(new_n689), .A3(new_n677), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n688), .B1(new_n690), .B2(G43gat), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n691), .A2(KEYINPUT105), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(KEYINPUT105), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n675), .A2(new_n658), .A3(new_n677), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G43gat), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n695), .A2(new_n687), .ZN(new_n696));
  OAI22_X1  g495(.A1(new_n692), .A2(new_n693), .B1(new_n696), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g496(.A(G50gat), .B1(new_n678), .B2(new_n399), .ZN(new_n698));
  INV_X1    g497(.A(G50gat), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n667), .A2(new_n699), .A3(new_n616), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n698), .A2(KEYINPUT48), .A3(new_n700), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n698), .A2(KEYINPUT106), .A3(new_n700), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT48), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(new_n698), .B2(KEYINPUT106), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n701), .B1(new_n702), .B2(new_n704), .ZN(G1331gat));
  NAND3_X1  g504(.A1(new_n283), .A2(new_n316), .A3(new_n251), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n336), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT107), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n671), .A2(new_n708), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n709), .A2(KEYINPUT108), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(KEYINPUT108), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n637), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g514(.A1(new_n712), .A2(new_n546), .ZN(new_n716));
  NOR2_X1   g515(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n717));
  AND2_X1   g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n716), .B2(new_n717), .ZN(G1333gat));
  NAND3_X1  g519(.A1(new_n713), .A2(G71gat), .A3(new_n658), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n255), .B1(new_n712), .B2(new_n647), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT50), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT50), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n721), .A2(new_n725), .A3(new_n722), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(G1334gat));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n399), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(new_n256), .ZN(G1335gat));
  NAND2_X1  g528(.A1(new_n248), .A2(new_n250), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n283), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n675), .A2(new_n637), .A3(new_n335), .A4(new_n731), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n732), .A2(G85gat), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n619), .A2(new_n615), .A3(new_n657), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n631), .B1(new_n624), .B2(KEYINPUT35), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n673), .B(new_n731), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT51), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n671), .A2(KEYINPUT51), .A3(new_n673), .A4(new_n731), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n736), .A2(KEYINPUT109), .A3(new_n737), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n741), .A2(new_n637), .A3(new_n335), .A4(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(G85gat), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n733), .A2(new_n744), .A3(KEYINPUT110), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n741), .A2(new_n742), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n747), .A2(new_n292), .A3(new_n637), .A4(new_n335), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n732), .A2(G85gat), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n746), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n745), .A2(new_n750), .ZN(G1336gat));
  NOR2_X1   g550(.A1(new_n546), .A2(G92gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n747), .A2(new_n335), .A3(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n675), .A2(new_n335), .A3(new_n582), .A4(new_n731), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n756), .A2(G92gat), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n336), .B1(new_n738), .B2(new_n739), .ZN(new_n758));
  AOI22_X1  g557(.A1(new_n756), .A2(G92gat), .B1(new_n752), .B2(new_n758), .ZN(new_n759));
  OAI22_X1  g558(.A1(new_n755), .A2(new_n757), .B1(new_n754), .B2(new_n759), .ZN(G1337gat));
  NOR2_X1   g559(.A1(new_n647), .A2(G99gat), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n747), .A2(new_n335), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n675), .A2(new_n335), .A3(new_n731), .ZN(new_n763));
  OAI21_X1  g562(.A(G99gat), .B1(new_n763), .B2(new_n659), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(G1338gat));
  NOR3_X1   g564(.A1(new_n399), .A2(G106gat), .A3(new_n336), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n747), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n675), .A2(new_n335), .A3(new_n616), .A4(new_n731), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(G106gat), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n738), .A2(new_n739), .ZN(new_n772));
  AOI22_X1  g571(.A1(new_n770), .A2(G106gat), .B1(new_n772), .B2(new_n766), .ZN(new_n773));
  OAI22_X1  g572(.A1(new_n769), .A2(new_n771), .B1(new_n773), .B2(new_n768), .ZN(G1339gat));
  NOR2_X1   g573(.A1(new_n706), .A2(new_n335), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n231), .A2(new_n232), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n225), .B1(new_n224), .B2(new_n228), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n239), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n248), .A2(new_n335), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n319), .A2(new_n320), .A3(new_n323), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n325), .A2(KEYINPUT54), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n323), .B1(new_n319), .B2(new_n320), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n331), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n782), .A2(KEYINPUT55), .A3(new_n785), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n334), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n248), .B2(new_n250), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n316), .B1(new_n780), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n790), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n673), .A2(new_n248), .A3(new_n793), .A4(new_n779), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n283), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n775), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n637), .A2(new_n546), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT111), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n647), .A2(new_n616), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n802), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT111), .B1(new_n799), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(G113gat), .B1(new_n806), .B2(new_n251), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n799), .A2(new_n622), .A3(new_n616), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n730), .A2(new_n422), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT112), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n807), .A2(new_n811), .ZN(G1340gat));
  OAI21_X1  g611(.A(G120gat), .B1(new_n806), .B2(new_n336), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n808), .B(new_n335), .C1(new_n417), .C2(new_n416), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(G1341gat));
  NAND4_X1  g614(.A1(new_n803), .A2(G127gat), .A3(new_n283), .A4(new_n805), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n816), .A2(KEYINPUT113), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n816), .A2(KEYINPUT113), .ZN(new_n818));
  AOI21_X1  g617(.A(G127gat), .B1(new_n808), .B2(new_n283), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(G1342gat));
  INV_X1    g619(.A(new_n797), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n673), .A2(new_n546), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(KEYINPUT114), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n637), .A3(new_n823), .ZN(new_n824));
  NOR4_X1   g623(.A1(new_n824), .A2(new_n409), .A3(new_n622), .A4(new_n616), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT56), .ZN(new_n826));
  OAI21_X1  g625(.A(G134gat), .B1(new_n806), .B2(new_n316), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(G1343gat));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n780), .B2(new_n791), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n730), .A2(new_n793), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n248), .A2(new_n335), .A3(new_n779), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(KEYINPUT116), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n830), .A2(new_n833), .A3(new_n316), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n283), .B1(new_n834), .B2(new_n794), .ZN(new_n835));
  OAI211_X1 g634(.A(KEYINPUT57), .B(new_n616), .C1(new_n835), .C2(new_n775), .ZN(new_n836));
  XOR2_X1   g635(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n837));
  OAI21_X1  g636(.A(new_n837), .B1(new_n797), .B2(new_n399), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n689), .A2(new_n798), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(new_n730), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n839), .A2(KEYINPUT117), .A3(new_n730), .A4(new_n840), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(G141gat), .A3(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT58), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n799), .A2(new_n399), .A3(new_n658), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n368), .A3(new_n730), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT118), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n841), .A2(G141gat), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n848), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT58), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n845), .A2(new_n854), .A3(new_n846), .A4(new_n848), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n850), .A2(new_n853), .A3(new_n855), .ZN(G1344gat));
  NAND3_X1  g655(.A1(new_n847), .A2(new_n370), .A3(new_n335), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n839), .A2(new_n840), .ZN(new_n858));
  AOI211_X1 g657(.A(KEYINPUT59), .B(new_n370), .C1(new_n858), .C2(new_n335), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n834), .A2(new_n794), .ZN(new_n861));
  OAI22_X1  g660(.A1(new_n861), .A2(new_n283), .B1(new_n340), .B2(new_n730), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT57), .B1(new_n862), .B2(new_n616), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n821), .A2(new_n616), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(new_n837), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n335), .B(new_n840), .C1(new_n863), .C2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n860), .B1(new_n866), .B2(G148gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n857), .B1(new_n859), .B2(new_n867), .ZN(G1345gat));
  NAND3_X1  g667(.A1(new_n858), .A2(G155gat), .A3(new_n283), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n847), .A2(new_n283), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n360), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  XOR2_X1   g671(.A(new_n872), .B(KEYINPUT119), .Z(G1346gat));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n673), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n658), .A2(new_n399), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n824), .A2(G162gat), .ZN(new_n876));
  AOI22_X1  g675(.A1(new_n874), .A2(G162gat), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT120), .ZN(G1347gat));
  NOR2_X1   g677(.A1(new_n797), .A2(new_n637), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n879), .A2(new_n623), .A3(new_n582), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n881), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(G169gat), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n885), .A3(new_n730), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n879), .A2(new_n582), .A3(new_n802), .ZN(new_n887));
  OAI21_X1  g686(.A(G169gat), .B1(new_n887), .B2(new_n251), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(G1348gat));
  INV_X1    g688(.A(G176gat), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n882), .A2(new_n890), .A3(new_n335), .A4(new_n883), .ZN(new_n891));
  OAI21_X1  g690(.A(G176gat), .B1(new_n887), .B2(new_n336), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n893), .B(new_n894), .ZN(G1349gat));
  NAND3_X1  g694(.A1(new_n880), .A2(new_n283), .A3(new_n494), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT60), .ZN(new_n898));
  OAI21_X1  g697(.A(G183gat), .B1(new_n887), .B2(new_n796), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n897), .A2(KEYINPUT60), .ZN(new_n901));
  XOR2_X1   g700(.A(new_n900), .B(new_n901), .Z(G1350gat));
  NAND3_X1  g701(.A1(new_n884), .A2(new_n495), .A3(new_n673), .ZN(new_n903));
  OAI21_X1  g702(.A(G190gat), .B1(new_n887), .B2(new_n316), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT61), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(G1351gat));
  AND3_X1   g705(.A1(new_n875), .A2(new_n582), .A3(new_n879), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT124), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n236), .A3(new_n730), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n658), .A2(new_n637), .A3(new_n546), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(new_n863), .B2(new_n865), .ZN(new_n911));
  OAI21_X1  g710(.A(G197gat), .B1(new_n911), .B2(new_n251), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n909), .A2(new_n912), .ZN(G1352gat));
  OAI211_X1 g712(.A(new_n335), .B(new_n910), .C1(new_n863), .C2(new_n865), .ZN(new_n914));
  XNOR2_X1  g713(.A(KEYINPUT125), .B(G204gat), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n336), .A2(new_n915), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n907), .A2(new_n917), .ZN(new_n918));
  XOR2_X1   g717(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n907), .B(new_n917), .C1(KEYINPUT126), .C2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n916), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT127), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n923), .B(new_n924), .ZN(G1353gat));
  NAND3_X1  g724(.A1(new_n908), .A2(new_n283), .A3(new_n345), .ZN(new_n926));
  INV_X1    g725(.A(new_n911), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n283), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT63), .B1(new_n928), .B2(G211gat), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT63), .ZN(new_n930));
  AOI211_X1 g729(.A(new_n930), .B(new_n270), .C1(new_n927), .C2(new_n283), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n926), .B1(new_n929), .B2(new_n931), .ZN(G1354gat));
  NAND3_X1  g731(.A1(new_n908), .A2(new_n346), .A3(new_n673), .ZN(new_n933));
  OAI21_X1  g732(.A(G218gat), .B1(new_n911), .B2(new_n316), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1355gat));
endmodule


