

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779;

  NAND2_X1 U365 ( .A1(n385), .A2(n389), .ZN(n470) );
  NOR2_X1 U366 ( .A1(n545), .A2(n544), .ZN(n546) );
  AND2_X1 U367 ( .A1(n377), .A2(n378), .ZN(n359) );
  XOR2_X1 U368 ( .A(G478), .B(n578), .Z(n590) );
  BUF_X1 U369 ( .A(G143), .Z(n422) );
  NOR2_X2 U370 ( .A1(G953), .A2(G237), .ZN(n556) );
  XNOR2_X1 U371 ( .A(n417), .B(G146), .ZN(n412) );
  INV_X1 U372 ( .A(G125), .ZN(n417) );
  XNOR2_X2 U373 ( .A(n562), .B(n529), .ZN(n764) );
  XNOR2_X2 U374 ( .A(n764), .B(n532), .ZN(n537) );
  NOR2_X2 U375 ( .A1(n633), .A2(n352), .ZN(n497) );
  XNOR2_X2 U376 ( .A(n370), .B(KEYINPUT0), .ZN(n633) );
  INV_X2 U377 ( .A(G143), .ZN(n472) );
  BUF_X1 U378 ( .A(G113), .Z(n451) );
  AND2_X1 U379 ( .A1(n588), .A2(n628), .ZN(n344) );
  AND2_X2 U380 ( .A1(n482), .A2(n434), .ZN(n423) );
  AND2_X1 U381 ( .A1(n471), .A2(n661), .ZN(n495) );
  XNOR2_X2 U382 ( .A(n505), .B(n504), .ZN(n507) );
  XNOR2_X2 U383 ( .A(n537), .B(n536), .ZN(n373) );
  XNOR2_X2 U384 ( .A(n604), .B(n477), .ZN(n650) );
  XNOR2_X2 U385 ( .A(n579), .B(KEYINPUT40), .ZN(n778) );
  NAND2_X2 U386 ( .A1(n374), .A2(n686), .ZN(n579) );
  XNOR2_X1 U387 ( .A(n621), .B(KEYINPUT86), .ZN(n663) );
  INV_X1 U388 ( .A(n602), .ZN(n345) );
  INV_X1 U389 ( .A(KEYINPUT68), .ZN(n504) );
  INV_X2 U390 ( .A(G953), .ZN(n768) );
  AND2_X1 U391 ( .A1(n396), .A2(n392), .ZN(n391) );
  AND2_X1 U392 ( .A1(n489), .A2(n487), .ZN(n452) );
  AND2_X1 U393 ( .A1(n488), .A2(n697), .ZN(n487) );
  AND2_X1 U394 ( .A1(n386), .A2(n388), .ZN(n385) );
  AND2_X1 U395 ( .A1(n383), .A2(n631), .ZN(n388) );
  XNOR2_X1 U396 ( .A(n380), .B(KEYINPUT41), .ZN(n729) );
  XNOR2_X1 U397 ( .A(n381), .B(KEYINPUT115), .ZN(n720) );
  OR2_X1 U398 ( .A1(n636), .A2(n635), .ZN(n352) );
  XNOR2_X1 U399 ( .A(n450), .B(n494), .ZN(n715) );
  NOR2_X1 U400 ( .A1(n639), .A2(n652), .ZN(n640) );
  OR2_X2 U401 ( .A1(n428), .A2(n425), .ZN(n652) );
  BUF_X1 U402 ( .A(n562), .Z(n399) );
  XNOR2_X1 U403 ( .A(n412), .B(KEYINPUT10), .ZN(n562) );
  XOR2_X1 U404 ( .A(KEYINPUT23), .B(KEYINPUT94), .Z(n535) );
  XNOR2_X1 U405 ( .A(G122), .B(KEYINPUT16), .ZN(n354) );
  XNOR2_X1 U406 ( .A(G902), .B(KEYINPUT15), .ZN(n660) );
  NOR2_X2 U407 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U408 ( .A1(n547), .A2(n354), .ZN(n348) );
  NAND2_X1 U409 ( .A1(n346), .A2(n347), .ZN(n349) );
  NAND2_X1 U410 ( .A1(n348), .A2(n349), .ZN(n410) );
  INV_X1 U411 ( .A(n547), .ZN(n346) );
  INV_X1 U412 ( .A(n354), .ZN(n347) );
  XNOR2_X2 U413 ( .A(n410), .B(n372), .ZN(n400) );
  BUF_X1 U414 ( .A(n369), .Z(n350) );
  AND2_X2 U415 ( .A1(n446), .A2(n495), .ZN(n752) );
  OR2_X1 U416 ( .A1(G237), .A2(G902), .ZN(n553) );
  INV_X1 U417 ( .A(G469), .ZN(n439) );
  NAND2_X1 U418 ( .A1(n591), .A2(KEYINPUT71), .ZN(n459) );
  XNOR2_X1 U419 ( .A(n694), .B(n424), .ZN(n611) );
  NOR2_X1 U420 ( .A1(n593), .A2(n460), .ZN(n614) );
  XNOR2_X1 U421 ( .A(n583), .B(n584), .ZN(n492) );
  INV_X1 U422 ( .A(n580), .ZN(n419) );
  XOR2_X1 U423 ( .A(KEYINPUT4), .B(G131), .Z(n501) );
  XNOR2_X1 U424 ( .A(n525), .B(n526), .ZN(n548) );
  INV_X1 U425 ( .A(G101), .ZN(n526) );
  NAND2_X1 U426 ( .A1(n715), .A2(n714), .ZN(n381) );
  INV_X1 U427 ( .A(KEYINPUT33), .ZN(n435) );
  NAND2_X1 U428 ( .A1(n652), .A2(n634), .ZN(n379) );
  NAND2_X1 U429 ( .A1(n540), .A2(n427), .ZN(n426) );
  INV_X1 U430 ( .A(G902), .ZN(n427) );
  NAND2_X1 U431 ( .A1(n373), .A2(n431), .ZN(n430) );
  XNOR2_X1 U432 ( .A(G116), .B(G107), .ZN(n566) );
  INV_X1 U433 ( .A(n575), .ZN(n448) );
  XNOR2_X1 U434 ( .A(KEYINPUT7), .B(KEYINPUT105), .ZN(n568) );
  AND2_X1 U435 ( .A1(n415), .A2(n345), .ZN(n588) );
  XNOR2_X1 U436 ( .A(n416), .B(KEYINPUT28), .ZN(n415) );
  INV_X1 U437 ( .A(n379), .ZN(n699) );
  AND2_X1 U438 ( .A1(n393), .A2(n741), .ZN(n392) );
  INV_X1 U439 ( .A(n483), .ZN(n394) );
  INV_X1 U440 ( .A(KEYINPUT75), .ZN(n402) );
  NOR2_X1 U441 ( .A1(n663), .A2(n502), .ZN(n659) );
  INV_X1 U442 ( .A(n755), .ZN(n741) );
  INV_X1 U443 ( .A(KEYINPUT87), .ZN(n424) );
  AND2_X1 U444 ( .A1(n344), .A2(n454), .ZN(n453) );
  NAND2_X1 U445 ( .A1(n344), .A2(n351), .ZN(n456) );
  XOR2_X1 U446 ( .A(KEYINPUT95), .B(KEYINPUT21), .Z(n543) );
  INV_X1 U447 ( .A(G134), .ZN(n503) );
  NOR2_X1 U448 ( .A1(n485), .A2(n414), .ZN(n413) );
  XNOR2_X1 U449 ( .A(G104), .B(G122), .ZN(n560) );
  INV_X1 U450 ( .A(G140), .ZN(n467) );
  XOR2_X1 U451 ( .A(KEYINPUT11), .B(n422), .Z(n555) );
  XNOR2_X1 U452 ( .A(n551), .B(n444), .ZN(n443) );
  XNOR2_X1 U453 ( .A(n552), .B(KEYINPUT17), .ZN(n444) );
  INV_X1 U454 ( .A(KEYINPUT38), .ZN(n494) );
  NOR2_X1 U455 ( .A1(n646), .A2(KEYINPUT34), .ZN(n387) );
  INV_X1 U456 ( .A(KEYINPUT72), .ZN(n629) );
  NAND2_X1 U457 ( .A1(n379), .A2(n420), .ZN(n377) );
  XNOR2_X1 U458 ( .A(KEYINPUT30), .B(KEYINPUT114), .ZN(n517) );
  XNOR2_X1 U459 ( .A(n564), .B(n463), .ZN(n597) );
  XNOR2_X1 U460 ( .A(n563), .B(G475), .ZN(n463) );
  INV_X1 U461 ( .A(KEYINPUT6), .ZN(n477) );
  INV_X1 U462 ( .A(n548), .ZN(n372) );
  XNOR2_X1 U463 ( .A(G119), .B(G128), .ZN(n530) );
  XNOR2_X1 U464 ( .A(n465), .B(n464), .ZN(n670) );
  XNOR2_X1 U465 ( .A(n399), .B(n466), .ZN(n465) );
  XNOR2_X1 U466 ( .A(n559), .B(n561), .ZN(n464) );
  XNOR2_X1 U467 ( .A(n560), .B(n467), .ZN(n466) );
  XNOR2_X1 U468 ( .A(n528), .B(n527), .ZN(n742) );
  XNOR2_X1 U469 ( .A(n548), .B(n449), .ZN(n527) );
  XNOR2_X1 U470 ( .A(n529), .B(n361), .ZN(n449) );
  INV_X1 U471 ( .A(KEYINPUT90), .ZN(n585) );
  NAND2_X1 U472 ( .A1(n713), .A2(KEYINPUT34), .ZN(n389) );
  XNOR2_X1 U473 ( .A(n597), .B(n462), .ZN(n589) );
  INV_X1 U474 ( .A(KEYINPUT103), .ZN(n462) );
  NAND2_X1 U475 ( .A1(n430), .A2(n429), .ZN(n428) );
  NAND2_X1 U476 ( .A1(n431), .A2(G902), .ZN(n429) );
  XNOR2_X1 U477 ( .A(n574), .B(n447), .ZN(n749) );
  XNOR2_X1 U478 ( .A(n448), .B(n573), .ZN(n447) );
  XNOR2_X1 U479 ( .A(n670), .B(KEYINPUT59), .ZN(n671) );
  NAND2_X1 U480 ( .A1(n729), .A2(n588), .ZN(n484) );
  NAND2_X1 U481 ( .A1(n391), .A2(n390), .ZN(n398) );
  INV_X1 U482 ( .A(KEYINPUT56), .ZN(n473) );
  AND2_X1 U483 ( .A1(n719), .A2(n366), .ZN(n351) );
  XOR2_X1 U484 ( .A(KEYINPUT74), .B(G107), .Z(n353) );
  XOR2_X1 U485 ( .A(n643), .B(KEYINPUT81), .Z(n355) );
  AND2_X1 U486 ( .A1(n469), .A2(n468), .ZN(n356) );
  AND2_X1 U487 ( .A1(n345), .A2(n418), .ZN(n357) );
  AND2_X1 U488 ( .A1(n699), .A2(n345), .ZN(n358) );
  NOR2_X1 U489 ( .A1(n589), .A2(n590), .ZN(n360) );
  INV_X1 U490 ( .A(n604), .ZN(n705) );
  AND2_X1 U491 ( .A1(G227), .A2(n768), .ZN(n361) );
  AND2_X1 U492 ( .A1(n553), .A2(G210), .ZN(n362) );
  INV_X1 U493 ( .A(n441), .ZN(n411) );
  XNOR2_X1 U494 ( .A(n443), .B(n442), .ZN(n441) );
  AND2_X1 U495 ( .A1(n638), .A2(KEYINPUT88), .ZN(n363) );
  INV_X1 U496 ( .A(n650), .ZN(n437) );
  XOR2_X1 U497 ( .A(n632), .B(KEYINPUT35), .Z(n364) );
  XOR2_X1 U498 ( .A(n637), .B(KEYINPUT22), .Z(n365) );
  INV_X1 U499 ( .A(n591), .ZN(n461) );
  AND2_X1 U500 ( .A1(n461), .A2(n458), .ZN(n366) );
  INV_X1 U501 ( .A(KEYINPUT77), .ZN(n420) );
  XOR2_X1 U502 ( .A(n740), .B(n739), .Z(n367) );
  AND2_X1 U503 ( .A1(n661), .A2(G478), .ZN(n368) );
  INV_X1 U504 ( .A(KEYINPUT71), .ZN(n458) );
  XNOR2_X1 U505 ( .A(n369), .B(n587), .ZN(n628) );
  NAND2_X1 U506 ( .A1(n615), .A2(n350), .ZN(n608) );
  XNOR2_X2 U507 ( .A(n479), .B(n585), .ZN(n369) );
  NAND2_X1 U508 ( .A1(n628), .A2(n627), .ZN(n370) );
  NAND2_X1 U509 ( .A1(n371), .A2(n659), .ZN(n403) );
  XNOR2_X2 U510 ( .A(n658), .B(KEYINPUT45), .ZN(n371) );
  NAND2_X1 U511 ( .A1(n767), .A2(n371), .ZN(n665) );
  NAND2_X1 U512 ( .A1(n371), .A2(n768), .ZN(n759) );
  XNOR2_X1 U513 ( .A(n400), .B(n441), .ZN(n738) );
  NOR2_X1 U514 ( .A1(n426), .A2(n373), .ZN(n425) );
  XNOR2_X1 U515 ( .A(n753), .B(n373), .ZN(n754) );
  NAND2_X1 U516 ( .A1(n374), .A2(n360), .ZN(n662) );
  XNOR2_X2 U517 ( .A(n432), .B(KEYINPUT39), .ZN(n374) );
  NAND2_X1 U518 ( .A1(n375), .A2(n420), .ZN(n378) );
  NAND2_X1 U519 ( .A1(n345), .A2(n419), .ZN(n375) );
  NAND2_X1 U520 ( .A1(n359), .A2(n376), .ZN(n544) );
  NAND2_X1 U521 ( .A1(n357), .A2(n699), .ZN(n376) );
  NAND2_X1 U522 ( .A1(n720), .A2(n718), .ZN(n380) );
  NAND2_X1 U523 ( .A1(n382), .A2(n705), .ZN(n710) );
  XNOR2_X1 U524 ( .A(n382), .B(KEYINPUT112), .ZN(n438) );
  XNOR2_X2 U525 ( .A(n630), .B(n629), .ZN(n382) );
  NAND2_X1 U526 ( .A1(n646), .A2(KEYINPUT34), .ZN(n383) );
  NAND2_X1 U527 ( .A1(n384), .A2(n387), .ZN(n386) );
  INV_X1 U528 ( .A(n713), .ZN(n384) );
  XNOR2_X2 U529 ( .A(n436), .B(n435), .ZN(n713) );
  OR2_X1 U530 ( .A1(n669), .A2(n483), .ZN(n390) );
  NAND2_X1 U531 ( .A1(n395), .A2(n394), .ZN(n393) );
  INV_X1 U532 ( .A(n666), .ZN(n395) );
  NAND2_X1 U533 ( .A1(n669), .A2(n397), .ZN(n396) );
  AND2_X1 U534 ( .A1(n666), .A2(n483), .ZN(n397) );
  XNOR2_X1 U535 ( .A(n398), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U536 ( .A(n668), .B(n667), .ZN(n483) );
  OR2_X2 U537 ( .A1(n668), .A2(G902), .ZN(n478) );
  INV_X1 U538 ( .A(n400), .ZN(n401) );
  XNOR2_X2 U539 ( .A(n403), .B(n402), .ZN(n446) );
  XNOR2_X1 U540 ( .A(n451), .B(G131), .ZN(n554) );
  BUF_X1 U541 ( .A(n752), .Z(n404) );
  NAND2_X1 U542 ( .A1(n475), .A2(n741), .ZN(n474) );
  XNOR2_X1 U543 ( .A(n476), .B(n367), .ZN(n475) );
  NOR2_X1 U544 ( .A1(n605), .A2(n604), .ZN(n416) );
  XNOR2_X1 U545 ( .A(n528), .B(n515), .ZN(n668) );
  XNOR2_X1 U546 ( .A(n644), .B(KEYINPUT32), .ZN(n405) );
  XNOR2_X1 U547 ( .A(n644), .B(KEYINPUT32), .ZN(n779) );
  BUF_X1 U548 ( .A(n766), .Z(n406) );
  AND2_X1 U549 ( .A1(n500), .A2(n638), .ZN(n407) );
  XNOR2_X1 U550 ( .A(n401), .B(n411), .ZN(n408) );
  XNOR2_X1 U551 ( .A(n497), .B(n365), .ZN(n421) );
  NAND2_X1 U552 ( .A1(n421), .A2(n639), .ZN(n651) );
  BUF_X1 U553 ( .A(n405), .Z(n409) );
  XNOR2_X2 U554 ( .A(n507), .B(n506), .ZN(n547) );
  XNOR2_X1 U555 ( .A(n401), .B(KEYINPUT124), .ZN(n760) );
  XNOR2_X1 U556 ( .A(n433), .B(n412), .ZN(n442) );
  NAND2_X1 U557 ( .A1(n491), .A2(n413), .ZN(n490) );
  INV_X1 U558 ( .A(n613), .ZN(n414) );
  NAND2_X1 U559 ( .A1(n701), .A2(n582), .ZN(n605) );
  NOR2_X1 U560 ( .A1(n580), .A2(n420), .ZN(n418) );
  AND2_X2 U561 ( .A1(n421), .A2(n355), .ZN(n644) );
  NAND2_X1 U562 ( .A1(n738), .A2(n660), .ZN(n445) );
  OR2_X2 U563 ( .A1(n742), .A2(G902), .ZN(n440) );
  NAND2_X1 U564 ( .A1(n423), .A2(n356), .ZN(n481) );
  NOR2_X2 U565 ( .A1(n689), .A2(n607), .ZN(n615) );
  NOR2_X2 U566 ( .A1(n610), .A2(n639), .ZN(n694) );
  INV_X1 U567 ( .A(n540), .ZN(n431) );
  NAND2_X1 U568 ( .A1(n599), .A2(n715), .ZN(n432) );
  XNOR2_X1 U569 ( .A(n546), .B(KEYINPUT76), .ZN(n599) );
  XNOR2_X2 U570 ( .A(n433), .B(n503), .ZN(n565) );
  XNOR2_X2 U571 ( .A(n472), .B(G128), .ZN(n433) );
  XNOR2_X1 U572 ( .A(n434), .B(G122), .ZN(G24) );
  XNOR2_X2 U573 ( .A(n470), .B(n364), .ZN(n434) );
  NAND2_X1 U574 ( .A1(n438), .A2(n437), .ZN(n436) );
  XNOR2_X2 U575 ( .A(n440), .B(n439), .ZN(n602) );
  XNOR2_X2 U576 ( .A(n766), .B(G146), .ZN(n528) );
  XNOR2_X2 U577 ( .A(n445), .B(n362), .ZN(n618) );
  NAND2_X1 U578 ( .A1(n446), .A2(n496), .ZN(n748) );
  AND2_X1 U579 ( .A1(n446), .A2(n661), .ZN(n669) );
  NAND2_X1 U580 ( .A1(n446), .A2(n471), .ZN(n734) );
  NAND2_X2 U581 ( .A1(n618), .A2(n714), .ZN(n479) );
  NOR2_X2 U582 ( .A1(n598), .A2(n597), .ZN(n718) );
  NAND2_X1 U583 ( .A1(n778), .A2(n777), .ZN(n583) );
  XNOR2_X2 U584 ( .A(n602), .B(n603), .ZN(n698) );
  NAND2_X1 U585 ( .A1(n752), .A2(G210), .ZN(n476) );
  NAND2_X1 U586 ( .A1(n405), .A2(KEYINPUT88), .ZN(n468) );
  BUF_X1 U587 ( .A(n618), .Z(n450) );
  NOR2_X2 U588 ( .A1(n663), .A2(n696), .ZN(n767) );
  NAND2_X1 U589 ( .A1(n452), .A2(n490), .ZN(n621) );
  NAND2_X1 U590 ( .A1(n455), .A2(n453), .ZN(n457) );
  NAND2_X1 U591 ( .A1(n459), .A2(n458), .ZN(n454) );
  NAND2_X1 U592 ( .A1(n719), .A2(n459), .ZN(n455) );
  NAND2_X1 U593 ( .A1(n457), .A2(n456), .ZN(n460) );
  NAND2_X1 U594 ( .A1(n500), .A2(n363), .ZN(n469) );
  XNOR2_X2 U595 ( .A(n651), .B(KEYINPUT111), .ZN(n500) );
  AND2_X1 U596 ( .A1(n471), .A2(n368), .ZN(n496) );
  AND2_X1 U597 ( .A1(n471), .A2(G472), .ZN(n666) );
  NAND2_X2 U598 ( .A1(n665), .A2(n664), .ZN(n471) );
  XNOR2_X1 U599 ( .A(n474), .B(n473), .ZN(G51) );
  XNOR2_X2 U600 ( .A(n478), .B(n516), .ZN(n604) );
  XNOR2_X1 U601 ( .A(n481), .B(n480), .ZN(n657) );
  INV_X1 U602 ( .A(KEYINPUT44), .ZN(n480) );
  NAND2_X1 U603 ( .A1(n499), .A2(n498), .ZN(n482) );
  XNOR2_X2 U604 ( .A(n484), .B(KEYINPUT42), .ZN(n777) );
  NAND2_X1 U605 ( .A1(n613), .A2(n614), .ZN(n493) );
  NAND2_X1 U606 ( .A1(n614), .A2(n486), .ZN(n485) );
  INV_X1 U607 ( .A(KEYINPUT48), .ZN(n486) );
  NAND2_X1 U608 ( .A1(n493), .A2(KEYINPUT48), .ZN(n488) );
  NAND2_X1 U609 ( .A1(n492), .A2(KEYINPUT48), .ZN(n489) );
  INV_X1 U610 ( .A(n492), .ZN(n491) );
  NAND2_X1 U611 ( .A1(n500), .A2(n638), .ZN(n499) );
  NOR2_X1 U612 ( .A1(n779), .A2(KEYINPUT88), .ZN(n498) );
  XOR2_X1 U613 ( .A(KEYINPUT83), .B(n622), .Z(n502) );
  INV_X1 U614 ( .A(n713), .ZN(n730) );
  INV_X1 U615 ( .A(n634), .ZN(n635) );
  XNOR2_X1 U616 ( .A(n518), .B(n517), .ZN(n545) );
  XNOR2_X1 U617 ( .A(n514), .B(n547), .ZN(n515) );
  XNOR2_X1 U618 ( .A(n539), .B(KEYINPUT25), .ZN(n540) );
  XNOR2_X1 U619 ( .A(n672), .B(n671), .ZN(n673) );
  NOR2_X1 U620 ( .A1(G952), .A2(n768), .ZN(n755) );
  XNOR2_X2 U621 ( .A(n565), .B(n501), .ZN(n766) );
  XNOR2_X2 U622 ( .A(G116), .B(G113), .ZN(n505) );
  XOR2_X1 U623 ( .A(KEYINPUT3), .B(G119), .Z(n506) );
  XOR2_X1 U624 ( .A(KEYINPUT5), .B(KEYINPUT97), .Z(n509) );
  NAND2_X1 U625 ( .A1(n556), .A2(G210), .ZN(n508) );
  XNOR2_X1 U626 ( .A(n509), .B(n508), .ZN(n513) );
  XOR2_X1 U627 ( .A(KEYINPUT98), .B(KEYINPUT73), .Z(n511) );
  XNOR2_X1 U628 ( .A(G101), .B(G137), .ZN(n510) );
  XNOR2_X1 U629 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U630 ( .A(n513), .B(n512), .Z(n514) );
  XOR2_X1 U631 ( .A(KEYINPUT116), .B(KEYINPUT62), .Z(n667) );
  XNOR2_X1 U632 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n584) );
  NAND2_X1 U633 ( .A1(G214), .A2(n553), .ZN(n714) );
  XNOR2_X1 U634 ( .A(G472), .B(KEYINPUT99), .ZN(n516) );
  NAND2_X1 U635 ( .A1(n714), .A2(n705), .ZN(n518) );
  NAND2_X1 U636 ( .A1(G234), .A2(G237), .ZN(n519) );
  XNOR2_X1 U637 ( .A(n519), .B(KEYINPUT14), .ZN(n520) );
  NAND2_X1 U638 ( .A1(G952), .A2(n520), .ZN(n728) );
  NOR2_X1 U639 ( .A1(G953), .A2(n728), .ZN(n624) );
  NAND2_X1 U640 ( .A1(n520), .A2(G902), .ZN(n521) );
  XNOR2_X1 U641 ( .A(n521), .B(KEYINPUT93), .ZN(n623) );
  NAND2_X1 U642 ( .A1(G953), .A2(n623), .ZN(n522) );
  NOR2_X1 U643 ( .A1(G900), .A2(n522), .ZN(n523) );
  NOR2_X1 U644 ( .A1(n624), .A2(n523), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G110), .B(G104), .ZN(n524) );
  XNOR2_X1 U646 ( .A(n353), .B(n524), .ZN(n525) );
  XOR2_X1 U647 ( .A(G137), .B(G140), .Z(n529) );
  XOR2_X1 U648 ( .A(KEYINPUT24), .B(G110), .Z(n531) );
  XNOR2_X1 U649 ( .A(n531), .B(n530), .ZN(n532) );
  NAND2_X1 U650 ( .A1(G234), .A2(n768), .ZN(n533) );
  XOR2_X1 U651 ( .A(KEYINPUT8), .B(n533), .Z(n572) );
  NAND2_X1 U652 ( .A1(G221), .A2(n572), .ZN(n534) );
  XNOR2_X1 U653 ( .A(n535), .B(n534), .ZN(n536) );
  NAND2_X1 U654 ( .A1(G234), .A2(n660), .ZN(n538) );
  XNOR2_X1 U655 ( .A(KEYINPUT20), .B(n538), .ZN(n541) );
  NAND2_X1 U656 ( .A1(G217), .A2(n541), .ZN(n539) );
  NAND2_X1 U657 ( .A1(n541), .A2(G221), .ZN(n542) );
  XNOR2_X1 U658 ( .A(n543), .B(n542), .ZN(n702) );
  XOR2_X1 U659 ( .A(n702), .B(KEYINPUT96), .Z(n634) );
  XOR2_X1 U660 ( .A(KEYINPUT92), .B(KEYINPUT18), .Z(n550) );
  XNOR2_X1 U661 ( .A(KEYINPUT4), .B(KEYINPUT79), .ZN(n549) );
  XNOR2_X1 U662 ( .A(n550), .B(n549), .ZN(n551) );
  NAND2_X1 U663 ( .A1(G224), .A2(n768), .ZN(n552) );
  XNOR2_X1 U664 ( .A(n555), .B(n554), .ZN(n561) );
  XOR2_X1 U665 ( .A(KEYINPUT12), .B(KEYINPUT101), .Z(n558) );
  NAND2_X1 U666 ( .A1(G214), .A2(n556), .ZN(n557) );
  XNOR2_X1 U667 ( .A(n558), .B(n557), .ZN(n559) );
  NOR2_X1 U668 ( .A1(G902), .A2(n670), .ZN(n564) );
  XNOR2_X1 U669 ( .A(KEYINPUT102), .B(KEYINPUT13), .ZN(n563) );
  INV_X1 U670 ( .A(n565), .ZN(n575) );
  XOR2_X1 U671 ( .A(KEYINPUT106), .B(G122), .Z(n567) );
  XNOR2_X1 U672 ( .A(n567), .B(n566), .ZN(n571) );
  XOR2_X1 U673 ( .A(KEYINPUT104), .B(KEYINPUT9), .Z(n569) );
  XNOR2_X1 U674 ( .A(n569), .B(n568), .ZN(n570) );
  XOR2_X1 U675 ( .A(n571), .B(n570), .Z(n574) );
  NAND2_X1 U676 ( .A1(G217), .A2(n572), .ZN(n573) );
  NOR2_X1 U677 ( .A1(G902), .A2(n749), .ZN(n577) );
  XNOR2_X1 U678 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n576) );
  XNOR2_X1 U679 ( .A(n577), .B(n576), .ZN(n578) );
  NAND2_X1 U680 ( .A1(n589), .A2(n590), .ZN(n689) );
  INV_X1 U681 ( .A(n689), .ZN(n686) );
  INV_X1 U682 ( .A(n652), .ZN(n701) );
  NOR2_X1 U683 ( .A1(n702), .A2(n580), .ZN(n581) );
  XOR2_X1 U684 ( .A(KEYINPUT67), .B(n581), .Z(n582) );
  INV_X1 U685 ( .A(n590), .ZN(n598) );
  XOR2_X1 U686 ( .A(KEYINPUT78), .B(KEYINPUT65), .Z(n586) );
  XOR2_X1 U687 ( .A(KEYINPUT19), .B(n586), .Z(n587) );
  INV_X1 U688 ( .A(n360), .ZN(n692) );
  NAND2_X1 U689 ( .A1(n689), .A2(n692), .ZN(n719) );
  INV_X1 U690 ( .A(n719), .ZN(n594) );
  XNOR2_X1 U691 ( .A(KEYINPUT66), .B(KEYINPUT47), .ZN(n591) );
  AND2_X1 U692 ( .A1(KEYINPUT47), .A2(n594), .ZN(n592) );
  NOR2_X1 U693 ( .A1(KEYINPUT84), .A2(n592), .ZN(n593) );
  NAND2_X1 U694 ( .A1(n594), .A2(KEYINPUT84), .ZN(n595) );
  NAND2_X1 U695 ( .A1(n595), .A2(n344), .ZN(n596) );
  NAND2_X1 U696 ( .A1(n596), .A2(KEYINPUT47), .ZN(n601) );
  AND2_X1 U697 ( .A1(n598), .A2(n597), .ZN(n631) );
  AND2_X1 U698 ( .A1(n599), .A2(n631), .ZN(n600) );
  NAND2_X1 U699 ( .A1(n450), .A2(n600), .ZN(n685) );
  NAND2_X1 U700 ( .A1(n601), .A2(n685), .ZN(n612) );
  INV_X1 U701 ( .A(KEYINPUT1), .ZN(n603) );
  INV_X1 U702 ( .A(n698), .ZN(n639) );
  XOR2_X1 U703 ( .A(KEYINPUT89), .B(KEYINPUT36), .Z(n609) );
  NOR2_X1 U704 ( .A1(n650), .A2(n605), .ZN(n606) );
  XNOR2_X1 U705 ( .A(n606), .B(KEYINPUT113), .ZN(n607) );
  XNOR2_X1 U706 ( .A(n609), .B(n608), .ZN(n610) );
  AND2_X1 U707 ( .A1(n639), .A2(n615), .ZN(n616) );
  NAND2_X1 U708 ( .A1(n616), .A2(n714), .ZN(n617) );
  XNOR2_X1 U709 ( .A(n617), .B(KEYINPUT43), .ZN(n620) );
  INV_X1 U710 ( .A(n450), .ZN(n619) );
  NAND2_X1 U711 ( .A1(n620), .A2(n619), .ZN(n697) );
  NAND2_X1 U712 ( .A1(KEYINPUT2), .A2(n662), .ZN(n622) );
  NOR2_X1 U713 ( .A1(G898), .A2(n768), .ZN(n761) );
  NAND2_X1 U714 ( .A1(n761), .A2(n623), .ZN(n626) );
  INV_X1 U715 ( .A(n624), .ZN(n625) );
  NAND2_X1 U716 ( .A1(n626), .A2(n625), .ZN(n627) );
  BUF_X2 U717 ( .A(n633), .Z(n646) );
  NAND2_X1 U718 ( .A1(n699), .A2(n698), .ZN(n630) );
  XOR2_X1 U719 ( .A(KEYINPUT80), .B(KEYINPUT85), .Z(n632) );
  INV_X1 U720 ( .A(n718), .ZN(n636) );
  XNOR2_X1 U721 ( .A(KEYINPUT70), .B(KEYINPUT69), .ZN(n637) );
  AND2_X1 U722 ( .A1(n701), .A2(n604), .ZN(n638) );
  XOR2_X1 U723 ( .A(KEYINPUT110), .B(n640), .Z(n642) );
  XOR2_X1 U724 ( .A(n650), .B(KEYINPUT82), .Z(n641) );
  NOR2_X1 U725 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U726 ( .A1(n646), .A2(n710), .ZN(n645) );
  XNOR2_X1 U727 ( .A(n645), .B(KEYINPUT31), .ZN(n691) );
  NOR2_X1 U728 ( .A1(n705), .A2(n646), .ZN(n647) );
  NAND2_X1 U729 ( .A1(n358), .A2(n647), .ZN(n648) );
  XNOR2_X1 U730 ( .A(KEYINPUT100), .B(n648), .ZN(n678) );
  NAND2_X1 U731 ( .A1(n691), .A2(n678), .ZN(n649) );
  NAND2_X1 U732 ( .A1(n649), .A2(n719), .ZN(n654) );
  NOR2_X1 U733 ( .A1(n437), .A2(n651), .ZN(n653) );
  NAND2_X1 U734 ( .A1(n653), .A2(n652), .ZN(n676) );
  NAND2_X1 U735 ( .A1(n654), .A2(n676), .ZN(n655) );
  XNOR2_X1 U736 ( .A(KEYINPUT109), .B(n655), .ZN(n656) );
  NAND2_X1 U737 ( .A1(n657), .A2(n656), .ZN(n658) );
  INV_X1 U738 ( .A(n660), .ZN(n661) );
  INV_X1 U739 ( .A(n662), .ZN(n696) );
  INV_X1 U740 ( .A(KEYINPUT2), .ZN(n664) );
  NAND2_X1 U741 ( .A1(n752), .A2(G475), .ZN(n672) );
  NAND2_X1 U742 ( .A1(n673), .A2(n741), .ZN(n675) );
  INV_X1 U743 ( .A(KEYINPUT60), .ZN(n674) );
  XNOR2_X1 U744 ( .A(n675), .B(n674), .ZN(G60) );
  XNOR2_X1 U745 ( .A(G101), .B(n676), .ZN(G3) );
  NOR2_X1 U746 ( .A1(n678), .A2(n689), .ZN(n677) );
  XOR2_X1 U747 ( .A(G104), .B(n677), .Z(G6) );
  NOR2_X1 U748 ( .A1(n678), .A2(n692), .ZN(n680) );
  XNOR2_X1 U749 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n679) );
  XNOR2_X1 U750 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U751 ( .A(G107), .B(n681), .ZN(G9) );
  XOR2_X1 U752 ( .A(G110), .B(n407), .Z(G12) );
  XOR2_X1 U753 ( .A(KEYINPUT29), .B(KEYINPUT117), .Z(n683) );
  NAND2_X1 U754 ( .A1(n360), .A2(n344), .ZN(n682) );
  XNOR2_X1 U755 ( .A(n683), .B(n682), .ZN(n684) );
  XOR2_X1 U756 ( .A(G128), .B(n684), .Z(G30) );
  XNOR2_X1 U757 ( .A(n422), .B(n685), .ZN(G45) );
  NAND2_X1 U758 ( .A1(n344), .A2(n686), .ZN(n687) );
  XNOR2_X1 U759 ( .A(n687), .B(KEYINPUT118), .ZN(n688) );
  XNOR2_X1 U760 ( .A(G146), .B(n688), .ZN(G48) );
  NOR2_X1 U761 ( .A1(n689), .A2(n691), .ZN(n690) );
  XOR2_X1 U762 ( .A(n451), .B(n690), .Z(G15) );
  NOR2_X1 U763 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U764 ( .A(G116), .B(n693), .Z(G18) );
  XNOR2_X1 U765 ( .A(G125), .B(n694), .ZN(n695) );
  XNOR2_X1 U766 ( .A(n695), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U767 ( .A(G134), .B(n696), .Z(G36) );
  XNOR2_X1 U768 ( .A(G140), .B(n697), .ZN(G42) );
  NOR2_X1 U769 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U770 ( .A(KEYINPUT50), .B(n700), .Z(n708) );
  XOR2_X1 U771 ( .A(KEYINPUT49), .B(KEYINPUT119), .Z(n704) );
  NAND2_X1 U772 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U773 ( .A(n704), .B(n703), .ZN(n706) );
  NOR2_X1 U774 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U775 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U776 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U777 ( .A(KEYINPUT51), .B(n711), .Z(n712) );
  NAND2_X1 U778 ( .A1(n729), .A2(n712), .ZN(n725) );
  NOR2_X1 U779 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U780 ( .A(KEYINPUT120), .B(n716), .Z(n717) );
  NAND2_X1 U781 ( .A1(n718), .A2(n717), .ZN(n722) );
  NAND2_X1 U782 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U783 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U784 ( .A1(n730), .A2(n723), .ZN(n724) );
  NAND2_X1 U785 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U786 ( .A(KEYINPUT52), .B(n726), .Z(n727) );
  NOR2_X1 U787 ( .A1(n728), .A2(n727), .ZN(n733) );
  AND2_X1 U788 ( .A1(n729), .A2(n730), .ZN(n731) );
  XOR2_X1 U789 ( .A(KEYINPUT121), .B(n731), .Z(n732) );
  NOR2_X1 U790 ( .A1(n733), .A2(n732), .ZN(n735) );
  NAND2_X1 U791 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U792 ( .A1(n736), .A2(G953), .ZN(n737) );
  XNOR2_X1 U793 ( .A(n737), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U794 ( .A(KEYINPUT91), .B(KEYINPUT55), .Z(n740) );
  XNOR2_X1 U795 ( .A(n408), .B(KEYINPUT54), .ZN(n739) );
  XNOR2_X1 U796 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n744) );
  XNOR2_X1 U797 ( .A(n742), .B(KEYINPUT57), .ZN(n743) );
  XNOR2_X1 U798 ( .A(n744), .B(n743), .ZN(n746) );
  NAND2_X1 U799 ( .A1(n752), .A2(G469), .ZN(n745) );
  XOR2_X1 U800 ( .A(n746), .B(n745), .Z(n747) );
  NOR2_X1 U801 ( .A1(n755), .A2(n747), .ZN(G54) );
  XNOR2_X1 U802 ( .A(n748), .B(KEYINPUT123), .ZN(n750) );
  XOR2_X1 U803 ( .A(n750), .B(n749), .Z(n751) );
  NOR2_X1 U804 ( .A1(n755), .A2(n751), .ZN(G63) );
  NAND2_X1 U805 ( .A1(G217), .A2(n404), .ZN(n753) );
  NOR2_X1 U806 ( .A1(n755), .A2(n754), .ZN(G66) );
  NAND2_X1 U807 ( .A1(G953), .A2(G224), .ZN(n756) );
  XNOR2_X1 U808 ( .A(KEYINPUT61), .B(n756), .ZN(n757) );
  NAND2_X1 U809 ( .A1(n757), .A2(G898), .ZN(n758) );
  NAND2_X1 U810 ( .A1(n759), .A2(n758), .ZN(n763) );
  NOR2_X1 U811 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U812 ( .A(n763), .B(n762), .ZN(G69) );
  XOR2_X1 U813 ( .A(n764), .B(KEYINPUT125), .Z(n765) );
  XNOR2_X1 U814 ( .A(n406), .B(n765), .ZN(n770) );
  XNOR2_X1 U815 ( .A(n770), .B(n767), .ZN(n769) );
  NAND2_X1 U816 ( .A1(n769), .A2(n768), .ZN(n775) );
  XNOR2_X1 U817 ( .A(G227), .B(n770), .ZN(n771) );
  NAND2_X1 U818 ( .A1(n771), .A2(G900), .ZN(n772) );
  XOR2_X1 U819 ( .A(KEYINPUT126), .B(n772), .Z(n773) );
  NAND2_X1 U820 ( .A1(G953), .A2(n773), .ZN(n774) );
  NAND2_X1 U821 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U822 ( .A(KEYINPUT127), .B(n776), .ZN(G72) );
  XNOR2_X1 U823 ( .A(G137), .B(n777), .ZN(G39) );
  XNOR2_X1 U824 ( .A(n778), .B(G131), .ZN(G33) );
  XOR2_X1 U825 ( .A(n409), .B(G119), .Z(G21) );
endmodule

