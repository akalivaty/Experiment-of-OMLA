

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U551 ( .A1(n596), .A2(n595), .ZN(n966) );
  OR2_X2 U552 ( .A1(KEYINPUT33), .A2(n765), .ZN(n518) );
  NOR2_X2 U553 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X2 U554 ( .A1(n697), .A2(n800), .ZN(n704) );
  NOR2_X2 U555 ( .A1(G164), .A2(G1384), .ZN(n800) );
  NOR2_X2 U556 ( .A1(n529), .A2(n528), .ZN(G164) );
  INV_X1 U557 ( .A(G2104), .ZN(n519) );
  OR2_X1 U558 ( .A1(n718), .A2(n977), .ZN(n516) );
  OR2_X1 U559 ( .A1(n766), .A2(n779), .ZN(n517) );
  NOR2_X1 U560 ( .A1(n731), .A2(n730), .ZN(n732) );
  AND2_X1 U561 ( .A1(n749), .A2(n748), .ZN(n751) );
  AND2_X1 U562 ( .A1(n983), .A2(n517), .ZN(n767) );
  INV_X1 U563 ( .A(n824), .ZN(n811) );
  NOR2_X1 U564 ( .A1(n821), .A2(n811), .ZN(n812) );
  INV_X1 U565 ( .A(KEYINPUT100), .ZN(n814) );
  INV_X1 U566 ( .A(KEYINPUT13), .ZN(n591) );
  NOR2_X1 U567 ( .A1(G651), .A2(G543), .ZN(n655) );
  NAND2_X1 U568 ( .A1(n519), .A2(n524), .ZN(n520) );
  XNOR2_X1 U569 ( .A(n815), .B(n814), .ZN(n817) );
  XNOR2_X2 U570 ( .A(n520), .B(KEYINPUT17), .ZN(n897) );
  NAND2_X1 U571 ( .A1(n897), .A2(G138), .ZN(n523) );
  INV_X1 U572 ( .A(G2105), .ZN(n524) );
  NOR2_X1 U573 ( .A1(G2104), .A2(n524), .ZN(n618) );
  NAND2_X1 U574 ( .A1(G126), .A2(n618), .ZN(n521) );
  XOR2_X1 U575 ( .A(KEYINPUT87), .B(n521), .Z(n522) );
  NAND2_X1 U576 ( .A1(n523), .A2(n522), .ZN(n529) );
  AND2_X1 U577 ( .A1(n524), .A2(G2104), .ZN(n898) );
  NAND2_X1 U578 ( .A1(G102), .A2(n898), .ZN(n527) );
  NAND2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n525) );
  XOR2_X1 U580 ( .A(KEYINPUT66), .B(n525), .Z(n615) );
  NAND2_X1 U581 ( .A1(G114), .A2(n615), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n527), .A2(n526), .ZN(n528) );
  NAND2_X1 U583 ( .A1(G91), .A2(n655), .ZN(n531) );
  XOR2_X1 U584 ( .A(KEYINPUT0), .B(G543), .Z(n646) );
  INV_X1 U585 ( .A(G651), .ZN(n536) );
  NOR2_X1 U586 ( .A1(n646), .A2(n536), .ZN(n653) );
  NAND2_X1 U587 ( .A1(G78), .A2(n653), .ZN(n530) );
  NAND2_X1 U588 ( .A1(n531), .A2(n530), .ZN(n535) );
  NOR2_X1 U589 ( .A1(G651), .A2(n646), .ZN(n532) );
  XNOR2_X2 U590 ( .A(KEYINPUT64), .B(n532), .ZN(n659) );
  NAND2_X1 U591 ( .A1(n659), .A2(G53), .ZN(n533) );
  XOR2_X1 U592 ( .A(KEYINPUT68), .B(n533), .Z(n534) );
  NOR2_X1 U593 ( .A1(n535), .A2(n534), .ZN(n539) );
  NOR2_X1 U594 ( .A1(G543), .A2(n536), .ZN(n537) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n537), .Z(n586) );
  NAND2_X1 U596 ( .A1(n586), .A2(G65), .ZN(n538) );
  NAND2_X1 U597 ( .A1(n539), .A2(n538), .ZN(G299) );
  XOR2_X1 U598 ( .A(G2438), .B(G2454), .Z(n541) );
  XNOR2_X1 U599 ( .A(G2435), .B(G2430), .ZN(n540) );
  XNOR2_X1 U600 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U601 ( .A(n542), .B(KEYINPUT102), .Z(n544) );
  XNOR2_X1 U602 ( .A(G1341), .B(G1348), .ZN(n543) );
  XNOR2_X1 U603 ( .A(n544), .B(n543), .ZN(n548) );
  XOR2_X1 U604 ( .A(G2427), .B(G2443), .Z(n546) );
  XNOR2_X1 U605 ( .A(G2451), .B(G2446), .ZN(n545) );
  XNOR2_X1 U606 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U607 ( .A(n548), .B(n547), .Z(n549) );
  AND2_X1 U608 ( .A1(G14), .A2(n549), .ZN(G401) );
  AND2_X1 U609 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U610 ( .A(G132), .ZN(G219) );
  INV_X1 U611 ( .A(G82), .ZN(G220) );
  NAND2_X1 U612 ( .A1(G88), .A2(n655), .ZN(n551) );
  NAND2_X1 U613 ( .A1(G75), .A2(n653), .ZN(n550) );
  NAND2_X1 U614 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U615 ( .A(KEYINPUT82), .B(n552), .ZN(n556) );
  NAND2_X1 U616 ( .A1(G62), .A2(n586), .ZN(n554) );
  NAND2_X1 U617 ( .A1(G50), .A2(n659), .ZN(n553) );
  NAND2_X1 U618 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U619 ( .A1(n556), .A2(n555), .ZN(G166) );
  NAND2_X1 U620 ( .A1(G64), .A2(n586), .ZN(n558) );
  NAND2_X1 U621 ( .A1(G52), .A2(n659), .ZN(n557) );
  NAND2_X1 U622 ( .A1(n558), .A2(n557), .ZN(n563) );
  NAND2_X1 U623 ( .A1(G90), .A2(n655), .ZN(n560) );
  NAND2_X1 U624 ( .A1(G77), .A2(n653), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U626 ( .A(KEYINPUT9), .B(n561), .Z(n562) );
  NOR2_X1 U627 ( .A1(n563), .A2(n562), .ZN(G171) );
  NAND2_X1 U628 ( .A1(G125), .A2(n618), .ZN(n564) );
  XOR2_X1 U629 ( .A(KEYINPUT65), .B(n564), .Z(n567) );
  NAND2_X1 U630 ( .A1(G101), .A2(n898), .ZN(n565) );
  XOR2_X1 U631 ( .A(KEYINPUT23), .B(n565), .Z(n566) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n695) );
  NAND2_X1 U633 ( .A1(G137), .A2(n897), .ZN(n569) );
  NAND2_X1 U634 ( .A1(G113), .A2(n615), .ZN(n568) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n693) );
  NOR2_X1 U636 ( .A1(n695), .A2(n693), .ZN(G160) );
  XNOR2_X1 U637 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n575) );
  NAND2_X1 U638 ( .A1(n655), .A2(G89), .ZN(n570) );
  XNOR2_X1 U639 ( .A(n570), .B(KEYINPUT4), .ZN(n572) );
  NAND2_X1 U640 ( .A1(G76), .A2(n653), .ZN(n571) );
  NAND2_X1 U641 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U642 ( .A(n573), .B(KEYINPUT5), .ZN(n574) );
  XNOR2_X1 U643 ( .A(n575), .B(n574), .ZN(n581) );
  NAND2_X1 U644 ( .A1(n586), .A2(G63), .ZN(n576) );
  XNOR2_X1 U645 ( .A(n576), .B(KEYINPUT74), .ZN(n578) );
  NAND2_X1 U646 ( .A1(G51), .A2(n659), .ZN(n577) );
  NAND2_X1 U647 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U648 ( .A(KEYINPUT6), .B(n579), .ZN(n580) );
  NOR2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U650 ( .A(KEYINPUT7), .B(n582), .Z(G168) );
  XOR2_X1 U651 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U652 ( .A1(G7), .A2(G661), .ZN(n583) );
  XNOR2_X1 U653 ( .A(n583), .B(KEYINPUT70), .ZN(n584) );
  XNOR2_X1 U654 ( .A(KEYINPUT10), .B(n584), .ZN(G223) );
  INV_X1 U655 ( .A(G223), .ZN(n833) );
  NAND2_X1 U656 ( .A1(n833), .A2(G567), .ZN(n585) );
  XOR2_X1 U657 ( .A(KEYINPUT11), .B(n585), .Z(G234) );
  NAND2_X1 U658 ( .A1(G56), .A2(n586), .ZN(n587) );
  XOR2_X1 U659 ( .A(KEYINPUT14), .B(n587), .Z(n594) );
  NAND2_X1 U660 ( .A1(G68), .A2(n653), .ZN(n590) );
  NAND2_X1 U661 ( .A1(n655), .A2(G81), .ZN(n588) );
  XNOR2_X1 U662 ( .A(n588), .B(KEYINPUT12), .ZN(n589) );
  NAND2_X1 U663 ( .A1(n590), .A2(n589), .ZN(n592) );
  XNOR2_X1 U664 ( .A(n592), .B(n591), .ZN(n593) );
  NAND2_X1 U665 ( .A1(G43), .A2(n659), .ZN(n595) );
  INV_X1 U666 ( .A(G860), .ZN(n609) );
  OR2_X1 U667 ( .A1(n966), .A2(n609), .ZN(G153) );
  NAND2_X1 U668 ( .A1(G868), .A2(G171), .ZN(n605) );
  NAND2_X1 U669 ( .A1(G79), .A2(n653), .ZN(n598) );
  NAND2_X1 U670 ( .A1(G54), .A2(n659), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U672 ( .A1(G66), .A2(n586), .ZN(n600) );
  NAND2_X1 U673 ( .A1(G92), .A2(n655), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U675 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X2 U676 ( .A(n603), .B(KEYINPUT15), .ZN(n977) );
  INV_X1 U677 ( .A(n977), .ZN(n627) );
  INV_X1 U678 ( .A(G868), .ZN(n674) );
  NAND2_X1 U679 ( .A1(n627), .A2(n674), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U681 ( .A(n606), .B(KEYINPUT71), .ZN(G284) );
  NOR2_X1 U682 ( .A1(G286), .A2(n674), .ZN(n608) );
  NOR2_X1 U683 ( .A1(G868), .A2(G299), .ZN(n607) );
  NOR2_X1 U684 ( .A1(n608), .A2(n607), .ZN(G297) );
  NAND2_X1 U685 ( .A1(n609), .A2(G559), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n610), .A2(n627), .ZN(n611) );
  XNOR2_X1 U687 ( .A(n611), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U688 ( .A1(G868), .A2(n966), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G868), .A2(n627), .ZN(n612) );
  NOR2_X1 U690 ( .A1(G559), .A2(n612), .ZN(n613) );
  NOR2_X1 U691 ( .A1(n614), .A2(n613), .ZN(G282) );
  BUF_X1 U692 ( .A(n615), .Z(n894) );
  NAND2_X1 U693 ( .A1(n894), .A2(G111), .ZN(n623) );
  NAND2_X1 U694 ( .A1(G135), .A2(n897), .ZN(n617) );
  NAND2_X1 U695 ( .A1(G99), .A2(n898), .ZN(n616) );
  NAND2_X1 U696 ( .A1(n617), .A2(n616), .ZN(n621) );
  BUF_X1 U697 ( .A(n618), .Z(n893) );
  NAND2_X1 U698 ( .A1(n893), .A2(G123), .ZN(n619) );
  XOR2_X1 U699 ( .A(KEYINPUT18), .B(n619), .Z(n620) );
  NOR2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U701 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U702 ( .A(n624), .B(KEYINPUT75), .ZN(n921) );
  XNOR2_X1 U703 ( .A(n921), .B(G2096), .ZN(n626) );
  INV_X1 U704 ( .A(G2100), .ZN(n625) );
  NAND2_X1 U705 ( .A1(n626), .A2(n625), .ZN(G156) );
  XNOR2_X1 U706 ( .A(n966), .B(KEYINPUT76), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n627), .A2(G559), .ZN(n628) );
  XNOR2_X1 U708 ( .A(n629), .B(n628), .ZN(n671) );
  NOR2_X1 U709 ( .A1(G860), .A2(n671), .ZN(n638) );
  NAND2_X1 U710 ( .A1(n655), .A2(G93), .ZN(n630) );
  XOR2_X1 U711 ( .A(KEYINPUT77), .B(n630), .Z(n632) );
  NAND2_X1 U712 ( .A1(n653), .A2(G80), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U714 ( .A(KEYINPUT78), .B(n633), .ZN(n637) );
  NAND2_X1 U715 ( .A1(G67), .A2(n586), .ZN(n635) );
  NAND2_X1 U716 ( .A1(G55), .A2(n659), .ZN(n634) );
  NAND2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U718 ( .A1(n637), .A2(n636), .ZN(n673) );
  XNOR2_X1 U719 ( .A(n638), .B(n673), .ZN(G145) );
  NAND2_X1 U720 ( .A1(G85), .A2(n655), .ZN(n640) );
  NAND2_X1 U721 ( .A1(G72), .A2(n653), .ZN(n639) );
  NAND2_X1 U722 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U723 ( .A1(G60), .A2(n586), .ZN(n641) );
  XNOR2_X1 U724 ( .A(KEYINPUT67), .B(n641), .ZN(n642) );
  NOR2_X1 U725 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U726 ( .A1(G47), .A2(n659), .ZN(n644) );
  NAND2_X1 U727 ( .A1(n645), .A2(n644), .ZN(G290) );
  NAND2_X1 U728 ( .A1(n646), .A2(G87), .ZN(n648) );
  NAND2_X1 U729 ( .A1(G49), .A2(n659), .ZN(n647) );
  NAND2_X1 U730 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U731 ( .A1(n586), .A2(n649), .ZN(n652) );
  NAND2_X1 U732 ( .A1(G74), .A2(G651), .ZN(n650) );
  XOR2_X1 U733 ( .A(KEYINPUT79), .B(n650), .Z(n651) );
  NAND2_X1 U734 ( .A1(n652), .A2(n651), .ZN(G288) );
  NAND2_X1 U735 ( .A1(G73), .A2(n653), .ZN(n654) );
  XNOR2_X1 U736 ( .A(n654), .B(KEYINPUT2), .ZN(n664) );
  NAND2_X1 U737 ( .A1(G61), .A2(n586), .ZN(n657) );
  NAND2_X1 U738 ( .A1(G86), .A2(n655), .ZN(n656) );
  NAND2_X1 U739 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U740 ( .A(KEYINPUT80), .B(n658), .ZN(n662) );
  NAND2_X1 U741 ( .A1(G48), .A2(n659), .ZN(n660) );
  XNOR2_X1 U742 ( .A(KEYINPUT81), .B(n660), .ZN(n661) );
  NOR2_X1 U743 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U744 ( .A1(n664), .A2(n663), .ZN(G305) );
  INV_X1 U745 ( .A(G299), .ZN(n716) );
  XNOR2_X1 U746 ( .A(n716), .B(n673), .ZN(n666) );
  XNOR2_X1 U747 ( .A(G290), .B(G166), .ZN(n665) );
  XNOR2_X1 U748 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U749 ( .A(KEYINPUT19), .B(n667), .ZN(n669) );
  XNOR2_X1 U750 ( .A(G288), .B(KEYINPUT83), .ZN(n668) );
  XNOR2_X1 U751 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U752 ( .A(n670), .B(G305), .ZN(n841) );
  XOR2_X1 U753 ( .A(n841), .B(n671), .Z(n672) );
  NOR2_X1 U754 ( .A1(n674), .A2(n672), .ZN(n676) );
  AND2_X1 U755 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U756 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U757 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XOR2_X1 U758 ( .A(KEYINPUT20), .B(n677), .Z(n678) );
  NAND2_X1 U759 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U760 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U761 ( .A1(n680), .A2(G2072), .ZN(n681) );
  XNOR2_X1 U762 ( .A(KEYINPUT84), .B(n681), .ZN(G158) );
  XNOR2_X1 U763 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U764 ( .A(KEYINPUT69), .B(G57), .ZN(G237) );
  NAND2_X1 U765 ( .A1(G661), .A2(G483), .ZN(n690) );
  NOR2_X1 U766 ( .A1(G220), .A2(G219), .ZN(n682) );
  XNOR2_X1 U767 ( .A(KEYINPUT22), .B(n682), .ZN(n683) );
  NAND2_X1 U768 ( .A1(n683), .A2(G96), .ZN(n684) );
  NOR2_X1 U769 ( .A1(n684), .A2(G218), .ZN(n685) );
  XNOR2_X1 U770 ( .A(n685), .B(KEYINPUT85), .ZN(n839) );
  NAND2_X1 U771 ( .A1(G2106), .A2(n839), .ZN(n689) );
  NAND2_X1 U772 ( .A1(G108), .A2(G120), .ZN(n686) );
  NOR2_X1 U773 ( .A1(G237), .A2(n686), .ZN(n687) );
  NAND2_X1 U774 ( .A1(G69), .A2(n687), .ZN(n838) );
  NAND2_X1 U775 ( .A1(G567), .A2(n838), .ZN(n688) );
  NAND2_X1 U776 ( .A1(n689), .A2(n688), .ZN(n840) );
  NOR2_X1 U777 ( .A1(n690), .A2(n840), .ZN(n691) );
  XNOR2_X1 U778 ( .A(n691), .B(KEYINPUT86), .ZN(n835) );
  NAND2_X1 U779 ( .A1(G36), .A2(n835), .ZN(G176) );
  INV_X1 U780 ( .A(G166), .ZN(G303) );
  INV_X1 U781 ( .A(G171), .ZN(G301) );
  INV_X1 U782 ( .A(G40), .ZN(n692) );
  OR2_X1 U783 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U784 ( .A1(n695), .A2(n694), .ZN(n697) );
  NAND2_X1 U785 ( .A1(G8), .A2(n704), .ZN(n779) );
  INV_X1 U786 ( .A(n704), .ZN(n726) );
  NAND2_X1 U787 ( .A1(n726), .A2(G2072), .ZN(n698) );
  XNOR2_X1 U788 ( .A(n698), .B(KEYINPUT27), .ZN(n700) );
  INV_X1 U789 ( .A(G1956), .ZN(n967) );
  NOR2_X1 U790 ( .A1(n967), .A2(n726), .ZN(n699) );
  NOR2_X1 U791 ( .A1(n700), .A2(n699), .ZN(n717) );
  NOR2_X1 U792 ( .A1(n716), .A2(n717), .ZN(n702) );
  XNOR2_X1 U793 ( .A(KEYINPUT28), .B(KEYINPUT93), .ZN(n701) );
  XNOR2_X1 U794 ( .A(n702), .B(n701), .ZN(n723) );
  XNOR2_X1 U795 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n710) );
  NOR2_X1 U796 ( .A1(G1996), .A2(n710), .ZN(n703) );
  NOR2_X1 U797 ( .A1(n703), .A2(n966), .ZN(n708) );
  NAND2_X1 U798 ( .A1(G1348), .A2(n704), .ZN(n706) );
  NAND2_X1 U799 ( .A1(G2067), .A2(n726), .ZN(n705) );
  NAND2_X1 U800 ( .A1(n706), .A2(n705), .ZN(n718) );
  NAND2_X1 U801 ( .A1(n977), .A2(n718), .ZN(n707) );
  NAND2_X1 U802 ( .A1(n708), .A2(n707), .ZN(n715) );
  INV_X1 U803 ( .A(G1341), .ZN(n996) );
  NAND2_X1 U804 ( .A1(n996), .A2(n710), .ZN(n709) );
  NAND2_X1 U805 ( .A1(n709), .A2(n704), .ZN(n713) );
  AND2_X1 U806 ( .A1(G1996), .A2(n726), .ZN(n711) );
  NAND2_X1 U807 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U809 ( .A1(n715), .A2(n714), .ZN(n721) );
  NAND2_X1 U810 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U811 ( .A1(n719), .A2(n516), .ZN(n720) );
  OR2_X1 U812 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U813 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U814 ( .A(n724), .B(KEYINPUT29), .ZN(n731) );
  XOR2_X1 U815 ( .A(KEYINPUT90), .B(G1961), .Z(n1011) );
  NAND2_X1 U816 ( .A1(n704), .A2(n1011), .ZN(n728) );
  XOR2_X1 U817 ( .A(G2078), .B(KEYINPUT91), .Z(n725) );
  XNOR2_X1 U818 ( .A(KEYINPUT25), .B(n725), .ZN(n952) );
  NAND2_X1 U819 ( .A1(n726), .A2(n952), .ZN(n727) );
  NAND2_X1 U820 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U821 ( .A(n729), .B(KEYINPUT92), .Z(n737) );
  NOR2_X1 U822 ( .A1(G301), .A2(n737), .ZN(n730) );
  XNOR2_X1 U823 ( .A(n732), .B(KEYINPUT95), .ZN(n742) );
  NOR2_X1 U824 ( .A1(G1966), .A2(n779), .ZN(n754) );
  NOR2_X1 U825 ( .A1(G2084), .A2(n704), .ZN(n755) );
  NOR2_X1 U826 ( .A1(n754), .A2(n755), .ZN(n733) );
  XNOR2_X1 U827 ( .A(KEYINPUT96), .B(n733), .ZN(n734) );
  NAND2_X1 U828 ( .A1(n734), .A2(G8), .ZN(n735) );
  XNOR2_X1 U829 ( .A(n735), .B(KEYINPUT30), .ZN(n736) );
  NOR2_X1 U830 ( .A1(G168), .A2(n736), .ZN(n739) );
  AND2_X1 U831 ( .A1(G301), .A2(n737), .ZN(n738) );
  NOR2_X1 U832 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U833 ( .A(KEYINPUT31), .B(n740), .Z(n741) );
  NAND2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n752) );
  NAND2_X1 U835 ( .A1(n752), .A2(G286), .ZN(n749) );
  INV_X1 U836 ( .A(G8), .ZN(n747) );
  NOR2_X1 U837 ( .A1(G1971), .A2(n779), .ZN(n744) );
  NOR2_X1 U838 ( .A1(G2090), .A2(n704), .ZN(n743) );
  NOR2_X1 U839 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U840 ( .A1(G303), .A2(n745), .ZN(n746) );
  OR2_X1 U841 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U842 ( .A(KEYINPUT32), .B(KEYINPUT97), .Z(n750) );
  XNOR2_X1 U843 ( .A(n751), .B(n750), .ZN(n768) );
  INV_X1 U844 ( .A(n752), .ZN(n753) );
  NOR2_X1 U845 ( .A1(n754), .A2(n753), .ZN(n757) );
  NAND2_X1 U846 ( .A1(G8), .A2(n755), .ZN(n756) );
  NAND2_X1 U847 ( .A1(n757), .A2(n756), .ZN(n769) );
  NAND2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n971) );
  AND2_X1 U849 ( .A1(n769), .A2(n971), .ZN(n758) );
  NAND2_X1 U850 ( .A1(n768), .A2(n758), .ZN(n763) );
  INV_X1 U851 ( .A(n971), .ZN(n761) );
  NOR2_X1 U852 ( .A1(G1976), .A2(G288), .ZN(n970) );
  NOR2_X1 U853 ( .A1(G1971), .A2(G303), .ZN(n759) );
  NOR2_X1 U854 ( .A1(n970), .A2(n759), .ZN(n760) );
  OR2_X1 U855 ( .A1(n761), .A2(n760), .ZN(n762) );
  AND2_X1 U856 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U857 ( .A1(n779), .A2(n764), .ZN(n765) );
  XOR2_X1 U858 ( .A(G1981), .B(G305), .Z(n983) );
  NAND2_X1 U859 ( .A1(n970), .A2(KEYINPUT33), .ZN(n766) );
  NAND2_X1 U860 ( .A1(n518), .A2(n767), .ZN(n775) );
  NAND2_X1 U861 ( .A1(n769), .A2(n768), .ZN(n772) );
  NOR2_X1 U862 ( .A1(G2090), .A2(G303), .ZN(n770) );
  NAND2_X1 U863 ( .A1(G8), .A2(n770), .ZN(n771) );
  NAND2_X1 U864 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U865 ( .A1(n773), .A2(n779), .ZN(n774) );
  NAND2_X1 U866 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U867 ( .A(n776), .B(KEYINPUT98), .ZN(n781) );
  NOR2_X1 U868 ( .A1(G1981), .A2(G305), .ZN(n777) );
  XOR2_X1 U869 ( .A(n777), .B(KEYINPUT24), .Z(n778) );
  NOR2_X1 U870 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U872 ( .A(n782), .B(KEYINPUT99), .ZN(n813) );
  NAND2_X1 U873 ( .A1(G131), .A2(n897), .ZN(n784) );
  NAND2_X1 U874 ( .A1(G95), .A2(n898), .ZN(n783) );
  NAND2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n788) );
  NAND2_X1 U876 ( .A1(G119), .A2(n893), .ZN(n786) );
  NAND2_X1 U877 ( .A1(G107), .A2(n894), .ZN(n785) );
  NAND2_X1 U878 ( .A1(n786), .A2(n785), .ZN(n787) );
  OR2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n885) );
  NAND2_X1 U880 ( .A1(G1991), .A2(n885), .ZN(n797) );
  NAND2_X1 U881 ( .A1(G141), .A2(n897), .ZN(n790) );
  NAND2_X1 U882 ( .A1(G117), .A2(n894), .ZN(n789) );
  NAND2_X1 U883 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U884 ( .A1(n898), .A2(G105), .ZN(n791) );
  XOR2_X1 U885 ( .A(KEYINPUT38), .B(n791), .Z(n792) );
  NOR2_X1 U886 ( .A1(n793), .A2(n792), .ZN(n795) );
  NAND2_X1 U887 ( .A1(n893), .A2(G129), .ZN(n794) );
  NAND2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n904) );
  NAND2_X1 U889 ( .A1(G1996), .A2(n904), .ZN(n796) );
  NAND2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U891 ( .A(KEYINPUT88), .B(n798), .Z(n922) );
  NAND2_X1 U892 ( .A1(G160), .A2(G40), .ZN(n799) );
  NOR2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n828) );
  XNOR2_X1 U894 ( .A(KEYINPUT89), .B(n828), .ZN(n801) );
  NOR2_X1 U895 ( .A1(n922), .A2(n801), .ZN(n821) );
  NAND2_X1 U896 ( .A1(G140), .A2(n897), .ZN(n803) );
  NAND2_X1 U897 ( .A1(G104), .A2(n898), .ZN(n802) );
  NAND2_X1 U898 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U899 ( .A(KEYINPUT34), .B(n804), .ZN(n809) );
  NAND2_X1 U900 ( .A1(G128), .A2(n893), .ZN(n806) );
  NAND2_X1 U901 ( .A1(G116), .A2(n894), .ZN(n805) );
  NAND2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U903 ( .A(KEYINPUT35), .B(n807), .Z(n808) );
  NOR2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U905 ( .A(KEYINPUT36), .B(n810), .ZN(n891) );
  XNOR2_X1 U906 ( .A(KEYINPUT37), .B(G2067), .ZN(n826) );
  NOR2_X1 U907 ( .A1(n891), .A2(n826), .ZN(n918) );
  NAND2_X1 U908 ( .A1(n828), .A2(n918), .ZN(n824) );
  NAND2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n815) );
  XNOR2_X1 U910 ( .A(G1986), .B(G290), .ZN(n979) );
  NAND2_X1 U911 ( .A1(n979), .A2(n828), .ZN(n816) );
  NAND2_X1 U912 ( .A1(n817), .A2(n816), .ZN(n831) );
  NOR2_X1 U913 ( .A1(G1996), .A2(n904), .ZN(n934) );
  NOR2_X1 U914 ( .A1(G1991), .A2(n885), .ZN(n925) );
  NOR2_X1 U915 ( .A1(G1986), .A2(G290), .ZN(n818) );
  XOR2_X1 U916 ( .A(n818), .B(KEYINPUT101), .Z(n819) );
  NOR2_X1 U917 ( .A1(n925), .A2(n819), .ZN(n820) );
  NOR2_X1 U918 ( .A1(n821), .A2(n820), .ZN(n822) );
  NOR2_X1 U919 ( .A1(n934), .A2(n822), .ZN(n823) );
  XNOR2_X1 U920 ( .A(n823), .B(KEYINPUT39), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n891), .A2(n826), .ZN(n917) );
  NAND2_X1 U923 ( .A1(n827), .A2(n917), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U926 ( .A(n832), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U929 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U931 ( .A1(n836), .A2(n835), .ZN(n837) );
  XOR2_X1 U932 ( .A(KEYINPUT103), .B(n837), .Z(G188) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G108), .ZN(G238) );
  INV_X1 U936 ( .A(G96), .ZN(G221) );
  INV_X1 U937 ( .A(G69), .ZN(G235) );
  NOR2_X1 U938 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  XOR2_X1 U940 ( .A(KEYINPUT104), .B(n840), .Z(G319) );
  XOR2_X1 U941 ( .A(KEYINPUT112), .B(n841), .Z(n843) );
  XNOR2_X1 U942 ( .A(G171), .B(G286), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n844), .B(n977), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n845), .B(n966), .ZN(n846) );
  NOR2_X1 U946 ( .A1(G37), .A2(n846), .ZN(G397) );
  XOR2_X1 U947 ( .A(G1971), .B(G1956), .Z(n848) );
  XNOR2_X1 U948 ( .A(G1981), .B(G1966), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(n858) );
  XOR2_X1 U950 ( .A(KEYINPUT41), .B(G2474), .Z(n850) );
  XNOR2_X1 U951 ( .A(G1996), .B(KEYINPUT107), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U953 ( .A(G1976), .B(G1961), .Z(n852) );
  XNOR2_X1 U954 ( .A(G1991), .B(G1986), .ZN(n851) );
  XNOR2_X1 U955 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U956 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U957 ( .A(KEYINPUT109), .B(KEYINPUT108), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U959 ( .A(n858), .B(n857), .Z(G229) );
  XOR2_X1 U960 ( .A(G2100), .B(KEYINPUT106), .Z(n860) );
  XNOR2_X1 U961 ( .A(KEYINPUT105), .B(KEYINPUT43), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U963 ( .A(KEYINPUT42), .B(G2072), .Z(n862) );
  XNOR2_X1 U964 ( .A(G2067), .B(G2090), .ZN(n861) );
  XNOR2_X1 U965 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U966 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U967 ( .A(G2678), .B(G2096), .ZN(n865) );
  XNOR2_X1 U968 ( .A(n866), .B(n865), .ZN(n868) );
  XOR2_X1 U969 ( .A(G2078), .B(G2084), .Z(n867) );
  XNOR2_X1 U970 ( .A(n868), .B(n867), .ZN(G227) );
  NAND2_X1 U971 ( .A1(n893), .A2(G124), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n869), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U973 ( .A1(G136), .A2(n897), .ZN(n870) );
  NAND2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U975 ( .A(KEYINPUT110), .B(n872), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G100), .A2(n898), .ZN(n874) );
  NAND2_X1 U977 ( .A1(G112), .A2(n894), .ZN(n873) );
  NAND2_X1 U978 ( .A1(n874), .A2(n873), .ZN(n875) );
  NOR2_X1 U979 ( .A1(n876), .A2(n875), .ZN(G162) );
  XNOR2_X1 U980 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n887) );
  NAND2_X1 U981 ( .A1(G139), .A2(n897), .ZN(n878) );
  NAND2_X1 U982 ( .A1(G103), .A2(n898), .ZN(n877) );
  NAND2_X1 U983 ( .A1(n878), .A2(n877), .ZN(n884) );
  NAND2_X1 U984 ( .A1(G127), .A2(n893), .ZN(n880) );
  NAND2_X1 U985 ( .A1(G115), .A2(n894), .ZN(n879) );
  NAND2_X1 U986 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U987 ( .A(KEYINPUT111), .B(n881), .ZN(n882) );
  XNOR2_X1 U988 ( .A(KEYINPUT47), .B(n882), .ZN(n883) );
  NOR2_X1 U989 ( .A1(n884), .A2(n883), .ZN(n928) );
  XNOR2_X1 U990 ( .A(n885), .B(n928), .ZN(n886) );
  XNOR2_X1 U991 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U992 ( .A(n888), .B(n921), .Z(n890) );
  XNOR2_X1 U993 ( .A(G160), .B(G162), .ZN(n889) );
  XNOR2_X1 U994 ( .A(n890), .B(n889), .ZN(n892) );
  XNOR2_X1 U995 ( .A(n892), .B(n891), .ZN(n908) );
  NAND2_X1 U996 ( .A1(G130), .A2(n893), .ZN(n896) );
  NAND2_X1 U997 ( .A1(G118), .A2(n894), .ZN(n895) );
  NAND2_X1 U998 ( .A1(n896), .A2(n895), .ZN(n903) );
  NAND2_X1 U999 ( .A1(G142), .A2(n897), .ZN(n900) );
  NAND2_X1 U1000 ( .A1(G106), .A2(n898), .ZN(n899) );
  NAND2_X1 U1001 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U1002 ( .A(n901), .B(KEYINPUT45), .Z(n902) );
  NOR2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1005 ( .A(G164), .B(n906), .Z(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n909), .ZN(G395) );
  INV_X1 U1008 ( .A(G319), .ZN(n910) );
  NOR2_X1 U1009 ( .A1(n910), .A2(G401), .ZN(n914) );
  NOR2_X1 U1010 ( .A1(G229), .A2(G227), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n911), .ZN(n912) );
  NOR2_X1 U1012 ( .A1(G397), .A2(n912), .ZN(n913) );
  NAND2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1014 ( .A1(n915), .A2(G395), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(n916), .B(KEYINPUT113), .ZN(G225) );
  XOR2_X1 U1016 ( .A(KEYINPUT114), .B(G225), .Z(G308) );
  INV_X1 U1017 ( .A(n917), .ZN(n919) );
  NOR2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n927) );
  XOR2_X1 U1019 ( .A(G2084), .B(G160), .Z(n920) );
  NOR2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n923) );
  NAND2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n939) );
  XNOR2_X1 U1024 ( .A(G2072), .B(n928), .ZN(n930) );
  XNOR2_X1 U1025 ( .A(G164), .B(G2078), .ZN(n929) );
  NAND2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(n931), .B(KEYINPUT50), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(n932), .B(KEYINPUT115), .ZN(n937) );
  XOR2_X1 U1029 ( .A(G2090), .B(G162), .Z(n933) );
  NOR2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1031 ( .A(KEYINPUT51), .B(n935), .Z(n936) );
  NAND2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1034 ( .A(KEYINPUT52), .B(n940), .ZN(n941) );
  XOR2_X1 U1035 ( .A(KEYINPUT55), .B(KEYINPUT116), .Z(n943) );
  NAND2_X1 U1036 ( .A1(n941), .A2(n943), .ZN(n942) );
  NAND2_X1 U1037 ( .A1(n942), .A2(G29), .ZN(n1027) );
  INV_X1 U1038 ( .A(G29), .ZN(n963) );
  XOR2_X1 U1039 ( .A(n943), .B(KEYINPUT117), .Z(n961) );
  XOR2_X1 U1040 ( .A(G2084), .B(G34), .Z(n944) );
  XNOR2_X1 U1041 ( .A(KEYINPUT54), .B(n944), .ZN(n959) );
  XNOR2_X1 U1042 ( .A(G2090), .B(G35), .ZN(n957) );
  XNOR2_X1 U1043 ( .A(G1996), .B(G32), .ZN(n946) );
  XNOR2_X1 U1044 ( .A(G33), .B(G2072), .ZN(n945) );
  NOR2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n951) );
  XOR2_X1 U1046 ( .A(G1991), .B(G25), .Z(n947) );
  NAND2_X1 U1047 ( .A1(n947), .A2(G28), .ZN(n949) );
  XNOR2_X1 U1048 ( .A(G26), .B(G2067), .ZN(n948) );
  NOR2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n954) );
  XOR2_X1 U1051 ( .A(G27), .B(n952), .Z(n953) );
  NOR2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1053 ( .A(KEYINPUT53), .B(n955), .ZN(n956) );
  NOR2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(n961), .B(n960), .ZN(n962) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n964), .A2(G11), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(n965), .B(KEYINPUT118), .ZN(n1025) );
  XNOR2_X1 U1060 ( .A(n996), .B(n966), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(G299), .B(n967), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n991) );
  XNOR2_X1 U1063 ( .A(G166), .B(G1971), .ZN(n975) );
  INV_X1 U1064 ( .A(n970), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1066 ( .A(KEYINPUT120), .B(n973), .Z(n974) );
  NAND2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1068 ( .A(n976), .B(KEYINPUT121), .ZN(n989) );
  XNOR2_X1 U1069 ( .A(G1348), .B(n977), .ZN(n978) );
  NOR2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n982) );
  XNOR2_X1 U1071 ( .A(G1961), .B(KEYINPUT119), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(n980), .B(G301), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n987) );
  XNOR2_X1 U1074 ( .A(G1966), .B(G168), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1076 ( .A(KEYINPUT57), .B(n985), .Z(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n993) );
  XOR2_X1 U1080 ( .A(G16), .B(KEYINPUT56), .Z(n992) );
  NOR2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n1022) );
  XOR2_X1 U1082 ( .A(G4), .B(KEYINPUT122), .Z(n995) );
  XNOR2_X1 U1083 ( .A(G1348), .B(KEYINPUT59), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(n995), .B(n994), .ZN(n1002) );
  XNOR2_X1 U1085 ( .A(G19), .B(n996), .ZN(n1000) );
  XNOR2_X1 U1086 ( .A(G1981), .B(G6), .ZN(n998) );
  XNOR2_X1 U1087 ( .A(G1956), .B(G20), .ZN(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(KEYINPUT60), .B(KEYINPUT123), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(n1004), .B(n1003), .ZN(n1017) );
  XNOR2_X1 U1093 ( .A(G1971), .B(G22), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(G23), .B(G1976), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  XOR2_X1 U1096 ( .A(G1986), .B(G24), .Z(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1010) );
  XOR2_X1 U1098 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n1009) );
  XNOR2_X1 U1099 ( .A(n1010), .B(n1009), .ZN(n1015) );
  XOR2_X1 U1100 ( .A(n1011), .B(G5), .Z(n1013) );
  XNOR2_X1 U1101 ( .A(G21), .B(G1966), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(KEYINPUT61), .B(KEYINPUT125), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(n1019), .B(n1018), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(G16), .A2(n1020), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1109 ( .A(KEYINPUT126), .B(n1023), .Z(n1024) );
  NOR2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(n1028), .B(KEYINPUT62), .ZN(n1029) );
  XNOR2_X1 U1113 ( .A(KEYINPUT127), .B(n1029), .ZN(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

