//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  AND2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(G353));
  NOR2_X1   g0007(.A1(G97), .A2(G107), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(new_n212), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(KEYINPUT65), .B(G77), .Z(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  AND2_X1   g0024(.A1(new_n224), .A2(G244), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G50), .A2(G226), .ZN(new_n229));
  NAND4_X1  g0029(.A1(new_n226), .A2(new_n227), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n214), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n217), .B(new_n222), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT66), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G169), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(new_n220), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  OAI211_X1 g0056(.A(G232), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT75), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT3), .B(G33), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT75), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n259), .A2(new_n260), .A3(G232), .A4(G1698), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G97), .ZN(new_n262));
  AND3_X1   g0062(.A1(new_n258), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  OAI211_X1 g0064(.A(G226), .B(new_n264), .C1(new_n255), .C2(new_n256), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT74), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n259), .A2(KEYINPUT74), .A3(G226), .A4(new_n264), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n254), .B1(new_n263), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT68), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(new_n252), .B2(new_n220), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n251), .A2(KEYINPUT68), .A3(G1), .A4(G13), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n272), .A2(new_n273), .A3(G238), .A4(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n211), .A2(G274), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(new_n271), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT67), .B(G41), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n277), .B1(new_n278), .B2(G45), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(KEYINPUT13), .B1(new_n270), .B2(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n267), .A2(new_n268), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n258), .A2(new_n261), .A3(new_n262), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n253), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT13), .ZN(new_n285));
  INV_X1    g0085(.A(new_n280), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n250), .B1(new_n281), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT14), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(KEYINPUT78), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n288), .B(new_n290), .ZN(new_n291));
  AND3_X1   g0091(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n285), .B1(new_n284), .B2(new_n286), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  NOR3_X1   g0094(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(KEYINPUT78), .B2(new_n289), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT71), .ZN(new_n298));
  NAND4_X1  g0098(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n299), .A2(new_n220), .ZN(new_n300));
  NAND3_X1  g0100(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT69), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(KEYINPUT70), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  AND4_X1   g0104(.A1(KEYINPUT70), .A2(new_n303), .A3(new_n220), .A4(new_n299), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n298), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n303), .A2(new_n220), .A3(new_n299), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT70), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n303), .A2(KEYINPUT70), .A3(new_n220), .A4(new_n299), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n309), .A2(KEYINPUT71), .A3(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(G20), .A2(G33), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n312), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n212), .A2(G33), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n313), .B1(new_n206), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n306), .A2(new_n311), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT11), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n306), .A2(KEYINPUT11), .A3(new_n311), .A4(new_n315), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(G68), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n321), .B(KEYINPUT12), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n212), .A2(G1), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(new_n309), .B2(new_n310), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n322), .B1(new_n324), .B2(G68), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n318), .A2(new_n319), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n297), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n272), .A2(new_n273), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n329), .A2(new_n274), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G244), .ZN(new_n331));
  OR2_X1    g0131(.A1(KEYINPUT3), .A2(G33), .ZN(new_n332));
  NAND2_X1  g0132(.A1(KEYINPUT3), .A2(G33), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n264), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n255), .A2(new_n256), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n334), .A2(G238), .B1(new_n335), .B2(G107), .ZN(new_n336));
  INV_X1    g0136(.A(G232), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n259), .A2(new_n264), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n253), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n331), .A2(new_n279), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n250), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n324), .A2(G77), .ZN(new_n343));
  XOR2_X1   g0143(.A(KEYINPUT8), .B(G58), .Z(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n312), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT15), .B(G87), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n345), .B1(new_n314), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(G20), .B2(new_n224), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n309), .A2(new_n310), .ZN(new_n349));
  OAI221_X1 g0149(.A(new_n343), .B1(new_n224), .B2(new_n320), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n342), .B(new_n350), .C1(G179), .C2(new_n341), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n341), .A2(G200), .ZN(new_n352));
  INV_X1    g0152(.A(G190), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n352), .B1(new_n353), .B2(new_n341), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n354), .A2(new_n350), .ZN(new_n355));
  AND3_X1   g0155(.A1(new_n327), .A2(new_n351), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n306), .A2(new_n311), .ZN(new_n357));
  INV_X1    g0157(.A(new_n323), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n357), .A2(new_n344), .A3(new_n320), .A4(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n344), .ZN(new_n360));
  INV_X1    g0160(.A(new_n320), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT7), .B1(new_n259), .B2(G20), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT7), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n335), .A2(new_n365), .A3(new_n212), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(new_n366), .A3(G68), .ZN(new_n367));
  XNOR2_X1  g0167(.A(G58), .B(G68), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n368), .A2(G20), .B1(G159), .B2(new_n312), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT16), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n367), .A2(KEYINPUT16), .A3(new_n369), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n304), .A2(new_n305), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n363), .A2(new_n377), .A3(KEYINPUT79), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n359), .B(new_n362), .C1(new_n349), .C2(new_n374), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT79), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n272), .A2(new_n273), .A3(G232), .A4(new_n274), .ZN(new_n382));
  MUX2_X1   g0182(.A(G223), .B(G226), .S(G1698), .Z(new_n383));
  AOI22_X1  g0183(.A1(new_n383), .A2(new_n259), .B1(G33), .B2(G87), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n382), .B(new_n279), .C1(new_n384), .C2(new_n254), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n385), .A2(new_n294), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(G169), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT80), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n386), .A2(KEYINPUT80), .A3(new_n387), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n378), .A2(new_n381), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT18), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT17), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n385), .A2(new_n353), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(G200), .B2(new_n385), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n395), .B1(new_n379), .B2(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n363), .A2(new_n377), .A3(KEYINPUT17), .A4(new_n397), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT18), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n378), .A2(new_n381), .A3(new_n392), .A4(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n394), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT76), .ZN(new_n406));
  INV_X1    g0206(.A(G200), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n292), .B2(new_n293), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n281), .A2(new_n353), .A3(new_n287), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n326), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n406), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI211_X1 g0212(.A(KEYINPUT76), .B(new_n326), .C1(new_n408), .C2(new_n409), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT77), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NOR3_X1   g0215(.A1(new_n292), .A2(new_n293), .A3(G190), .ZN(new_n416));
  AOI21_X1  g0216(.A(G200), .B1(new_n281), .B2(new_n287), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n411), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT76), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n410), .A2(new_n406), .A3(new_n411), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT77), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n356), .B(new_n405), .C1(new_n415), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n330), .A2(G226), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n279), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n224), .A2(new_n335), .B1(G223), .B2(new_n334), .ZN(new_n425));
  INV_X1    g0225(.A(G222), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n425), .B1(new_n426), .B2(new_n338), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n424), .B1(new_n253), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n294), .ZN(new_n429));
  XOR2_X1   g0229(.A(new_n429), .B(KEYINPUT73), .Z(new_n430));
  INV_X1    g0230(.A(new_n357), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n312), .A2(G150), .ZN(new_n432));
  OAI221_X1 g0232(.A(new_n432), .B1(new_n360), .B2(new_n314), .C1(new_n205), .C2(new_n212), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n357), .A2(G50), .A3(new_n320), .A4(new_n358), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n361), .A2(new_n201), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n435), .A2(KEYINPUT72), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT72), .B1(new_n435), .B2(new_n436), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n434), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n430), .B(new_n439), .C1(G169), .C2(new_n428), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(KEYINPUT9), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT9), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n442), .B(new_n434), .C1(new_n437), .C2(new_n438), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT10), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n428), .A2(new_n407), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n446), .B1(G190), .B2(new_n428), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n444), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n445), .B1(new_n444), .B2(new_n447), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n440), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n422), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n334), .A2(G264), .ZN(new_n452));
  INV_X1    g0252(.A(G303), .ZN(new_n453));
  INV_X1    g0253(.A(G257), .ZN(new_n454));
  OAI221_X1 g0254(.A(new_n452), .B1(new_n453), .B2(new_n259), .C1(new_n454), .C2(new_n338), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n253), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT5), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n211), .B(G45), .C1(new_n457), .C2(G41), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n458), .B1(new_n278), .B2(new_n457), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n459), .A2(G274), .A3(new_n272), .A4(new_n273), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G270), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n328), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT84), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT84), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n328), .A2(new_n459), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G270), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n465), .B1(new_n467), .B2(new_n460), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n456), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(G20), .B1(G33), .B2(G283), .ZN(new_n470));
  INV_X1    g0270(.A(G33), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G97), .ZN(new_n472));
  INV_X1    g0272(.A(G116), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n470), .A2(new_n472), .B1(G20), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n307), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT20), .ZN(new_n476));
  XNOR2_X1  g0276(.A(new_n475), .B(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n471), .A2(G1), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n349), .A2(G116), .A3(new_n320), .A4(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n320), .A2(G116), .ZN(new_n481));
  XNOR2_X1  g0281(.A(new_n481), .B(KEYINPUT85), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n477), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n469), .A2(KEYINPUT21), .A3(G169), .A4(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT21), .ZN(new_n485));
  OAI21_X1  g0285(.A(KEYINPUT84), .B1(new_n461), .B2(new_n463), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n467), .A2(new_n465), .A3(new_n460), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n486), .A2(new_n487), .B1(new_n253), .B2(new_n455), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n483), .A2(G169), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(G179), .A3(new_n483), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n484), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(G190), .B(new_n456), .C1(new_n464), .C2(new_n468), .ZN(new_n493));
  INV_X1    g0293(.A(new_n483), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n493), .B(new_n494), .C1(new_n488), .C2(new_n407), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n458), .ZN(new_n498));
  AND2_X1   g0298(.A1(KEYINPUT67), .A2(G41), .ZN(new_n499));
  NOR2_X1   g0299(.A1(KEYINPUT67), .A2(G41), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n457), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n502), .A2(G264), .A3(new_n272), .A4(new_n273), .ZN(new_n503));
  OAI211_X1 g0303(.A(G250), .B(new_n264), .C1(new_n255), .C2(new_n256), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G294), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT87), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n334), .A2(new_n507), .A3(G257), .ZN(new_n508));
  OAI211_X1 g0308(.A(G257), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT87), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n506), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n503), .B(new_n460), .C1(new_n511), .C2(new_n254), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(new_n353), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n513), .B1(G200), .B2(new_n512), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n357), .A2(G107), .A3(new_n320), .A4(new_n479), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n212), .B(G87), .C1(new_n255), .C2(new_n256), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT22), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT22), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n259), .A2(new_n518), .A3(new_n212), .A4(G87), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT24), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n471), .A2(new_n473), .A3(G20), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT23), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n212), .B2(G107), .ZN(new_n524));
  INV_X1    g0324(.A(G107), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(KEYINPUT23), .A3(G20), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n522), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n520), .A2(new_n521), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n521), .B1(new_n520), .B2(new_n527), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n376), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n361), .A2(KEYINPUT25), .A3(new_n525), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT86), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT25), .B1(new_n361), .B2(new_n525), .ZN(new_n533));
  XOR2_X1   g0333(.A(new_n532), .B(new_n533), .Z(new_n534));
  NAND3_X1  g0334(.A1(new_n515), .A2(new_n530), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n514), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT88), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n512), .A2(new_n538), .A3(G169), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n508), .A2(new_n510), .ZN(new_n540));
  INV_X1    g0340(.A(new_n506), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n253), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n543), .A2(G179), .A3(new_n460), .A4(new_n503), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n538), .B1(new_n512), .B2(G169), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n535), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n537), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n320), .A2(G97), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT6), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT81), .ZN(new_n551));
  INV_X1    g0351(.A(G97), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT6), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G97), .A2(G107), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n209), .A2(new_n551), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  AND2_X1   g0355(.A1(G97), .A2(G107), .ZN(new_n556));
  OAI211_X1 g0356(.A(KEYINPUT81), .B(new_n550), .C1(new_n556), .C2(new_n208), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G20), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n364), .A2(new_n366), .A3(G107), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n312), .A2(G77), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n549), .B1(new_n562), .B2(new_n376), .ZN(new_n563));
  AND3_X1   g0363(.A1(new_n309), .A2(KEYINPUT71), .A3(new_n310), .ZN(new_n564));
  AOI21_X1  g0364(.A(KEYINPUT71), .B1(new_n309), .B2(new_n310), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n320), .B(new_n479), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n563), .B1(new_n566), .B2(new_n552), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(G274), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n328), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n466), .A2(G257), .B1(new_n570), .B2(new_n459), .ZN(new_n571));
  OAI211_X1 g0371(.A(G244), .B(new_n264), .C1(new_n255), .C2(new_n256), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT4), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n259), .A2(KEYINPUT4), .A3(G244), .A4(new_n264), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G33), .A2(G283), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n259), .A2(G250), .A3(G1698), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n574), .A2(new_n575), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n578), .A2(KEYINPUT82), .A3(new_n253), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT82), .B1(new_n578), .B2(new_n253), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n571), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G200), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n578), .A2(new_n253), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n329), .A2(G257), .A3(new_n502), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n583), .A2(G190), .A3(new_n460), .A4(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT83), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n571), .A2(KEYINPUT83), .A3(G190), .A4(new_n583), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n568), .A2(new_n582), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n259), .A2(new_n212), .A3(G68), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT19), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n212), .B1(new_n262), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(G87), .B2(new_n209), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n591), .B1(new_n314), .B2(new_n552), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n590), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n376), .A2(new_n595), .B1(new_n361), .B2(new_n346), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  AOI211_X1 g0397(.A(new_n361), .B(new_n478), .C1(new_n306), .C2(new_n311), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n597), .B1(new_n598), .B2(G87), .ZN(new_n599));
  OAI211_X1 g0399(.A(G238), .B(new_n264), .C1(new_n255), .C2(new_n256), .ZN(new_n600));
  OAI211_X1 g0400(.A(G244), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n600), .B(new_n601), .C1(new_n471), .C2(new_n473), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n253), .ZN(new_n603));
  INV_X1    g0403(.A(G45), .ZN(new_n604));
  OAI21_X1  g0404(.A(G250), .B1(new_n604), .B2(G1), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n604), .B2(new_n276), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n329), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n407), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n603), .A2(new_n607), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n608), .B1(new_n610), .B2(G190), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n596), .B1(new_n566), .B2(new_n346), .ZN(new_n612));
  AOI21_X1  g0412(.A(G169), .B1(new_n603), .B2(new_n607), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(new_n610), .B2(new_n294), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n599), .A2(new_n611), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n571), .A2(new_n583), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n250), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n294), .B(new_n571), .C1(new_n579), .C2(new_n580), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n567), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n589), .A2(new_n615), .A3(new_n619), .ZN(new_n620));
  AND4_X1   g0420(.A1(new_n451), .A2(new_n497), .A3(new_n548), .A4(new_n620), .ZN(G372));
  AND3_X1   g0421(.A1(new_n567), .A2(new_n617), .A3(new_n618), .ZN(new_n622));
  INV_X1    g0422(.A(new_n580), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n578), .A2(KEYINPUT82), .A3(new_n253), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n407), .B1(new_n625), .B2(new_n571), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n587), .A2(new_n588), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n622), .B1(new_n628), .B2(new_n568), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n547), .A2(new_n484), .A3(new_n490), .A4(new_n491), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n514), .A2(new_n536), .B1(new_n599), .B2(new_n611), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n612), .A2(new_n614), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n610), .A2(G190), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n357), .A2(G87), .A3(new_n320), .A4(new_n479), .ZN(new_n635));
  INV_X1    g0435(.A(new_n608), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n634), .A2(new_n635), .A3(new_n596), .A4(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(KEYINPUT26), .B1(new_n638), .B2(new_n619), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n632), .A2(new_n633), .A3(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT89), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n638), .B1(new_n641), .B2(new_n619), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n567), .A2(new_n617), .A3(new_n618), .A4(KEYINPUT89), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n451), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n440), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n327), .A2(new_n351), .ZN(new_n649));
  INV_X1    g0449(.A(new_n327), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n419), .A2(new_n420), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n649), .B(new_n401), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n379), .A2(new_n388), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(KEYINPUT18), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n379), .A2(new_n402), .A3(new_n388), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n448), .A2(new_n449), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n648), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n647), .A2(new_n659), .ZN(G369));
  NAND3_X1  g0460(.A1(new_n211), .A2(new_n212), .A3(G13), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  XOR2_X1   g0462(.A(new_n662), .B(KEYINPUT90), .Z(new_n663));
  INV_X1    g0463(.A(G213), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(new_n661), .B2(KEYINPUT27), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(new_n494), .ZN(new_n670));
  MUX2_X1   g0470(.A(new_n497), .B(new_n492), .S(new_n670), .Z(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G330), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n548), .B1(new_n536), .B2(new_n669), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n547), .B2(new_n669), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n492), .A2(new_n669), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n548), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n547), .A2(new_n668), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n676), .A2(new_n681), .ZN(G399));
  INV_X1    g0482(.A(new_n215), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(new_n278), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n209), .A2(G87), .A3(G116), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G1), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n218), .B2(new_n685), .ZN(new_n688));
  XOR2_X1   g0488(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n689));
  XNOR2_X1  g0489(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n646), .A2(KEYINPUT93), .A3(new_n669), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT29), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n669), .B1(new_n640), .B2(new_n645), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT93), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n691), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT94), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n642), .A2(new_n697), .A3(KEYINPUT26), .A4(new_n644), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n619), .A2(new_n641), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n699), .A2(new_n615), .A3(KEYINPUT26), .A4(new_n644), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n643), .B1(new_n638), .B2(new_n619), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(KEYINPUT94), .A3(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n698), .A2(new_n702), .A3(new_n633), .A4(new_n632), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(KEYINPUT29), .A3(new_n669), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n696), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(G330), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT31), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n497), .A2(new_n620), .A3(new_n548), .A4(new_n669), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n488), .A2(G179), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n542), .A2(new_n253), .B1(new_n466), .B2(G264), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(new_n610), .A3(new_n571), .A4(new_n583), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT92), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT30), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  OAI211_X1 g0514(.A(KEYINPUT92), .B(new_n714), .C1(new_n709), .C2(new_n711), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n610), .A2(G179), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n469), .A2(new_n512), .A3(new_n581), .A4(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n713), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n668), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n707), .B1(new_n708), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(KEYINPUT31), .B1(new_n718), .B2(new_n668), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n706), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n705), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n690), .B1(new_n727), .B2(G1), .ZN(G364));
  AND2_X1   g0528(.A1(new_n212), .A2(G13), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n211), .B1(new_n729), .B2(G45), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n684), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n673), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(G330), .B2(new_n671), .ZN(new_n734));
  INV_X1    g0534(.A(new_n732), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n220), .B1(G20), .B2(new_n250), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n212), .A2(G190), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n739), .A2(new_n294), .A3(G200), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n741), .A2(KEYINPUT96), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(KEYINPUT96), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n224), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G179), .A2(G200), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT97), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n739), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G159), .ZN(new_n750));
  XOR2_X1   g0550(.A(new_n750), .B(KEYINPUT32), .Z(new_n751));
  OAI21_X1  g0551(.A(G20), .B1(new_n748), .B2(new_n353), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G97), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n212), .A2(new_n353), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n407), .A2(G179), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n757), .A2(G87), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n754), .A2(G179), .A3(new_n407), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n294), .A2(new_n407), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(new_n738), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n759), .A2(new_n202), .B1(new_n761), .B2(new_n203), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n738), .A2(new_n755), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n259), .B1(new_n763), .B2(new_n525), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n754), .A2(new_n760), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n201), .ZN(new_n766));
  NOR4_X1   g0566(.A1(new_n758), .A2(new_n762), .A3(new_n764), .A4(new_n766), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n746), .A2(new_n751), .A3(new_n753), .A4(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G326), .ZN(new_n769));
  INV_X1    g0569(.A(G283), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n765), .A2(new_n769), .B1(new_n763), .B2(new_n770), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n259), .B(new_n771), .C1(G311), .C2(new_n740), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n756), .A2(new_n453), .ZN(new_n773));
  INV_X1    g0573(.A(G317), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n774), .A2(KEYINPUT33), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(KEYINPUT33), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n761), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n759), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n773), .B(new_n777), .C1(G322), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n752), .A2(G294), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n749), .A2(G329), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n772), .A2(new_n779), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n737), .B1(new_n768), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G13), .A2(G33), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n736), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n215), .A2(new_n259), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT95), .Z(new_n789));
  INV_X1    g0589(.A(G355), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n789), .A2(new_n790), .B1(G116), .B2(new_n215), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n683), .A2(new_n259), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(G45), .B2(new_n218), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(G45), .B2(new_n248), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n735), .B(new_n783), .C1(new_n787), .C2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n786), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n796), .B1(new_n671), .B2(new_n797), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n734), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(G396));
  NOR2_X1   g0600(.A1(new_n351), .A2(new_n668), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n350), .A2(new_n668), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n802), .A2(KEYINPUT100), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(KEYINPUT100), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n355), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n801), .B1(new_n805), .B2(new_n351), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n691), .A2(new_n695), .A3(new_n807), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n808), .A2(KEYINPUT101), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(KEYINPUT101), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n806), .B(new_n669), .C1(new_n640), .C2(new_n645), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n732), .B1(new_n812), .B2(new_n725), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n725), .B2(new_n812), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n736), .A2(new_n784), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n735), .B1(new_n206), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n765), .ZN(new_n817));
  INV_X1    g0617(.A(new_n763), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n817), .A2(G303), .B1(new_n818), .B2(G87), .ZN(new_n819));
  INV_X1    g0619(.A(G294), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n819), .B1(new_n770), .B2(new_n761), .C1(new_n820), .C2(new_n759), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n259), .B(new_n821), .C1(G107), .C2(new_n757), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n745), .A2(G116), .B1(G311), .B2(new_n749), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n822), .A2(new_n753), .A3(new_n823), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT98), .Z(new_n825));
  OAI21_X1  g0625(.A(new_n259), .B1(new_n756), .B2(new_n201), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(G68), .B2(new_n818), .ZN(new_n827));
  INV_X1    g0627(.A(new_n749), .ZN(new_n828));
  INV_X1    g0628(.A(G132), .ZN(new_n829));
  INV_X1    g0629(.A(new_n752), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n827), .B1(new_n828), .B2(new_n829), .C1(new_n202), .C2(new_n830), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n778), .A2(G143), .B1(new_n817), .B2(G137), .ZN(new_n832));
  INV_X1    g0632(.A(G150), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(new_n761), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n745), .B2(G159), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n831), .B1(new_n835), .B2(KEYINPUT34), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(KEYINPUT34), .B2(new_n835), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n825), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(KEYINPUT99), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n736), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n838), .A2(KEYINPUT99), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n816), .B1(new_n785), .B2(new_n806), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n814), .A2(new_n842), .ZN(G384));
  OAI211_X1 g0643(.A(G116), .B(new_n221), .C1(new_n558), .C2(KEYINPUT35), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT102), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n558), .A2(KEYINPUT35), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(KEYINPUT103), .B(KEYINPUT36), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n849), .B(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n224), .B(new_n219), .C1(new_n202), .C2(new_n203), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n201), .A2(G68), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n211), .B(G13), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n451), .A2(new_n724), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n411), .A2(new_n669), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n327), .A2(new_n651), .A3(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT104), .ZN(new_n860));
  INV_X1    g0660(.A(new_n297), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n415), .B2(new_n421), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n860), .B1(new_n862), .B2(new_n857), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n414), .B1(new_n412), .B2(new_n413), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n419), .A2(KEYINPUT77), .A3(new_n420), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n297), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n866), .A2(KEYINPUT104), .A3(new_n858), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n859), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n666), .B(KEYINPUT105), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n378), .A2(new_n381), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n653), .B1(new_n379), .B2(new_n398), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT37), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n379), .A2(new_n398), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n378), .A2(new_n381), .A3(new_n869), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n393), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n401), .A2(new_n654), .A3(new_n655), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n870), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n359), .A2(new_n362), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n431), .B2(new_n375), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n884), .A2(new_n666), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n404), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n666), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n388), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT37), .B1(new_n889), .B2(new_n873), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n876), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n886), .A2(KEYINPUT38), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n882), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n806), .B1(new_n720), .B2(new_n722), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n868), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n862), .A2(new_n860), .A3(new_n857), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT104), .B1(new_n866), .B2(new_n858), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n894), .B1(new_n899), .B2(new_n859), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n886), .A2(new_n891), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n881), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT40), .B1(new_n902), .B2(new_n892), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n896), .A2(KEYINPUT40), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n856), .B1(new_n904), .B2(new_n706), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT106), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n868), .A2(new_n903), .A3(new_n895), .ZN(new_n907));
  INV_X1    g0707(.A(new_n859), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n897), .B2(new_n898), .ZN(new_n909));
  AOI221_X4 g0709(.A(new_n881), .B1(new_n876), .B2(new_n890), .C1(new_n404), .C2(new_n885), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT38), .B1(new_n877), .B2(new_n879), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n909), .A2(new_n912), .A3(new_n894), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT40), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n907), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI211_X1 g0715(.A(new_n450), .B(new_n422), .C1(new_n721), .C2(new_n723), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n906), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT39), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n893), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n327), .A2(new_n668), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n902), .A2(KEYINPUT39), .A3(new_n892), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n902), .A2(new_n892), .ZN(new_n923));
  INV_X1    g0723(.A(new_n801), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n811), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n868), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n656), .A2(new_n869), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n922), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n696), .A2(new_n451), .A3(new_n704), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n659), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n928), .B(new_n930), .Z(new_n931));
  OAI22_X1  g0731(.A1(new_n917), .A2(new_n931), .B1(new_n211), .B2(new_n729), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n917), .A2(new_n931), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n855), .B1(new_n932), .B2(new_n933), .ZN(G367));
  AOI21_X1  g0734(.A(new_n259), .B1(new_n818), .B2(G97), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n757), .A2(KEYINPUT46), .A3(G116), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT46), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n756), .B2(new_n473), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n759), .A2(new_n453), .B1(new_n761), .B2(new_n820), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(G311), .B2(new_n817), .ZN(new_n941));
  OAI221_X1 g0741(.A(new_n941), .B1(new_n774), .B2(new_n828), .C1(new_n744), .C2(new_n770), .ZN(new_n942));
  AOI211_X1 g0742(.A(new_n939), .B(new_n942), .C1(G107), .C2(new_n752), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT109), .Z(new_n944));
  XOR2_X1   g0744(.A(KEYINPUT111), .B(G137), .Z(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n259), .B1(new_n223), .B2(new_n763), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT110), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n749), .A2(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n948), .B2(new_n947), .ZN(new_n950));
  INV_X1    g0750(.A(new_n761), .ZN(new_n951));
  AOI22_X1  g0751(.A1(G143), .A2(new_n817), .B1(new_n951), .B2(G159), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n952), .B1(new_n202), .B2(new_n756), .C1(new_n833), .C2(new_n759), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n745), .B2(G50), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n203), .B2(new_n830), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n944), .B1(new_n950), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT113), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n956), .B(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n736), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n792), .A2(new_n241), .ZN(new_n961));
  INV_X1    g0761(.A(new_n787), .ZN(new_n962));
  INV_X1    g0762(.A(new_n346), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n962), .B1(new_n683), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n735), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n615), .B1(new_n599), .B2(new_n669), .ZN(new_n966));
  OR3_X1    g0766(.A1(new_n633), .A2(new_n599), .A3(new_n669), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n960), .B(new_n965), .C1(new_n797), .C2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n629), .B1(new_n568), .B2(new_n669), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n622), .A2(new_n668), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n681), .A2(new_n972), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT45), .Z(new_n974));
  NOR2_X1   g0774(.A1(new_n681), .A2(new_n972), .ZN(new_n975));
  XNOR2_X1  g0775(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n975), .B(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n676), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n978), .B(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n679), .B1(new_n675), .B2(new_n678), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(KEYINPUT108), .B2(new_n672), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n672), .A2(KEYINPUT108), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n982), .B(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n727), .B1(new_n980), .B2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n684), .B(KEYINPUT41), .Z(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n731), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n972), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n989), .A2(new_n679), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT42), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n619), .B1(new_n970), .B2(new_n547), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n669), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n991), .A2(new_n993), .B1(KEYINPUT43), .B2(new_n968), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n994), .B(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n676), .A2(new_n989), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n996), .B(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n969), .B1(new_n988), .B2(new_n998), .ZN(G387));
  OAI21_X1  g0799(.A(new_n792), .B1(new_n238), .B2(new_n604), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n686), .B2(new_n789), .ZN(new_n1001));
  OR3_X1    g0801(.A1(new_n360), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1002));
  OAI21_X1  g0802(.A(KEYINPUT50), .B1(new_n360), .B2(G50), .ZN(new_n1003));
  AOI21_X1  g0803(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1002), .A2(new_n686), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n1001), .A2(new_n1005), .B1(new_n525), .B2(new_n683), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n732), .B1(new_n1006), .B2(new_n962), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n201), .A2(new_n759), .B1(new_n223), .B2(new_n756), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n335), .B(new_n1008), .C1(G97), .C2(new_n818), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n752), .A2(new_n963), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n749), .A2(G150), .ZN(new_n1011));
  INV_X1    g0811(.A(G159), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n360), .A2(new_n761), .B1(new_n1012), .B2(new_n765), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(G68), .B2(new_n740), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1014), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G322), .A2(new_n817), .B1(new_n951), .B2(G311), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n774), .B2(new_n759), .C1(new_n744), .C2(new_n453), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1018), .A2(KEYINPUT48), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(KEYINPUT48), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n752), .A2(G283), .B1(G294), .B2(new_n757), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT49), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n335), .B1(new_n473), .B2(new_n763), .C1(new_n828), .C2(new_n769), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1015), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1007), .B1(new_n1028), .B2(new_n736), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n675), .B2(new_n797), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n726), .A2(new_n984), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n684), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n726), .A2(new_n984), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1030), .B1(new_n730), .B2(new_n984), .C1(new_n1033), .C2(new_n1034), .ZN(G393));
  XNOR2_X1  g0835(.A(new_n978), .B(new_n676), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n1031), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n980), .A2(new_n1032), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n1038), .A3(new_n684), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1036), .A2(new_n731), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n972), .A2(new_n797), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT114), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n787), .B1(new_n552), .B2(new_n215), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n792), .B2(new_n245), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n778), .A2(G311), .B1(new_n817), .B2(G317), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT52), .Z(new_n1046));
  INV_X1    g0846(.A(G322), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1046), .B1(new_n1047), .B2(new_n828), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n741), .A2(new_n820), .B1(new_n453), .B2(new_n761), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G283), .B2(new_n757), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n259), .B1(new_n818), .B2(G107), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(new_n473), .C2(new_n830), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n749), .A2(G143), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n778), .A2(G159), .B1(new_n817), .B2(G150), .ZN(new_n1054));
  XOR2_X1   g0854(.A(KEYINPUT115), .B(KEYINPUT51), .Z(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1053), .B1(new_n1054), .B2(new_n1056), .C1(new_n744), .C2(new_n360), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n752), .A2(G77), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n335), .B1(new_n818), .B2(G87), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G50), .A2(new_n951), .B1(new_n757), .B2(G68), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n1048), .A2(new_n1052), .B1(new_n1057), .B2(new_n1062), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n735), .B(new_n1044), .C1(new_n1063), .C2(new_n736), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1042), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1039), .A2(new_n1040), .A3(new_n1065), .ZN(G390));
  OAI211_X1 g0866(.A(G330), .B(new_n806), .C1(new_n720), .C2(new_n722), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n868), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n925), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n909), .A2(new_n1071), .B1(new_n327), .B2(new_n668), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n919), .A2(new_n921), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n920), .B1(new_n882), .B2(new_n892), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n805), .A2(new_n351), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n703), .A2(new_n669), .A3(new_n1075), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1076), .A2(new_n924), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1074), .B1(new_n909), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT116), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g0880(.A(KEYINPUT116), .B(new_n1074), .C1(new_n909), .C2(new_n1077), .ZN(new_n1081));
  AOI221_X4 g0881(.A(new_n1070), .B1(new_n1072), .B2(new_n1073), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1069), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n909), .A2(new_n1067), .ZN(new_n1086));
  AND3_X1   g0886(.A1(new_n1069), .A2(new_n1077), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT117), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n868), .B2(new_n1068), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1071), .B1(new_n1089), .B2(new_n1086), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n909), .A2(new_n1088), .A3(new_n1067), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1087), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n929), .A2(new_n856), .A3(new_n659), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n1082), .A2(new_n1085), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1069), .A2(KEYINPUT117), .A3(new_n1086), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1095), .A2(new_n925), .A3(new_n1091), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1069), .A2(new_n1077), .A3(new_n1086), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1093), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1076), .A2(new_n924), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n868), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(KEYINPUT116), .B1(new_n1100), .B2(new_n1074), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1081), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1084), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n1070), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1083), .A2(new_n1084), .A3(new_n1069), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1098), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1094), .A2(new_n1106), .A3(new_n684), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n745), .A2(G97), .B1(G294), .B2(new_n749), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n759), .A2(new_n473), .B1(new_n765), .B2(new_n770), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n761), .A2(new_n525), .B1(new_n763), .B2(new_n203), .ZN(new_n1110));
  NOR4_X1   g0910(.A1(new_n758), .A2(new_n1109), .A3(new_n1110), .A4(new_n259), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1108), .A2(new_n1059), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n749), .A2(G125), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n259), .B1(new_n763), .B2(new_n201), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT118), .Z(new_n1115));
  XNOR2_X1  g0915(.A(KEYINPUT54), .B(G143), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1113), .B(new_n1115), .C1(new_n744), .C2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n756), .A2(new_n833), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT53), .ZN(new_n1119));
  INV_X1    g0919(.A(G128), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n759), .A2(new_n829), .B1(new_n765), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n951), .B2(new_n946), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1119), .B(new_n1122), .C1(new_n1012), .C2(new_n830), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n1117), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n737), .B1(new_n1112), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n815), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n732), .B1(new_n344), .B2(new_n1126), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1125), .B(new_n1127), .C1(new_n1073), .C2(new_n784), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1128), .B1(new_n1129), .B2(new_n731), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1107), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(G378));
  INV_X1    g0932(.A(new_n1093), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1106), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n928), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n439), .A2(new_n887), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n658), .A2(new_n440), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1137), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n450), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1136), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1138), .A2(new_n1140), .A3(new_n1136), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n904), .A2(new_n1144), .A3(new_n706), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1143), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1146), .A2(new_n1141), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n915), .B2(G330), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1135), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT122), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1144), .B1(new_n904), .B2(new_n706), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n915), .A2(G330), .A3(new_n1147), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(new_n1152), .A3(new_n928), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1149), .A2(new_n1150), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n928), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(KEYINPUT122), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1134), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT57), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1158), .B1(new_n1149), .B2(new_n1153), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n685), .B1(new_n1160), .B2(new_n1134), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1154), .A2(new_n731), .A3(new_n1156), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n732), .B1(G50), .B2(new_n1126), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT121), .Z(new_n1165));
  AOI22_X1  g0965(.A1(new_n778), .A2(G107), .B1(new_n817), .B2(G116), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n202), .B2(new_n763), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n741), .A2(new_n346), .B1(new_n223), .B2(new_n756), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n259), .A2(new_n278), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n552), .B2(new_n761), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1167), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1171), .B1(new_n203), .B2(new_n830), .C1(new_n770), .C2(new_n828), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT119), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT58), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1176));
  INV_X1    g0976(.A(G41), .ZN(new_n1177));
  AOI211_X1 g0977(.A(G50), .B(new_n1169), .C1(new_n471), .C2(new_n1177), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n759), .A2(new_n1120), .B1(new_n761), .B2(new_n829), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G125), .B2(new_n817), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1116), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n740), .A2(G137), .B1(new_n757), .B2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1180), .B(new_n1182), .C1(new_n833), .C2(new_n830), .ZN(new_n1183));
  XOR2_X1   g0983(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1184));
  XNOR2_X1  g0984(.A(new_n1183), .B(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n471), .B(new_n1177), .C1(new_n763), .C2(new_n1012), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n749), .B2(G124), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1178), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1175), .A2(new_n1176), .A3(new_n1188), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1165), .B1(new_n737), .B2(new_n1189), .C1(new_n1144), .C2(new_n785), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1163), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1162), .A2(new_n1192), .ZN(G375));
  INV_X1    g0993(.A(new_n1098), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1096), .A2(new_n1093), .A3(new_n1097), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(new_n987), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n909), .A2(new_n784), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT123), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n732), .B1(G68), .B2(new_n1126), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n741), .A2(new_n833), .B1(new_n761), .B2(new_n1116), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n765), .A2(new_n829), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n259), .B1(new_n763), .B2(new_n202), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n759), .A2(new_n945), .B1(new_n756), .B2(new_n1012), .ZN(new_n1203));
  NOR4_X1   g1003(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n201), .B2(new_n830), .C1(new_n1120), .C2(new_n828), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n745), .A2(G107), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n259), .B1(new_n778), .B2(G283), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n761), .A2(new_n473), .B1(new_n763), .B2(new_n206), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G294), .B2(new_n817), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1206), .A2(new_n1010), .A3(new_n1207), .A4(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n749), .A2(G303), .B1(G97), .B2(new_n757), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT124), .Z(new_n1212));
  OAI21_X1  g1012(.A(new_n1205), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1199), .B1(new_n1213), .B2(new_n736), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1198), .A2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1092), .B2(new_n730), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1196), .A2(new_n1217), .ZN(G381));
  AOI21_X1  g1018(.A(new_n1191), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n1131), .ZN(new_n1220));
  INV_X1    g1020(.A(G387), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n814), .A2(new_n842), .ZN(new_n1222));
  INV_X1    g1022(.A(G390), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(G393), .A2(G396), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  OR3_X1    g1025(.A1(new_n1220), .A2(G381), .A3(new_n1225), .ZN(G407));
  NOR2_X1   g1026(.A1(G375), .A2(G378), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n664), .A2(G343), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(G407), .A2(G213), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(KEYINPUT125), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT125), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(G407), .A2(new_n1232), .A3(G213), .A4(new_n1229), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(G409));
  XNOR2_X1  g1034(.A(G393), .B(new_n799), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  AND2_X1   g1036(.A1(G387), .A2(new_n1223), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(G387), .A2(new_n1223), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1236), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1221), .A2(G390), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(G387), .A2(new_n1223), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1240), .A2(new_n1235), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1239), .A2(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1096), .A2(KEYINPUT60), .A3(new_n1093), .A4(new_n1097), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n684), .ZN(new_n1245));
  OAI21_X1  g1045(.A(KEYINPUT60), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1245), .B1(new_n1195), .B2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1222), .B1(new_n1247), .B2(new_n1216), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT60), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1195), .B1(new_n1098), .B2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1250), .A2(new_n684), .A3(new_n1244), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1251), .A2(G384), .A3(new_n1217), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1248), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  AND3_X1   g1054(.A1(new_n1151), .A2(new_n928), .A3(new_n1152), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n731), .B1(new_n1255), .B2(new_n1155), .ZN(new_n1256));
  AND4_X1   g1056(.A1(new_n1107), .A2(new_n1256), .A3(new_n1130), .A4(new_n1190), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1134), .A2(new_n1154), .A3(new_n987), .A4(new_n1156), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1228), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1254), .B(new_n1259), .C1(new_n1219), .C2(new_n1131), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT127), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1260), .A2(new_n1261), .A3(KEYINPUT62), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT61), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1248), .A2(KEYINPUT126), .A3(new_n1252), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1228), .A2(G2897), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT126), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1253), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1253), .A2(new_n1268), .A3(new_n1266), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1131), .B1(new_n1162), .B2(new_n1192), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1228), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1270), .B(new_n1271), .C1(new_n1272), .C2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1262), .A2(new_n1263), .A3(new_n1276), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1261), .A2(KEYINPUT62), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1261), .A2(KEYINPUT62), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1260), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1243), .B1(new_n1277), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT63), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1243), .B1(new_n1282), .B2(new_n1260), .ZN(new_n1283));
  OR2_X1    g1083(.A1(new_n1260), .A2(new_n1282), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1283), .A2(new_n1263), .A3(new_n1276), .A4(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1281), .A2(new_n1285), .ZN(G405));
  OAI21_X1  g1086(.A(new_n1254), .B1(new_n1227), .B2(new_n1272), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1272), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(new_n1220), .A3(new_n1253), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1243), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1290), .B(new_n1291), .ZN(G402));
endmodule


