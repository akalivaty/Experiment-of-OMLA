//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 0 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT71), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G119), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT71), .A3(G116), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(G119), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT2), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G113), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n195), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(new_n199), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n202), .A2(new_n191), .A3(new_n193), .A4(new_n194), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT72), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n201), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n195), .A2(new_n200), .A3(KEYINPUT72), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G104), .ZN(new_n209));
  NOR3_X1   g023(.A1(new_n209), .A2(KEYINPUT3), .A3(G107), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G104), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT80), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(G104), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n214), .B1(new_n215), .B2(KEYINPUT3), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n214), .B(KEYINPUT3), .C1(new_n209), .C2(G107), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n213), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G101), .ZN(new_n220));
  INV_X1    g034(.A(G101), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n213), .B(new_n221), .C1(new_n216), .C2(new_n218), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(KEYINPUT4), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n219), .A2(new_n224), .A3(G101), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n208), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT87), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(G110), .B(G122), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT5), .A4(new_n194), .ZN(new_n230));
  NOR3_X1   g044(.A1(new_n190), .A2(KEYINPUT5), .A3(G119), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(new_n196), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT88), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n230), .A2(new_n232), .A3(KEYINPUT88), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n235), .A2(new_n203), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT82), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT81), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n209), .A2(G107), .ZN(new_n240));
  AOI211_X1 g054(.A(new_n239), .B(new_n221), .C1(new_n215), .C2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n221), .B1(new_n215), .B2(new_n240), .ZN(new_n243));
  OR2_X1    g057(.A1(new_n243), .A2(KEYINPUT81), .ZN(new_n244));
  AND4_X1   g058(.A1(new_n238), .A2(new_n222), .A3(new_n242), .A4(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n243), .A2(KEYINPUT81), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n246), .A2(new_n241), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n238), .B1(new_n247), .B2(new_n222), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n237), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n208), .A2(new_n223), .A3(KEYINPUT87), .A4(new_n225), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n228), .A2(new_n229), .A3(new_n249), .A4(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G224), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n253), .A2(KEYINPUT7), .ZN(new_n254));
  INV_X1    g068(.A(G146), .ZN(new_n255));
  AND2_X1   g069(.A1(KEYINPUT66), .A2(G143), .ZN(new_n256));
  NOR2_X1   g070(.A1(KEYINPUT66), .A2(G143), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n255), .A2(G143), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n255), .A2(G143), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT1), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n258), .A2(new_n260), .B1(new_n262), .B2(G128), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT66), .ZN(new_n264));
  INV_X1    g078(.A(G143), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(KEYINPUT66), .A2(G143), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(G146), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G128), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(KEYINPUT1), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n261), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n268), .A2(KEYINPUT70), .A3(new_n261), .A4(new_n270), .ZN(new_n274));
  AOI211_X1 g088(.A(G125), .B(new_n263), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT90), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n254), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n258), .A2(new_n260), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(KEYINPUT0), .A2(G128), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT65), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OR2_X1    g096(.A1(KEYINPUT0), .A2(G128), .ZN(new_n283));
  NAND3_X1  g097(.A1(KEYINPUT65), .A2(KEYINPUT0), .A3(G128), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n268), .A2(new_n261), .ZN(new_n286));
  OAI22_X1  g100(.A1(new_n279), .A2(new_n285), .B1(new_n286), .B2(new_n280), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G125), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n273), .A2(new_n274), .ZN(new_n289));
  INV_X1    g103(.A(new_n263), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n288), .B(KEYINPUT90), .C1(new_n291), .C2(G125), .ZN(new_n292));
  INV_X1    g106(.A(G125), .ZN(new_n293));
  OR2_X1    g107(.A1(new_n286), .A2(new_n280), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n278), .A2(new_n282), .A3(new_n284), .A4(new_n283), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n275), .A2(new_n296), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n277), .A2(new_n292), .B1(new_n297), .B2(new_n254), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n229), .B(KEYINPUT8), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n233), .A2(new_n203), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n222), .A2(new_n244), .A3(new_n242), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT82), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n247), .A2(new_n238), .A3(new_n222), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n301), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n237), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n299), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n251), .A2(new_n298), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G902), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT91), .ZN(new_n311));
  INV_X1    g125(.A(new_n229), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n226), .A2(new_n227), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n249), .A2(new_n250), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT6), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n316), .A2(KEYINPUT89), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(new_n251), .A3(new_n317), .ZN(new_n318));
  OAI221_X1 g132(.A(new_n312), .B1(KEYINPUT89), .B2(new_n316), .C1(new_n313), .C2(new_n314), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n297), .B(new_n253), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT91), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n308), .A2(new_n322), .A3(new_n309), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n311), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(G210), .B1(G237), .B2(G902), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n311), .A2(new_n321), .A3(new_n325), .A4(new_n323), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n188), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(G110), .B(G140), .ZN(new_n330));
  INV_X1    g144(.A(G227), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(G953), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n330), .B(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT69), .ZN(new_n334));
  INV_X1    g148(.A(G137), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(KEYINPUT11), .A3(G134), .ZN(new_n336));
  INV_X1    g150(.A(G134), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G137), .ZN(new_n338));
  AOI21_X1  g152(.A(KEYINPUT11), .B1(new_n335), .B2(G134), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n336), .B(new_n338), .C1(new_n339), .C2(KEYINPUT67), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT11), .ZN(new_n341));
  OAI211_X1 g155(.A(KEYINPUT67), .B(new_n341), .C1(new_n337), .C2(G137), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n334), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n336), .A2(new_n338), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT67), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n337), .A2(G137), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n346), .B1(new_n347), .B2(KEYINPUT11), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n345), .A2(new_n348), .A3(KEYINPUT69), .A4(new_n342), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n344), .A2(G131), .A3(new_n349), .ZN(new_n350));
  XOR2_X1   g164(.A(KEYINPUT68), .B(G131), .Z(new_n351));
  NAND4_X1  g165(.A1(new_n345), .A2(new_n348), .A3(new_n351), .A4(new_n342), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT84), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(G146), .B1(new_n266), .B2(new_n267), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT1), .ZN(new_n357));
  OAI21_X1  g171(.A(G128), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n273), .A2(new_n274), .B1(new_n358), .B2(new_n286), .ZN(new_n359));
  OR2_X1    g173(.A1(new_n359), .A2(new_n301), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n263), .B1(new_n273), .B2(new_n274), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n302), .A2(new_n361), .A3(new_n303), .ZN(new_n362));
  AOI211_X1 g176(.A(KEYINPUT12), .B(new_n355), .C1(new_n360), .C2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT12), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n360), .ZN(new_n365));
  INV_X1    g179(.A(new_n355), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n350), .A2(KEYINPUT83), .A3(new_n352), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT83), .B1(new_n350), .B2(new_n352), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(KEYINPUT10), .B(new_n291), .C1(new_n245), .C2(new_n248), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n373), .B1(new_n359), .B2(new_n301), .ZN(new_n374));
  INV_X1    g188(.A(new_n287), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(new_n223), .A3(new_n225), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n371), .A2(new_n372), .A3(new_n374), .A4(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT85), .B1(new_n368), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n359), .A2(new_n301), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n245), .A2(new_n248), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n379), .B1(new_n380), .B2(new_n361), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT12), .B1(new_n381), .B2(new_n355), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n365), .A2(new_n364), .A3(new_n366), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n382), .A2(KEYINPUT85), .A3(new_n377), .A4(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n333), .B1(new_n378), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n333), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n377), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT86), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n372), .A2(new_n374), .A3(new_n376), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n353), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT86), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n388), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n390), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n386), .A2(G469), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G469), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n397), .A2(new_n309), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n387), .B1(new_n392), .B2(new_n377), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n382), .A2(new_n377), .A3(new_n387), .A4(new_n383), .ZN(new_n401));
  AOI21_X1  g215(.A(G902), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n398), .B1(new_n402), .B2(new_n397), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n396), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT9), .B(G234), .ZN(new_n405));
  OAI21_X1  g219(.A(G221), .B1(new_n405), .B2(G902), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n329), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G217), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n408), .B1(G234), .B2(new_n309), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n252), .A2(G221), .A3(G234), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT79), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT22), .B(G137), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n411), .B(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT74), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n192), .B2(G128), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT23), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n269), .A2(G119), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT23), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n192), .A2(G128), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n417), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n418), .A2(new_n421), .ZN(new_n423));
  XOR2_X1   g237(.A(KEYINPUT24), .B(G110), .Z(new_n424));
  OAI22_X1  g238(.A1(new_n422), .A2(G110), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT76), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT16), .ZN(new_n427));
  INV_X1    g241(.A(G140), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n426), .A2(new_n427), .A3(new_n428), .A4(G125), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n293), .A2(KEYINPUT16), .A3(G140), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n429), .B1(new_n430), .B2(new_n426), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n428), .A2(G125), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n293), .A2(G140), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n433), .A3(KEYINPUT16), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n431), .A2(G146), .A3(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(G125), .B(G140), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n255), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n425), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT77), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n434), .A2(G146), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n427), .A2(new_n428), .A3(G125), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n293), .A2(G140), .ZN(new_n442));
  NOR2_X1   g256(.A1(KEYINPUT76), .A2(KEYINPUT16), .ZN(new_n443));
  AOI22_X1  g257(.A1(KEYINPUT76), .A2(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n439), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n431), .A2(KEYINPUT77), .A3(G146), .A4(new_n434), .ZN(new_n446));
  AOI21_X1  g260(.A(G146), .B1(new_n431), .B2(new_n434), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n445), .A2(new_n446), .B1(new_n447), .B2(KEYINPUT78), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT78), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n441), .A2(KEYINPUT76), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n450), .A2(new_n429), .B1(new_n436), .B2(KEYINPUT16), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n449), .B1(new_n451), .B2(G146), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n417), .A2(new_n420), .A3(KEYINPUT75), .A4(new_n421), .ZN(new_n454));
  INV_X1    g268(.A(G110), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT75), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n455), .B1(new_n422), .B2(new_n456), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n454), .A2(new_n457), .B1(new_n423), .B2(new_n424), .ZN(new_n458));
  AOI211_X1 g272(.A(new_n414), .B(new_n438), .C1(new_n453), .C2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n453), .A2(new_n458), .ZN(new_n460));
  INV_X1    g274(.A(new_n438), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n413), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(KEYINPUT25), .B1(new_n463), .B2(new_n309), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT25), .ZN(new_n465));
  NOR4_X1   g279(.A1(new_n459), .A2(new_n462), .A3(new_n465), .A4(G902), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n409), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n463), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n409), .A2(G902), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n467), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n353), .A2(new_n375), .ZN(new_n472));
  INV_X1    g286(.A(new_n338), .ZN(new_n473));
  OAI21_X1  g287(.A(G131), .B1(new_n473), .B2(new_n347), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n352), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n291), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n472), .A2(KEYINPUT30), .A3(new_n477), .ZN(new_n478));
  XOR2_X1   g292(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n287), .B1(new_n350), .B2(new_n352), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n361), .A2(new_n475), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n478), .A2(new_n483), .A3(new_n208), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n472), .A2(new_n207), .A3(new_n477), .ZN(new_n485));
  INV_X1    g299(.A(G237), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n252), .A3(G210), .ZN(new_n487));
  XOR2_X1   g301(.A(new_n487), .B(KEYINPUT27), .Z(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT26), .B(G101), .ZN(new_n489));
  XOR2_X1   g303(.A(new_n488), .B(new_n489), .Z(new_n490));
  NAND3_X1  g304(.A1(new_n484), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT31), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n484), .A2(KEYINPUT31), .A3(new_n485), .A4(new_n490), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n208), .B1(new_n481), .B2(new_n482), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n485), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT28), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT28), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n485), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n490), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n495), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT32), .ZN(new_n505));
  NOR2_X1   g319(.A1(G472), .A2(G902), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n493), .A2(new_n494), .B1(new_n501), .B2(new_n502), .ZN(new_n508));
  INV_X1    g322(.A(new_n506), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT32), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n484), .A2(new_n485), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n502), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n498), .A2(new_n500), .A3(new_n490), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT29), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT73), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n517), .B1(new_n485), .B2(new_n496), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n472), .A2(new_n477), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT73), .B1(new_n519), .B2(new_n208), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT28), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n500), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n490), .A2(KEYINPUT29), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n516), .B(new_n309), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G472), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n471), .B1(new_n511), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n445), .A2(new_n446), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n447), .A2(KEYINPUT78), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT92), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n486), .A2(new_n252), .A3(G143), .A4(G214), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n266), .A2(new_n267), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n486), .A2(new_n252), .A3(G214), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n529), .B(new_n530), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n530), .A2(new_n529), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n351), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n533), .A2(new_n535), .A3(KEYINPUT17), .A4(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n527), .A2(new_n452), .A3(new_n528), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT96), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n530), .A2(new_n529), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n256), .A2(new_n257), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n486), .A2(new_n252), .A3(G214), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n534), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT93), .B1(new_n544), .B2(new_n536), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n533), .A2(new_n535), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT93), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n547), .A3(new_n351), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT17), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n544), .A2(new_n536), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n545), .A2(new_n548), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT96), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n448), .A2(new_n552), .A3(new_n452), .A4(new_n537), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n539), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n544), .A2(KEYINPUT18), .A3(G131), .ZN(new_n555));
  NAND2_X1  g369(.A1(KEYINPUT18), .A2(G131), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n546), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n436), .B(new_n255), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(G113), .B(G122), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT95), .B(G104), .ZN(new_n561));
  XOR2_X1   g375(.A(new_n560), .B(new_n561), .Z(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n554), .A2(new_n559), .A3(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT19), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n436), .B1(KEYINPUT94), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n566), .B1(new_n436), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n435), .B1(new_n568), .B2(G146), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n548), .A2(new_n550), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n569), .B1(new_n570), .B2(new_n545), .ZN(new_n571));
  INV_X1    g385(.A(new_n559), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n562), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n564), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT20), .ZN(new_n575));
  NOR2_X1   g389(.A1(G475), .A2(G902), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT97), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n574), .A2(KEYINPUT97), .A3(new_n575), .A4(new_n576), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n574), .A2(new_n576), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT20), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT98), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n554), .A2(new_n559), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n562), .ZN(new_n586));
  AOI21_X1  g400(.A(G902), .B1(new_n586), .B2(new_n564), .ZN(new_n587));
  INV_X1    g401(.A(G475), .ZN(new_n588));
  OR2_X1    g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n583), .A2(new_n584), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n584), .B1(new_n583), .B2(new_n589), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n265), .A2(G128), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n592), .B1(new_n541), .B2(G128), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n337), .ZN(new_n594));
  XNOR2_X1  g408(.A(G116), .B(G122), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(new_n211), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n593), .A2(KEYINPUT13), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n541), .A2(G128), .ZN(new_n598));
  OAI21_X1  g412(.A(G134), .B1(new_n598), .B2(KEYINPUT13), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n594), .B(new_n596), .C1(new_n597), .C2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n593), .B(new_n337), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n595), .A2(new_n211), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT14), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n595), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n190), .A2(KEYINPUT14), .A3(G122), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(G107), .A3(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT99), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n600), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n405), .A2(new_n408), .A3(G953), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n600), .B(new_n610), .C1(new_n603), .C2(new_n608), .ZN(new_n613));
  AOI21_X1  g427(.A(G902), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(G478), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(KEYINPUT15), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n614), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(G234), .A2(G237), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n618), .A2(G902), .A3(G953), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT21), .B(G898), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n618), .A2(G952), .A3(new_n252), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n617), .A2(new_n624), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n590), .A2(new_n591), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n407), .A2(new_n526), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT100), .B(G101), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G3));
  NAND2_X1  g443(.A1(new_n327), .A2(new_n328), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(new_n624), .A3(new_n187), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n576), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n564), .B2(new_n573), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n580), .B1(new_n575), .B2(new_n634), .ZN(new_n635));
  AOI211_X1 g449(.A(KEYINPUT20), .B(new_n633), .C1(new_n564), .C2(new_n573), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(KEYINPUT97), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n589), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT98), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n583), .A2(new_n584), .A3(new_n589), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n612), .A2(new_n613), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT33), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n612), .A2(new_n644), .A3(new_n613), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n643), .A2(G478), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n615), .A2(new_n309), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n614), .B2(new_n615), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n646), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n647), .B1(new_n646), .B2(new_n649), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT102), .B1(new_n641), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n655));
  AOI211_X1 g469(.A(new_n655), .B(new_n652), .C1(new_n639), .C2(new_n640), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n509), .B1(new_n495), .B2(new_n503), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n504), .A2(new_n309), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n658), .B1(new_n659), .B2(G472), .ZN(new_n660));
  INV_X1    g474(.A(new_n406), .ZN(new_n661));
  AOI211_X1 g475(.A(new_n661), .B(new_n471), .C1(new_n396), .C2(new_n403), .ZN(new_n662));
  AND4_X1   g476(.A1(new_n632), .A2(new_n657), .A3(new_n660), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT34), .B(G104), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  INV_X1    g479(.A(new_n471), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n404), .A2(new_n660), .A3(new_n666), .A4(new_n406), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n634), .A2(new_n575), .ZN(new_n668));
  OAI22_X1  g482(.A1(new_n668), .A2(new_n636), .B1(new_n587), .B2(new_n588), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n617), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n329), .A2(new_n624), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT35), .B(G107), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G9));
  NAND2_X1  g488(.A1(new_n460), .A2(new_n461), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT103), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n414), .A2(KEYINPUT36), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n469), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n467), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n660), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n407), .A2(new_n626), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT37), .B(G110), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  OR2_X1    g499(.A1(new_n464), .A2(new_n466), .ZN(new_n686));
  AOI22_X1  g500(.A1(new_n686), .A2(new_n409), .B1(new_n678), .B2(new_n469), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n511), .B2(new_n525), .ZN(new_n688));
  INV_X1    g502(.A(G900), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n622), .B1(new_n619), .B2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n670), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n661), .B1(new_n396), .B2(new_n403), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n688), .A2(new_n693), .A3(new_n329), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  XOR2_X1   g510(.A(new_n690), .B(KEYINPUT39), .Z(new_n697));
  NAND2_X1  g511(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT40), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT106), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT40), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n698), .B(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OR2_X1    g518(.A1(new_n518), .A2(new_n520), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n309), .B1(new_n705), .B2(new_n490), .ZN(new_n706));
  INV_X1    g520(.A(new_n512), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n502), .ZN(new_n708));
  OAI21_X1  g522(.A(G472), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n511), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n511), .A2(KEYINPUT105), .A3(new_n709), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n630), .B(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n590), .A2(new_n591), .ZN(new_n717));
  INV_X1    g531(.A(new_n617), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n687), .A2(new_n718), .A3(new_n187), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n716), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n700), .A2(new_n704), .A3(new_n714), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n531), .ZN(G45));
  AOI21_X1  g536(.A(new_n505), .B1(new_n504), .B2(new_n506), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n508), .A2(KEYINPUT32), .A3(new_n509), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n525), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AND4_X1   g539(.A1(new_n725), .A2(new_n694), .A3(new_n329), .A4(new_n680), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n653), .B(new_n691), .C1(new_n590), .C2(new_n591), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G146), .ZN(G48));
  AOI22_X1  g544(.A1(new_n507), .A2(new_n510), .B1(new_n524), .B2(G472), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n399), .B1(new_n368), .B2(new_n389), .ZN(new_n732));
  OAI21_X1  g546(.A(G469), .B1(new_n732), .B2(G902), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n402), .A2(new_n397), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n734), .A3(new_n406), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n731), .A2(new_n471), .A3(new_n735), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n632), .B(new_n736), .C1(new_n654), .C2(new_n656), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT41), .B(G113), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G15));
  AND3_X1   g553(.A1(new_n329), .A2(new_n624), .A3(new_n670), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G116), .ZN(G18));
  AND3_X1   g556(.A1(new_n733), .A2(new_n734), .A3(new_n406), .ZN(new_n743));
  AND4_X1   g557(.A1(new_n725), .A2(new_n329), .A3(new_n680), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n626), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G119), .ZN(G21));
  NAND3_X1  g560(.A1(new_n641), .A2(new_n718), .A3(new_n329), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT108), .ZN(new_n748));
  AOI22_X1  g562(.A1(new_n522), .A2(new_n502), .B1(new_n493), .B2(new_n494), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n506), .B(KEYINPUT107), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n748), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n495), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n490), .B1(new_n521), .B2(new_n500), .ZN(new_n754));
  OAI211_X1 g568(.A(KEYINPUT108), .B(new_n750), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n752), .A2(new_n755), .B1(G472), .B2(new_n659), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n756), .A2(new_n666), .A3(new_n624), .A4(new_n743), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n747), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G122), .ZN(G24));
  NAND2_X1  g573(.A1(new_n329), .A2(new_n743), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n752), .A2(new_n755), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n659), .A2(G472), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n763), .A3(new_n680), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n728), .A2(new_n761), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G125), .ZN(G27));
  NAND3_X1  g581(.A1(new_n382), .A2(new_n377), .A3(new_n383), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT85), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n384), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT109), .B1(new_n771), .B2(new_n333), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT109), .ZN(new_n773));
  AOI211_X1 g587(.A(new_n773), .B(new_n387), .C1(new_n770), .C2(new_n384), .ZN(new_n774));
  OAI211_X1 g588(.A(G469), .B(new_n395), .C1(new_n772), .C2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n403), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n776), .A2(new_n526), .A3(new_n406), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n327), .A2(new_n187), .A3(new_n328), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n727), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(new_n779), .A3(KEYINPUT42), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT42), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n661), .B1(new_n775), .B2(new_n403), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n526), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n327), .A2(new_n187), .A3(new_n328), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n641), .A2(new_n653), .A3(new_n691), .A4(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n781), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n780), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G131), .ZN(G33));
  NOR2_X1   g602(.A1(new_n692), .A2(new_n778), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n782), .A2(new_n526), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(KEYINPUT110), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT110), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n782), .A2(new_n792), .A3(new_n789), .A4(new_n526), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G134), .ZN(G36));
  AOI21_X1  g609(.A(KEYINPUT45), .B1(new_n386), .B2(new_n395), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n397), .ZN(new_n797));
  OAI211_X1 g611(.A(KEYINPUT45), .B(new_n395), .C1(new_n772), .C2(new_n774), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n398), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n799), .A2(KEYINPUT46), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n734), .B1(new_n799), .B2(KEYINPUT46), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(new_n406), .A3(new_n697), .A4(new_n784), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT43), .B1(new_n717), .B2(KEYINPUT111), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n717), .A2(new_n653), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n660), .A2(new_n687), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT44), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n803), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT44), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n806), .A2(new_n807), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G137), .ZN(G39));
  OAI21_X1  g627(.A(new_n406), .B1(new_n800), .B2(new_n801), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT47), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n779), .A2(new_n731), .A3(new_n471), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT112), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G140), .ZN(G42));
  INV_X1    g634(.A(new_n714), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n653), .A2(new_n666), .A3(new_n187), .A4(new_n406), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n733), .A2(new_n734), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n823), .A2(KEYINPUT49), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(KEYINPUT49), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n821), .A2(new_n826), .A3(new_n717), .A4(new_n716), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT42), .B1(new_n777), .B2(new_n779), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n783), .A2(new_n785), .A3(new_n781), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n744), .A2(new_n626), .B1(new_n736), .B2(new_n740), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n737), .A2(new_n832), .A3(new_n758), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n694), .A2(new_n329), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n639), .A2(new_n640), .A3(new_n624), .A4(new_n617), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n835), .A2(new_n836), .A3(new_n681), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n639), .A2(new_n640), .A3(new_n718), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n667), .A2(new_n838), .A3(new_n631), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n837), .A2(new_n839), .A3(KEYINPUT114), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n653), .B1(new_n590), .B2(new_n591), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT113), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n667), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n641), .A2(KEYINPUT113), .A3(new_n653), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n843), .A2(new_n844), .A3(new_n845), .A4(new_n632), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n627), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n590), .A2(new_n591), .A3(new_n617), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n632), .A2(new_n849), .A3(new_n662), .A4(new_n660), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n848), .B1(new_n850), .B2(new_n683), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n840), .A2(new_n847), .A3(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n669), .A2(new_n718), .A3(new_n690), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n688), .A2(new_n694), .A3(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n776), .A2(new_n406), .A3(new_n680), .A4(new_n756), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n854), .B1(new_n855), .B2(new_n727), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n784), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n794), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n834), .A2(new_n852), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n630), .A2(new_n718), .A3(new_n187), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n717), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n680), .A2(new_n690), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n714), .A2(new_n862), .A3(new_n782), .A4(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(new_n695), .A3(new_n729), .A4(new_n766), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT52), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n828), .B1(new_n860), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT115), .B1(new_n831), .B2(new_n833), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n688), .A2(new_n329), .A3(new_n743), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n526), .A2(new_n743), .ZN(new_n871));
  OAI22_X1  g685(.A1(new_n870), .A2(new_n836), .B1(new_n871), .B2(new_n671), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n747), .A2(new_n757), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT115), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n787), .A2(new_n874), .A3(new_n875), .A4(new_n737), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT114), .B1(new_n837), .B2(new_n839), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n850), .A2(new_n683), .A3(new_n848), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n878), .A2(new_n627), .A3(new_n879), .A4(new_n846), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n756), .A2(new_n329), .A3(new_n680), .A4(new_n743), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n695), .B1(new_n727), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT52), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT53), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n880), .A2(new_n858), .A3(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT52), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n865), .B(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n877), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n867), .A2(new_n868), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n787), .A2(new_n874), .A3(new_n737), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n890), .A2(new_n880), .A3(new_n858), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n883), .A2(new_n828), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(new_n887), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n868), .B1(new_n867), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n806), .A2(new_n622), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n756), .A2(new_n666), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n823), .A2(new_n406), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n784), .B(new_n898), .C1(new_n816), .C2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n897), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n716), .A2(new_n188), .A3(new_n743), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n806), .A2(new_n622), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT116), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT50), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n903), .A2(new_n904), .A3(KEYINPUT50), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n778), .A2(new_n735), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n910), .A2(new_n471), .A3(new_n623), .ZN(new_n911));
  AND4_X1   g725(.A1(new_n717), .A2(new_n911), .A3(new_n652), .A4(new_n821), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n896), .A2(new_n910), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n912), .B1(new_n913), .B2(new_n765), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n900), .A2(new_n907), .A3(new_n908), .A4(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT51), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n657), .A2(new_n821), .A3(new_n911), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(G952), .A3(new_n252), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n898), .B2(new_n761), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT48), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n913), .B2(new_n526), .ZN(new_n922));
  INV_X1    g736(.A(new_n526), .ZN(new_n923));
  NOR4_X1   g737(.A1(new_n896), .A2(KEYINPUT48), .A3(new_n923), .A4(new_n910), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n920), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n915), .B2(new_n916), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n895), .A2(new_n917), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(G952), .A2(G953), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n827), .B1(new_n927), .B2(new_n928), .ZN(G75));
  NOR2_X1   g743(.A1(new_n252), .A2(G952), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT117), .Z(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n309), .B1(new_n867), .B2(new_n888), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT56), .B1(new_n933), .B2(G210), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n318), .A2(new_n319), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n320), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT55), .Z(new_n937));
  OR2_X1    g751(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n934), .A2(new_n937), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n932), .B1(new_n938), .B2(new_n939), .ZN(G51));
  XNOR2_X1  g754(.A(new_n398), .B(KEYINPUT57), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n868), .B1(new_n867), .B2(new_n888), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n941), .B1(new_n889), .B2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n732), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n933), .A2(new_n798), .A3(new_n797), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n930), .B1(new_n945), .B2(new_n946), .ZN(G54));
  NAND3_X1  g761(.A1(new_n933), .A2(KEYINPUT58), .A3(G475), .ZN(new_n948));
  INV_X1    g762(.A(new_n574), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n950), .A2(new_n951), .A3(new_n930), .ZN(G60));
  INV_X1    g766(.A(KEYINPUT119), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n643), .A2(new_n645), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  XOR2_X1   g769(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(new_n648), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n877), .A2(new_n885), .A3(new_n887), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT53), .B1(new_n891), .B2(new_n887), .ZN(new_n961));
  OAI21_X1  g775(.A(KEYINPUT54), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n867), .A2(new_n868), .A3(new_n888), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n953), .B1(new_n964), .B2(new_n932), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n958), .B1(new_n889), .B2(new_n942), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n966), .A2(KEYINPUT119), .A3(new_n931), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n955), .B1(new_n895), .B2(new_n957), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n965), .A2(new_n967), .A3(new_n968), .ZN(G63));
  INV_X1    g783(.A(KEYINPUT121), .ZN(new_n970));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT60), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n867), .B2(new_n888), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n970), .B1(new_n973), .B2(new_n463), .ZN(new_n974));
  INV_X1    g788(.A(new_n972), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(new_n960), .B2(new_n961), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n976), .A2(KEYINPUT121), .A3(new_n468), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n678), .B(new_n975), .C1(new_n960), .C2(new_n961), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n931), .A2(KEYINPUT61), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n974), .A2(new_n977), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n932), .B1(new_n976), .B2(new_n468), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT120), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n973), .A2(new_n982), .A3(new_n678), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n978), .A2(KEYINPUT120), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n981), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n980), .B1(new_n985), .B2(KEYINPUT61), .ZN(G66));
  INV_X1    g800(.A(G224), .ZN(new_n987));
  OAI21_X1  g801(.A(G953), .B1(new_n620), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n880), .A2(new_n833), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n988), .B1(new_n989), .B2(G953), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n935), .B1(G898), .B2(new_n252), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT122), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n990), .B(new_n992), .ZN(G69));
  NAND2_X1  g807(.A1(new_n478), .A2(new_n483), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT123), .Z(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(new_n568), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n849), .B1(new_n843), .B2(new_n845), .ZN(new_n997));
  OR4_X1    g811(.A1(new_n923), .A2(new_n997), .A3(new_n698), .A4(new_n778), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n812), .A2(new_n819), .A3(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT62), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n882), .B1(new_n726), .B2(new_n728), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n721), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT124), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1000), .B1(new_n721), .B2(new_n1001), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT125), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n999), .A2(new_n252), .A3(new_n1003), .A4(new_n1006), .ZN(new_n1007));
  NAND3_X1  g821(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n996), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n331), .A2(G900), .A3(G953), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n802), .A2(new_n406), .A3(new_n697), .ZN(new_n1011));
  NOR3_X1   g825(.A1(new_n1011), .A2(new_n923), .A3(new_n747), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1001), .A2(new_n787), .A3(new_n794), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1014), .A2(new_n812), .A3(new_n819), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(KEYINPUT126), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT126), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n1014), .A2(new_n812), .A3(new_n819), .A4(new_n1017), .ZN(new_n1018));
  AND2_X1   g832(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1010), .B1(new_n1019), .B2(G953), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1009), .B1(new_n1020), .B2(new_n996), .ZN(G72));
  NAND2_X1  g835(.A1(new_n707), .A2(new_n502), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1016), .A2(new_n989), .A3(new_n1018), .ZN(new_n1023));
  XNOR2_X1  g837(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1024));
  NAND2_X1  g838(.A1(G472), .A2(G902), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1024), .B(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1022), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(new_n708), .ZN(new_n1028));
  NAND4_X1  g842(.A1(new_n999), .A2(new_n989), .A3(new_n1003), .A4(new_n1006), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1028), .B1(new_n1029), .B2(new_n1026), .ZN(new_n1030));
  AND2_X1   g844(.A1(new_n867), .A2(new_n893), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n513), .A2(new_n491), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1032), .A2(new_n1026), .ZN(new_n1033));
  OAI22_X1  g847(.A1(new_n1031), .A2(new_n1033), .B1(G952), .B2(new_n252), .ZN(new_n1034));
  NOR3_X1   g848(.A1(new_n1027), .A2(new_n1030), .A3(new_n1034), .ZN(G57));
endmodule


