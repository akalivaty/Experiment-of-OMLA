//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1264, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(new_n204), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G107), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n206), .B1(new_n219), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n209), .B1(new_n212), .B2(new_n213), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT64), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  INV_X1    g0040(.A(G50), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n215), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n240), .B(new_n246), .Z(G351));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n210), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n204), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G150), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  OAI22_X1  g0054(.A1(new_n250), .A2(new_n251), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G58), .A2(G68), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n204), .B1(new_n256), .B2(new_n241), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n249), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n249), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n203), .A2(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(new_n241), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n261), .A2(new_n264), .B1(new_n241), .B2(new_n260), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT9), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n266), .B1(KEYINPUT69), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(KEYINPUT69), .B2(new_n267), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT69), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n266), .A2(new_n270), .A3(KEYINPUT9), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(G1), .A3(G13), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G274), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n273), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(new_n277), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n279), .B1(G226), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT3), .B(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G222), .A2(G1698), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(G223), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n283), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n287), .B(new_n280), .C1(G77), .C2(new_n283), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n282), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT65), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n282), .A2(KEYINPUT65), .A3(new_n288), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n269), .A2(new_n271), .B1(G190), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT68), .B(G200), .ZN(new_n295));
  OAI21_X1  g0095(.A(KEYINPUT70), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT70), .ZN(new_n297));
  INV_X1    g0097(.A(new_n295), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n291), .A2(new_n297), .A3(new_n298), .A4(new_n292), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n294), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT10), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT10), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n294), .A2(new_n302), .A3(new_n296), .A4(new_n299), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G179), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n293), .A2(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n306), .B(new_n266), .C1(G169), .C2(new_n293), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n283), .A2(G232), .A3(new_n285), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT66), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n309), .B(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G33), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT3), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT3), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G33), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NOR3_X1   g0116(.A1(new_n316), .A2(new_n216), .A3(new_n285), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(G107), .B2(new_n316), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n273), .B1(new_n311), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G274), .ZN(new_n320));
  INV_X1    g0120(.A(new_n210), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n272), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n277), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n278), .A2(new_n273), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(new_n222), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n319), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n305), .ZN(new_n327));
  INV_X1    g0127(.A(new_n250), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n328), .A2(new_n253), .B1(G20), .B2(G77), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT15), .B(G87), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n329), .B1(new_n251), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT67), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n259), .B(new_n332), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n331), .A2(new_n249), .B1(new_n221), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G13), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n335), .A2(G1), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(new_n332), .A3(G20), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n259), .A2(KEYINPUT67), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n249), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n339), .A2(G77), .A3(new_n262), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G169), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n319), .B2(new_n325), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n327), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n341), .B1(new_n326), .B2(G190), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n298), .B1(new_n319), .B2(new_n325), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G232), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G1698), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n283), .B(new_n350), .C1(G226), .C2(G1698), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G33), .A2(G97), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n280), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n279), .B1(G238), .B2(new_n281), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT13), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n273), .B1(new_n351), .B2(new_n352), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n323), .B1(new_n324), .B2(new_n216), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT13), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G190), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n339), .A2(G68), .A3(new_n262), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT71), .ZN(new_n365));
  XOR2_X1   g0165(.A(KEYINPUT72), .B(KEYINPUT12), .Z(new_n366));
  NAND2_X1  g0166(.A1(new_n337), .A2(new_n338), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n366), .B1(new_n367), .B2(G68), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n215), .A2(G20), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT12), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n336), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n368), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  OAI221_X1 g0172(.A(new_n369), .B1(new_n251), .B2(new_n221), .C1(new_n254), .C2(new_n241), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n249), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n374), .B(KEYINPUT11), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n365), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G200), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(new_n357), .B2(new_n360), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n363), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n361), .A2(G169), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT14), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n357), .A2(G179), .A3(new_n360), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT14), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n361), .A2(new_n383), .A3(G169), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n379), .B1(new_n385), .B2(new_n376), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT73), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n345), .B(new_n348), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n386), .A2(new_n387), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n308), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n323), .B1(new_n324), .B2(new_n349), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n362), .A2(KEYINPUT77), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n362), .A2(KEYINPUT77), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n314), .A2(G33), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT74), .B1(new_n312), .B2(KEYINPUT3), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT74), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n398), .A2(new_n314), .A3(G33), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n396), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  MUX2_X1   g0200(.A(G223), .B(G226), .S(G1698), .Z(new_n401));
  AOI22_X1  g0201(.A1(new_n400), .A2(new_n401), .B1(G33), .B2(G87), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n392), .B(new_n395), .C1(new_n402), .C2(new_n273), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n402), .A2(new_n273), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n404), .A2(new_n391), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n403), .B1(new_n405), .B2(G200), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n250), .A2(new_n263), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n407), .A2(new_n261), .B1(new_n260), .B2(new_n250), .ZN(new_n408));
  INV_X1    g0208(.A(G58), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n409), .A2(new_n215), .ZN(new_n410));
  OAI21_X1  g0210(.A(G20), .B1(new_n410), .B2(new_n256), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n253), .A2(G159), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT16), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n398), .B1(new_n314), .B2(G33), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n312), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n313), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT7), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n420), .A3(new_n204), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT7), .B1(new_n400), .B2(G20), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n422), .A3(G68), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT75), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n397), .A2(new_n399), .ZN(new_n425));
  AOI21_X1  g0225(.A(G20), .B1(new_n425), .B2(new_n313), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n215), .B1(new_n426), .B2(new_n420), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT75), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(new_n428), .A3(new_n422), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n416), .B1(new_n424), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n420), .A2(new_n204), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n283), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT76), .B1(new_n314), .B2(G33), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT76), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n434), .A2(new_n312), .A3(KEYINPUT3), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n435), .A3(new_n315), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n204), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n432), .B1(new_n437), .B2(KEYINPUT7), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n413), .B1(new_n438), .B2(G68), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n249), .B1(new_n439), .B2(KEYINPUT16), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n406), .B(new_n408), .C1(new_n430), .C2(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(KEYINPUT78), .A2(KEYINPUT17), .ZN(new_n442));
  NAND2_X1  g0242(.A1(KEYINPUT78), .A2(KEYINPUT17), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n441), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n408), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n428), .B1(new_n427), .B2(new_n422), .ZN(new_n447));
  AND4_X1   g0247(.A1(new_n428), .A2(new_n421), .A3(new_n422), .A4(G68), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n415), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n249), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n437), .A2(KEYINPUT7), .ZN(new_n451));
  INV_X1    g0251(.A(new_n432), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n451), .A2(G68), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n413), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n450), .B1(new_n455), .B2(new_n414), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n446), .B1(new_n449), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(new_n406), .A3(new_n443), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n445), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n408), .B1(new_n430), .B2(new_n440), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n405), .A2(G179), .ZN(new_n461));
  OAI21_X1  g0261(.A(G169), .B1(new_n404), .B2(new_n391), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT18), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT18), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n460), .A2(new_n466), .A3(new_n463), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n459), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n390), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n259), .A2(G97), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n203), .A2(G33), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n450), .A2(new_n259), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n472), .B1(new_n475), .B2(G97), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n438), .A2(G107), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT6), .ZN(new_n479));
  INV_X1    g0279(.A(G97), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n479), .A2(new_n480), .A3(G107), .ZN(new_n481));
  XNOR2_X1  g0281(.A(G97), .B(G107), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(new_n479), .ZN(new_n483));
  OAI22_X1  g0283(.A1(new_n483), .A2(new_n204), .B1(new_n221), .B2(new_n254), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n478), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n477), .B1(new_n486), .B2(new_n249), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n313), .A2(new_n315), .A3(G250), .A4(G1698), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G33), .A2(G283), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n222), .A2(G1698), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n425), .A2(new_n313), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT4), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g0294(.A1(KEYINPUT4), .A2(G244), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n313), .A2(new_n315), .A3(new_n495), .A4(new_n285), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT79), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n283), .A2(KEYINPUT79), .A3(new_n285), .A4(new_n495), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n273), .B1(new_n494), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n276), .A2(G1), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G41), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT80), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(new_n503), .B2(G41), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n503), .A2(G41), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT80), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n505), .A2(new_n322), .A3(new_n507), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n502), .A2(new_n504), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n273), .B(G257), .C1(new_n511), .C2(new_n508), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n501), .A2(G190), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n492), .A2(new_n493), .ZN(new_n515));
  INV_X1    g0315(.A(new_n490), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n500), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n280), .ZN(new_n518));
  INV_X1    g0318(.A(new_n513), .ZN(new_n519));
  AOI21_X1  g0319(.A(G200), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n487), .B1(new_n514), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT22), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(new_n217), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n425), .A2(new_n204), .A3(new_n313), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n204), .A2(G87), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n522), .B1(new_n316), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n204), .A2(G33), .A3(G116), .ZN(new_n527));
  OAI21_X1  g0327(.A(KEYINPUT23), .B1(new_n204), .B2(G107), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT23), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(new_n223), .A3(G20), .ZN(new_n530));
  NAND2_X1  g0330(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n531));
  AND4_X1   g0331(.A1(new_n527), .A2(new_n528), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n524), .A2(new_n526), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n524), .A2(new_n534), .A3(new_n532), .A4(new_n526), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n450), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n259), .A2(G107), .ZN(new_n540));
  XNOR2_X1  g0340(.A(KEYINPUT84), .B(KEYINPUT25), .ZN(new_n541));
  XNOR2_X1  g0341(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n474), .A2(new_n223), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n273), .B(G264), .C1(new_n511), .C2(new_n508), .ZN(new_n545));
  MUX2_X1   g0345(.A(G250), .B(G257), .S(G1698), .Z(new_n546));
  AOI22_X1  g0346(.A1(new_n400), .A2(new_n546), .B1(G33), .B2(G294), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n510), .B(new_n545), .C1(new_n547), .C2(new_n273), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n548), .A2(new_n377), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(G190), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n539), .B(new_n544), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n484), .B1(new_n438), .B2(G107), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n476), .B1(new_n552), .B2(new_n450), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n518), .A2(new_n305), .A3(new_n519), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n342), .B1(new_n501), .B2(new_n513), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n521), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(G116), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n558), .B1(new_n203), .B2(G33), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n339), .A2(new_n559), .B1(new_n333), .B2(new_n558), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n489), .B(new_n204), .C1(G33), .C2(new_n480), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT20), .ZN(new_n562));
  AOI22_X1  g0362(.A1(KEYINPUT82), .A2(new_n562), .B1(new_n558), .B2(G20), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n563), .A3(new_n249), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(KEYINPUT82), .B2(new_n562), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n562), .A2(KEYINPUT82), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n561), .A2(new_n563), .A3(new_n249), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n560), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n273), .B(G270), .C1(new_n511), .C2(new_n508), .ZN(new_n570));
  NOR2_X1   g0370(.A1(G257), .A2(G1698), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n571), .B1(new_n224), .B2(G1698), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n400), .A2(new_n572), .B1(G303), .B2(new_n316), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n510), .B(new_n570), .C1(new_n573), .C2(new_n273), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n569), .A2(G169), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT21), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n342), .B1(new_n560), .B2(new_n568), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n578), .A2(KEYINPUT21), .A3(new_n574), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n400), .A2(new_n572), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n316), .A2(G303), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n273), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n510), .A2(new_n570), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n569), .A2(new_n584), .A3(G179), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n577), .A2(new_n579), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n544), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n538), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n545), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n400), .A2(new_n546), .ZN(new_n590));
  NAND2_X1  g0390(.A1(G33), .A2(G294), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n589), .B1(new_n592), .B2(new_n280), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(new_n305), .A3(new_n510), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n548), .A2(new_n342), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n588), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n586), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n330), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n367), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n400), .A2(new_n204), .A3(G68), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT19), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n251), .B2(new_n480), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n602), .B1(new_n352), .B2(new_n204), .ZN(new_n604));
  NOR4_X1   g0404(.A1(KEYINPUT81), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT81), .ZN(new_n606));
  NOR2_X1   g0406(.A1(G87), .A2(G97), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n606), .B1(new_n607), .B2(new_n223), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n604), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n601), .A2(new_n603), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n600), .B1(new_n610), .B2(new_n249), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n475), .A2(new_n599), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n502), .A2(new_n320), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n218), .B1(new_n276), .B2(G1), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(new_n273), .A3(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(G238), .A2(G1698), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n222), .B2(G1698), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n400), .A2(new_n618), .B1(G33), .B2(G116), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n616), .B1(new_n619), .B2(new_n273), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n342), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n425), .A2(new_n618), .A3(new_n313), .ZN(new_n622));
  NAND2_X1  g0422(.A1(G33), .A2(G116), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n273), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n616), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n305), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n613), .A2(new_n621), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n620), .A2(new_n295), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n362), .B(new_n616), .C1(new_n619), .C2(new_n273), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n474), .A2(new_n217), .ZN(new_n632));
  AOI211_X1 g0432(.A(new_n600), .B(new_n632), .C1(new_n610), .C2(new_n249), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n628), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n584), .A2(new_n377), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n574), .A2(new_n395), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n636), .A2(new_n637), .A3(new_n569), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  AND4_X1   g0439(.A1(new_n471), .A2(new_n557), .A3(new_n598), .A4(new_n639), .ZN(G372));
  NAND2_X1  g0440(.A1(new_n385), .A2(new_n376), .ZN(new_n641));
  INV_X1    g0441(.A(new_n379), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n344), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n459), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n304), .B1(new_n644), .B2(new_n468), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n645), .A2(new_n307), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n635), .A2(new_n556), .A3(new_n647), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n649));
  INV_X1    g0449(.A(new_n632), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n611), .A2(KEYINPUT85), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(KEYINPUT85), .B1(new_n611), .B2(new_n650), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n631), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n649), .A2(new_n653), .A3(new_n628), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n648), .B1(new_n647), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n653), .B1(new_n586), .B2(new_n597), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n521), .A2(new_n551), .A3(new_n556), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n628), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n646), .B1(new_n470), .B2(new_n659), .ZN(G369));
  NAND2_X1  g0460(.A1(new_n336), .A2(new_n204), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  OAI21_X1  g0466(.A(KEYINPUT86), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT86), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n664), .A2(new_n668), .A3(G343), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n569), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n586), .B(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G330), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n672), .A2(new_n673), .A3(new_n638), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n588), .A2(new_n596), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n670), .B1(new_n538), .B2(new_n587), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(new_n551), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n597), .A2(new_n670), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n680), .A2(KEYINPUT87), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(KEYINPUT87), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n667), .A2(new_n669), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n586), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n677), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n597), .B2(new_n685), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n684), .A2(new_n688), .ZN(G399));
  INV_X1    g0489(.A(new_n207), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OR3_X1    g0492(.A1(new_n605), .A2(new_n608), .A3(G116), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n692), .A2(G1), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n213), .B2(new_n692), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT88), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT29), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n685), .B1(new_n655), .B2(new_n658), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n699), .B1(new_n700), .B2(KEYINPUT90), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n611), .A2(new_n650), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT85), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n633), .A2(KEYINPUT85), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n704), .A2(new_n705), .B1(new_n629), .B2(new_n630), .ZN(new_n706));
  INV_X1    g0506(.A(new_n628), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n708), .A2(KEYINPUT26), .A3(new_n649), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n647), .B1(new_n635), .B2(new_n556), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT91), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI211_X1 g0512(.A(KEYINPUT91), .B(new_n647), .C1(new_n635), .C2(new_n556), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n709), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n685), .B1(new_n714), .B2(new_n658), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT90), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n700), .A2(new_n716), .ZN(new_n717));
  AOI22_X1  g0517(.A1(new_n701), .A2(new_n715), .B1(new_n717), .B2(new_n699), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n557), .A2(new_n598), .A3(new_n639), .A4(new_n685), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n584), .A2(new_n626), .A3(new_n593), .A4(G179), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n518), .A2(new_n519), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(KEYINPUT89), .B1(new_n624), .B2(new_n625), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT89), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n725), .B(new_n616), .C1(new_n619), .C2(new_n273), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n548), .A2(new_n574), .A3(new_n305), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(new_n728), .A3(new_n722), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n501), .A2(new_n513), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n574), .A2(new_n305), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n545), .B1(new_n547), .B2(new_n273), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n620), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n730), .A2(new_n731), .A3(new_n733), .A4(KEYINPUT30), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n723), .A2(new_n729), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n670), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT31), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n670), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n719), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G330), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n718), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n698), .B1(new_n743), .B2(G1), .ZN(G364));
  AOI21_X1  g0544(.A(new_n210), .B1(G20), .B2(new_n342), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n204), .A2(G190), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n298), .A2(new_n305), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n223), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n204), .A2(new_n305), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G200), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n395), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(G190), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n751), .A2(G50), .B1(new_n752), .B2(G68), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G179), .A2(G200), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n204), .B1(new_n754), .B2(G190), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G97), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n749), .A2(new_n377), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G190), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n753), .B(new_n757), .C1(new_n221), .C2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT32), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n746), .A2(new_n754), .ZN(new_n763));
  INV_X1    g0563(.A(G159), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n763), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n766), .A2(KEYINPUT32), .A3(G159), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n748), .B(new_n761), .C1(new_n765), .C2(new_n767), .ZN(new_n768));
  NOR4_X1   g0568(.A1(new_n295), .A2(new_n204), .A3(G179), .A4(new_n362), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n316), .B1(new_n769), .B2(G87), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT96), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n395), .A2(new_n758), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n772), .A2(KEYINPUT95), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(KEYINPUT95), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n768), .B(new_n771), .C1(new_n409), .C2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT97), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n769), .ZN(new_n779));
  INV_X1    g0579(.A(G303), .ZN(new_n780));
  INV_X1    g0580(.A(G283), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n779), .A2(new_n780), .B1(new_n781), .B2(new_n747), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n283), .B1(new_n766), .B2(G329), .ZN(new_n783));
  INV_X1    g0583(.A(G311), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n783), .B1(new_n760), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n752), .ZN(new_n786));
  XOR2_X1   g0586(.A(KEYINPUT33), .B(G317), .Z(new_n787));
  INV_X1    g0587(.A(G294), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n786), .A2(new_n787), .B1(new_n788), .B2(new_n755), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n782), .A2(new_n785), .A3(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G322), .ZN(new_n791));
  INV_X1    g0591(.A(G326), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n751), .B(KEYINPUT98), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n790), .B1(new_n791), .B2(new_n775), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n778), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n776), .A2(new_n777), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n745), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n335), .A2(G20), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n203), .B1(new_n798), .B2(G45), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n691), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n207), .A2(new_n283), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(KEYINPUT93), .B2(G355), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(KEYINPUT93), .B2(G355), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n246), .A2(new_n276), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n690), .A2(new_n400), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(G45), .B2(new_n213), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n805), .B1(G116), .B2(new_n207), .C1(new_n806), .C2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G13), .A2(G33), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(G20), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n745), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT94), .Z(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n802), .B1(new_n809), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n672), .A2(new_n638), .ZN(new_n817));
  INV_X1    g0617(.A(new_n812), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n797), .B(new_n816), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT92), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n674), .B(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n802), .B1(new_n817), .B2(G330), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n819), .B1(new_n821), .B2(new_n822), .ZN(G396));
  NAND3_X1  g0623(.A1(new_n345), .A2(new_n348), .A3(new_n685), .ZN(new_n824));
  AND3_X1   g0624(.A1(new_n577), .A2(new_n579), .A3(new_n585), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n706), .B1(new_n825), .B2(new_n675), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n707), .B1(new_n826), .B2(new_n557), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n654), .A2(new_n647), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n649), .A2(KEYINPUT26), .A3(new_n634), .A4(new_n628), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n824), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n685), .A2(new_n327), .A3(new_n341), .A4(new_n343), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n346), .A2(new_n347), .B1(new_n341), .B2(new_n670), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(new_n344), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n831), .B1(new_n700), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n801), .B1(new_n836), .B2(new_n741), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n836), .A2(new_n741), .ZN(new_n839));
  INV_X1    g0639(.A(new_n834), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n811), .ZN(new_n841));
  INV_X1    g0641(.A(new_n745), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n811), .ZN(new_n843));
  INV_X1    g0643(.A(new_n747), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(G87), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n283), .B1(new_n766), .B2(G311), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n845), .A2(new_n757), .A3(new_n846), .ZN(new_n847));
  AOI22_X1  g0647(.A1(G116), .A2(new_n759), .B1(new_n752), .B2(G283), .ZN(new_n848));
  INV_X1    g0648(.A(new_n751), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n848), .B1(new_n780), .B2(new_n849), .C1(new_n775), .C2(new_n788), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n847), .B(new_n850), .C1(G107), .C2(new_n769), .ZN(new_n851));
  INV_X1    g0651(.A(G132), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n400), .B1(new_n409), .B2(new_n755), .C1(new_n852), .C2(new_n763), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n844), .A2(G68), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n241), .B2(new_n779), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n751), .A2(G137), .B1(new_n759), .B2(G159), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n252), .B2(new_n786), .ZN(new_n857));
  INV_X1    g0657(.A(new_n775), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n857), .B1(new_n858), .B2(G143), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n853), .B(new_n855), .C1(new_n859), .C2(KEYINPUT34), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n859), .A2(KEYINPUT34), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n851), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n801), .B1(G77), .B2(new_n843), .C1(new_n862), .C2(new_n842), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT99), .Z(new_n864));
  OAI22_X1  g0664(.A1(new_n838), .A2(new_n839), .B1(new_n841), .B2(new_n864), .ZN(G384));
  NOR2_X1   g0665(.A1(new_n798), .A2(new_n203), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n646), .B1(new_n718), .B2(new_n470), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT103), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT39), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n460), .A2(new_n664), .ZN(new_n871));
  AND4_X1   g0671(.A1(new_n870), .A2(new_n464), .A3(new_n871), .A4(new_n441), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n449), .A2(new_n249), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n424), .A2(new_n429), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT16), .B1(new_n874), .B2(new_n454), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n408), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n664), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n463), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n877), .A2(new_n878), .A3(new_n441), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n872), .B1(new_n879), .B2(KEYINPUT37), .ZN(new_n880));
  INV_X1    g0680(.A(new_n467), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n466), .B1(new_n460), .B2(new_n463), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n445), .A2(new_n458), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n877), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n880), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n463), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n441), .B1(new_n457), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n890), .A2(KEYINPUT102), .A3(new_n870), .A4(new_n871), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n464), .A2(new_n871), .A3(new_n870), .A4(new_n441), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT102), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n457), .A2(new_n665), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT37), .B1(new_n889), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n891), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n895), .B1(new_n459), .B2(new_n468), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n869), .B1(new_n887), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n385), .A2(new_n376), .A3(new_n685), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n886), .B1(new_n880), .B2(new_n885), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n454), .B1(new_n447), .B2(new_n448), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n414), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n450), .B1(new_n874), .B2(new_n415), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n446), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n441), .B1(new_n907), .B2(new_n888), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n907), .A2(new_n665), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT37), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n892), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n909), .B1(new_n459), .B2(new_n468), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n911), .A2(KEYINPUT38), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n903), .A2(new_n913), .A3(KEYINPUT39), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n900), .A2(new_n902), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n903), .A2(new_n913), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n376), .A2(new_n670), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n641), .A2(new_n642), .A3(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n376), .B(new_n670), .C1(new_n385), .C2(new_n379), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n345), .A2(new_n348), .A3(new_n685), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n655), .B2(new_n658), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n832), .B(KEYINPUT101), .Z(new_n923));
  AOI21_X1  g0723(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n916), .A2(new_n924), .B1(new_n468), .B2(new_n665), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n915), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n868), .B(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n739), .A2(KEYINPUT104), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT104), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n735), .A2(new_n929), .A3(KEYINPUT31), .A4(new_n670), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n719), .A2(new_n928), .A3(new_n738), .A4(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n834), .B1(new_n918), .B2(new_n919), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT105), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n931), .A2(new_n932), .A3(KEYINPUT105), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT38), .B1(new_n911), .B2(new_n912), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n935), .B(new_n936), .C1(new_n887), .C2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT40), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AND3_X1   g0740(.A1(new_n931), .A2(new_n932), .A3(KEYINPUT40), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n887), .B2(new_n899), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n931), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n470), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n673), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n943), .B2(new_n945), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n866), .B1(new_n927), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n927), .B2(new_n947), .ZN(new_n949));
  INV_X1    g0749(.A(new_n483), .ZN(new_n950));
  OAI211_X1 g0750(.A(G116), .B(new_n211), .C1(new_n950), .C2(KEYINPUT35), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(KEYINPUT100), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(KEYINPUT35), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(KEYINPUT100), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT36), .ZN(new_n956));
  OAI21_X1  g0756(.A(G77), .B1(new_n409), .B2(new_n215), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n242), .B1(new_n957), .B2(new_n213), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n958), .A2(G1), .A3(new_n335), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n949), .A2(new_n956), .A3(new_n959), .ZN(G367));
  INV_X1    g0760(.A(G137), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n283), .B1(new_n961), .B2(new_n763), .C1(new_n786), .C2(new_n764), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n779), .A2(new_n409), .B1(new_n221), .B2(new_n747), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n760), .A2(new_n241), .B1(new_n755), .B2(new_n215), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(G143), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n965), .B1(new_n966), .B2(new_n793), .C1(new_n252), .C2(new_n775), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT46), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n769), .A2(G116), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n858), .A2(G303), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n970), .B1(new_n968), .B2(new_n969), .C1(new_n784), .C2(new_n793), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n747), .A2(new_n480), .ZN(new_n972));
  INV_X1    g0772(.A(G317), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n419), .B1(new_n973), .B2(new_n763), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n759), .A2(G283), .B1(G107), .B2(new_n756), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n975), .B(new_n976), .C1(new_n788), .C2(new_n786), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n967), .B1(new_n971), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n979));
  XNOR2_X1  g0779(.A(new_n978), .B(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n745), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n814), .B1(new_n690), .B2(new_n599), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n807), .A2(new_n236), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n802), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n704), .A2(new_n670), .A3(new_n705), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n708), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n628), .ZN(new_n987));
  OR3_X1    g0787(.A1(new_n986), .A2(KEYINPUT106), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(KEYINPUT106), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n981), .B(new_n984), .C1(new_n991), .C2(new_n818), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n521), .B(new_n556), .C1(new_n487), .C2(new_n685), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n649), .A2(new_n670), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n688), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT44), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n688), .A2(new_n995), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT45), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(new_n684), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n679), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n687), .B1(new_n1003), .B2(new_n686), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n821), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n674), .B2(new_n1004), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n742), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n691), .B(KEYINPUT41), .Z(new_n1008));
  OAI21_X1  g0808(.A(new_n799), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n687), .A2(new_n995), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1010), .A2(KEYINPUT42), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT107), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n993), .A2(new_n675), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n670), .B1(new_n1013), .B2(new_n556), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(KEYINPUT42), .B2(new_n1010), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1012), .A2(new_n1015), .B1(new_n991), .B2(KEYINPUT43), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n683), .A2(new_n995), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1021), .B(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT108), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1009), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1025), .B1(new_n1009), .B2(new_n1024), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n992), .B1(new_n1027), .B2(new_n1028), .ZN(G387));
  OAI21_X1  g0829(.A(new_n807), .B1(new_n233), .B2(new_n276), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n694), .B2(new_n803), .ZN(new_n1031));
  OR3_X1    g0831(.A1(new_n250), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1032));
  OAI21_X1  g0832(.A(KEYINPUT50), .B1(new_n250), .B2(G50), .ZN(new_n1033));
  AOI21_X1  g0833(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n694), .A2(new_n1032), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1031), .A2(new_n1035), .B1(new_n223), .B2(new_n690), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n801), .B1(new_n1036), .B2(new_n814), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n858), .A2(G50), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n769), .A2(G77), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n419), .B(new_n972), .C1(G150), .C2(new_n766), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n849), .A2(new_n764), .B1(new_n330), .B2(new_n755), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n250), .A2(new_n786), .B1(new_n760), .B2(new_n215), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .A4(new_n1043), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n769), .A2(G294), .B1(G283), .B2(new_n756), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G303), .A2(new_n759), .B1(new_n752), .B2(G311), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n793), .B2(new_n791), .C1(new_n973), .C2(new_n775), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT48), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1045), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT110), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT49), .Z(new_n1053));
  OAI221_X1 g0853(.A(new_n419), .B1(new_n792), .B2(new_n763), .C1(new_n747), .C2(new_n558), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT111), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1044), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1037), .B1(new_n1056), .B2(new_n745), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n1057), .A2(KEYINPUT112), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1057), .A2(KEYINPUT112), .B1(new_n1003), .B2(new_n812), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n1058), .A2(new_n1059), .B1(new_n800), .B2(new_n1006), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1006), .A2(new_n743), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1006), .A2(new_n743), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n691), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1060), .B1(new_n1061), .B2(new_n1063), .ZN(G393));
  INV_X1    g0864(.A(new_n1002), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n1062), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1062), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n692), .B1(new_n1002), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n807), .A2(new_n240), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n815), .B(new_n1070), .C1(new_n480), .C2(new_n207), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n802), .B1(new_n1071), .B2(KEYINPUT113), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(KEYINPUT113), .B2(new_n1071), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n756), .A2(G77), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1074), .B1(new_n760), .B2(new_n250), .C1(new_n241), .C2(new_n786), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1076), .A2(KEYINPUT114), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1076), .A2(KEYINPUT114), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n419), .B1(G143), .B2(new_n766), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n845), .B(new_n1079), .C1(new_n215), .C2(new_n779), .ZN(new_n1080));
  OR3_X1    g0880(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n775), .A2(new_n764), .B1(new_n252), .B2(new_n849), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT51), .Z(new_n1083));
  OAI22_X1  g0883(.A1(new_n775), .A2(new_n784), .B1(new_n973), .B2(new_n849), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT52), .Z(new_n1085));
  AOI21_X1  g0885(.A(new_n748), .B1(G283), .B2(new_n769), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n316), .B1(new_n763), .B2(new_n791), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G303), .B2(new_n752), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n759), .A2(G294), .B1(G116), .B2(new_n756), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1086), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n1081), .A2(new_n1083), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1073), .B1(new_n1091), .B2(new_n745), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n995), .B2(new_n818), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1069), .B(new_n1093), .C1(new_n799), .C2(new_n1065), .ZN(G390));
  OAI21_X1  g0894(.A(new_n896), .B1(new_n893), .B2(new_n892), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n892), .A2(new_n893), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n898), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n886), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n913), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n709), .A2(new_n712), .A3(new_n713), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n670), .B1(new_n1100), .B2(new_n827), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n833), .A2(new_n344), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1101), .A2(new_n1103), .B1(new_n344), .B2(new_n685), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1099), .B(new_n901), .C1(new_n920), .C2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n918), .A2(new_n919), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n740), .A2(G330), .A3(new_n1106), .A4(new_n840), .ZN(new_n1107));
  AOI21_X1  g0907(.A(KEYINPUT39), .B1(new_n1098), .B2(new_n913), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n903), .A2(KEYINPUT39), .A3(new_n913), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT115), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n924), .B2(new_n902), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n923), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1106), .B1(new_n831), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1114), .A2(KEYINPUT115), .A3(new_n901), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1105), .B(new_n1107), .C1(new_n1110), .C2(new_n1116), .ZN(new_n1117));
  NOR3_X1   g0917(.A1(new_n924), .A2(new_n1111), .A3(new_n902), .ZN(new_n1118));
  AOI21_X1  g0918(.A(KEYINPUT115), .B1(new_n1114), .B2(new_n901), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n900), .A2(new_n914), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1104), .A2(new_n920), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n902), .B1(new_n1098), .B2(new_n913), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1120), .A2(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n931), .A2(new_n932), .A3(G330), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1117), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n685), .B(new_n1103), .C1(new_n714), .C2(new_n658), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1127), .A2(new_n1107), .A3(new_n832), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n931), .A2(G330), .A3(new_n840), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n920), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n740), .A2(new_n840), .A3(G330), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n920), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n1125), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n922), .A2(new_n923), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1128), .A2(new_n1130), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n944), .A2(new_n673), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1136), .A2(new_n469), .A3(new_n390), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n646), .B(new_n1137), .C1(new_n718), .C2(new_n470), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1126), .A2(new_n1140), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1117), .B(new_n1139), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(new_n691), .A3(new_n1142), .ZN(new_n1143));
  OR2_X1    g0943(.A1(new_n1126), .A2(new_n799), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n801), .B1(new_n328), .B2(new_n843), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n858), .A2(G116), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n849), .A2(new_n781), .B1(new_n760), .B2(new_n480), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(G107), .B2(new_n752), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1074), .B(new_n316), .C1(new_n788), .C2(new_n763), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G87), .B2(new_n769), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1146), .A2(new_n854), .A3(new_n1148), .A4(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(G125), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT54), .B(G143), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n283), .B1(new_n763), .B2(new_n1152), .C1(new_n760), .C2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(G50), .B2(new_n844), .ZN(new_n1155));
  INV_X1    g0955(.A(G128), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n849), .A2(new_n1156), .B1(new_n764), .B2(new_n755), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G137), .B2(new_n752), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1155), .B(new_n1158), .C1(new_n852), .C2(new_n775), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n769), .A2(G150), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT53), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1151), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1145), .B1(new_n1162), .B2(new_n745), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n1110), .B2(new_n811), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1143), .A2(new_n1144), .A3(new_n1164), .ZN(G378));
  INV_X1    g0965(.A(new_n926), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n931), .A2(new_n932), .A3(KEYINPUT105), .ZN(new_n1167));
  AOI21_X1  g0967(.A(KEYINPUT105), .B1(new_n931), .B2(new_n932), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(KEYINPUT40), .B1(new_n1169), .B2(new_n916), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n942), .A2(G330), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n266), .A2(new_n664), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n304), .A2(new_n307), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1174), .B1(new_n304), .B2(new_n307), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1173), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1177), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(new_n1175), .A3(new_n1172), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1170), .A2(new_n1171), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1181), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n673), .B1(new_n1099), .B2(new_n941), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1183), .B1(new_n940), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1166), .B1(new_n1182), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1181), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n940), .A2(new_n1184), .A3(new_n1183), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n1188), .A3(new_n926), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n799), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1183), .A2(new_n810), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n801), .B1(G50), .B2(new_n843), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n747), .A2(new_n409), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1193), .A2(G41), .A3(new_n400), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1194), .B(new_n1039), .C1(new_n781), .C2(new_n763), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT116), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n759), .A2(new_n599), .B1(G68), .B2(new_n756), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1197), .B1(new_n480), .B2(new_n786), .C1(new_n558), .C2(new_n849), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G107), .B2(new_n858), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1196), .A2(new_n1199), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT117), .Z(new_n1201));
  OR2_X1    g1001(.A1(new_n1201), .A2(KEYINPUT58), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(KEYINPUT58), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(G33), .A2(G41), .ZN(new_n1204));
  AOI211_X1 g1004(.A(G50), .B(new_n1204), .C1(new_n419), .C2(new_n275), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n849), .A2(new_n1152), .B1(new_n760), .B2(new_n961), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n786), .A2(new_n852), .B1(new_n252), .B2(new_n755), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n779), .B2(new_n1153), .C1(new_n1156), .C2(new_n775), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1209), .A2(KEYINPUT59), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n766), .A2(G124), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1204), .B(new_n1211), .C1(new_n747), .C2(new_n764), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1209), .B2(KEYINPUT59), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1205), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1202), .A2(new_n1203), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1192), .B1(new_n1215), .B2(new_n745), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1190), .B1(new_n1191), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT118), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n926), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1220), .A2(KEYINPUT118), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1138), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1142), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(KEYINPUT57), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1222), .A2(new_n1225), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1142), .A2(new_n1223), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n691), .B1(new_n1227), .B2(KEYINPUT57), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1217), .B1(new_n1226), .B2(new_n1228), .ZN(G375));
  INV_X1    g1029(.A(new_n1008), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1140), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1135), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n920), .A2(new_n810), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n801), .B1(G68), .B2(new_n843), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n858), .A2(G137), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n769), .A2(G159), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n419), .B(new_n1193), .C1(G128), .C2(new_n766), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n849), .A2(new_n852), .B1(new_n760), .B2(new_n252), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n786), .A2(new_n1153), .B1(new_n241), .B2(new_n755), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .A4(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n858), .A2(G283), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n769), .A2(G97), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n849), .A2(new_n788), .B1(new_n760), .B2(new_n223), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G116), .B2(new_n752), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n316), .B1(new_n763), .B2(new_n780), .C1(new_n330), .C2(new_n755), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G77), .B2(new_n844), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1243), .A2(new_n1244), .A3(new_n1246), .A4(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1242), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1235), .B1(new_n1250), .B2(new_n745), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1233), .A2(new_n800), .B1(new_n1234), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1232), .A2(new_n1252), .ZN(new_n1253));
  XOR2_X1   g1053(.A(new_n1253), .B(KEYINPUT119), .Z(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(G381));
  INV_X1    g1055(.A(G384), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1093), .B1(new_n1065), .B2(new_n799), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1068), .B2(new_n1066), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(G393), .A2(G396), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1254), .A2(new_n1256), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  NOR4_X1   g1060(.A1(new_n1260), .A2(G387), .A3(G375), .A4(G378), .ZN(new_n1261));
  XOR2_X1   g1061(.A(new_n1261), .B(KEYINPUT120), .Z(G407));
  INV_X1    g1062(.A(G378), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n666), .ZN(new_n1264));
  OAI211_X1 g1064(.A(G407), .B(G213), .C1(G375), .C2(new_n1264), .ZN(G409));
  INV_X1    g1065(.A(G213), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1266), .A2(G343), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1142), .A2(new_n1223), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1187), .A2(new_n1188), .A3(new_n926), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1230), .B1(new_n1269), .B2(new_n1220), .ZN(new_n1270));
  OAI21_X1  g1070(.A(KEYINPUT121), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1191), .A2(new_n1216), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n800), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1008), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT121), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n1275), .A3(new_n1224), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .A4(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(KEYINPUT122), .A3(new_n1263), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G378), .B(new_n1217), .C1(new_n1226), .C2(new_n1228), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1277), .A2(new_n1263), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT122), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1267), .B1(new_n1280), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT126), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT60), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1233), .A2(new_n1223), .A3(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1287), .A2(new_n692), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1231), .B1(new_n1139), .B2(new_n1286), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(G384), .A3(new_n1252), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(G384), .B1(new_n1290), .B2(new_n1252), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1284), .A2(new_n1285), .A3(KEYINPUT63), .A4(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1267), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT122), .B1(new_n1277), .B2(new_n1263), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1294), .B(new_n1296), .C1(new_n1297), .C2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT63), .ZN(new_n1300));
  OAI21_X1  g1100(.A(KEYINPUT126), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1295), .A2(new_n1301), .ZN(new_n1302));
  XOR2_X1   g1102(.A(G393), .B(G396), .Z(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1009), .A2(new_n1024), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(KEYINPUT108), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1026), .ZN(new_n1307));
  AOI21_X1  g1107(.A(G390), .B1(new_n1307), .B2(new_n992), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n992), .ZN(new_n1309));
  AOI211_X1 g1109(.A(new_n1309), .B(new_n1258), .C1(new_n1306), .C2(new_n1026), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1304), .B1(new_n1308), .B2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT61), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(G387), .A2(new_n1258), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1307), .A2(new_n992), .A3(G390), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1313), .A2(new_n1314), .A3(new_n1303), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1311), .A2(new_n1312), .A3(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT125), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1267), .A2(G2897), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1294), .A2(new_n1318), .ZN(new_n1319));
  OAI211_X1 g1119(.A(G2897), .B(new_n1267), .C1(new_n1292), .C2(new_n1293), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1283), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1321), .B1(new_n1322), .B2(new_n1296), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1316), .B1(new_n1317), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1299), .A2(KEYINPUT123), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT123), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1322), .A2(new_n1326), .A3(new_n1294), .A4(new_n1296), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1325), .A2(new_n1327), .A3(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(KEYINPUT125), .B1(new_n1284), .B2(new_n1321), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1302), .A2(new_n1324), .A3(new_n1329), .A4(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1311), .A2(new_n1315), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1296), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1321), .ZN(new_n1334));
  AOI21_X1  g1134(.A(KEYINPUT62), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1299), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1312), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(KEYINPUT62), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1332), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1331), .A2(new_n1339), .ZN(G405));
  XNOR2_X1  g1140(.A(G375), .B(G378), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1294), .ZN(new_n1342));
  OR2_X1    g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT127), .ZN(new_n1345));
  OAI211_X1 g1145(.A(new_n1343), .B(new_n1344), .C1(new_n1345), .C2(new_n1332), .ZN(new_n1346));
  AOI21_X1  g1146(.A(KEYINPUT127), .B1(new_n1311), .B2(new_n1315), .ZN(new_n1347));
  XNOR2_X1  g1147(.A(new_n1346), .B(new_n1347), .ZN(G402));
endmodule


