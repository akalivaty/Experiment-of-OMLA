

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U546 ( .A(n755), .ZN(n733) );
  NOR2_X2 U547 ( .A1(G2105), .A2(G2104), .ZN(n530) );
  XNOR2_X1 U548 ( .A(n718), .B(n717), .ZN(n728) );
  NAND2_X1 U549 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U550 ( .A(KEYINPUT69), .B(n531), .Z(n532) );
  AND2_X1 U551 ( .A1(G1341), .A2(n755), .ZN(n513) );
  AND2_X1 U552 ( .A1(G125), .A2(n859), .ZN(n514) );
  XNOR2_X1 U553 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n717) );
  NOR2_X1 U554 ( .A1(n932), .A2(n513), .ZN(n727) );
  NOR2_X1 U555 ( .A1(G168), .A2(n749), .ZN(n750) );
  INV_X1 U556 ( .A(n711), .ZN(n716) );
  INV_X1 U557 ( .A(G2105), .ZN(n535) );
  XNOR2_X1 U558 ( .A(KEYINPUT15), .B(n604), .ZN(n933) );
  AND2_X1 U559 ( .A1(G2105), .A2(G2104), .ZN(n858) );
  NOR2_X1 U560 ( .A1(n645), .A2(G651), .ZN(n656) );
  NAND2_X1 U561 ( .A1(n540), .A2(n539), .ZN(n541) );
  INV_X1 U562 ( .A(G651), .ZN(n521) );
  NOR2_X1 U563 ( .A1(G543), .A2(n521), .ZN(n515) );
  XOR2_X1 U564 ( .A(KEYINPUT1), .B(n515), .Z(n649) );
  NAND2_X1 U565 ( .A1(G63), .A2(n649), .ZN(n517) );
  XOR2_X1 U566 ( .A(KEYINPUT0), .B(G543), .Z(n645) );
  NAND2_X1 U567 ( .A1(G51), .A2(n656), .ZN(n516) );
  NAND2_X1 U568 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U569 ( .A(KEYINPUT6), .B(n518), .ZN(n527) );
  NOR2_X1 U570 ( .A1(G543), .A2(G651), .ZN(n652) );
  NAND2_X1 U571 ( .A1(G89), .A2(n652), .ZN(n519) );
  XNOR2_X1 U572 ( .A(n519), .B(KEYINPUT76), .ZN(n520) );
  XNOR2_X1 U573 ( .A(n520), .B(KEYINPUT4), .ZN(n523) );
  NOR2_X2 U574 ( .A1(n645), .A2(n521), .ZN(n648) );
  NAND2_X1 U575 ( .A1(G76), .A2(n648), .ZN(n522) );
  NAND2_X1 U576 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U577 ( .A(KEYINPUT5), .B(n524), .ZN(n525) );
  XNOR2_X1 U578 ( .A(KEYINPUT77), .B(n525), .ZN(n526) );
  NOR2_X1 U579 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U580 ( .A(KEYINPUT7), .B(n528), .Z(G168) );
  NOR2_X1 U581 ( .A1(n535), .A2(G2104), .ZN(n529) );
  XNOR2_X2 U582 ( .A(n529), .B(KEYINPUT66), .ZN(n859) );
  XOR2_X2 U583 ( .A(KEYINPUT17), .B(n530), .Z(n862) );
  NAND2_X1 U584 ( .A1(n862), .A2(G137), .ZN(n533) );
  NAND2_X1 U585 ( .A1(G113), .A2(n858), .ZN(n531) );
  NOR2_X1 U586 ( .A1(n514), .A2(n534), .ZN(n540) );
  XOR2_X1 U587 ( .A(KEYINPUT68), .B(KEYINPUT23), .Z(n538) );
  NAND2_X1 U588 ( .A1(n535), .A2(G2104), .ZN(n536) );
  XNOR2_X2 U589 ( .A(n536), .B(KEYINPUT67), .ZN(n863) );
  NAND2_X1 U590 ( .A1(G101), .A2(n863), .ZN(n537) );
  XNOR2_X1 U591 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X2 U592 ( .A(n541), .B(KEYINPUT65), .ZN(G160) );
  XNOR2_X1 U593 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  INV_X1 U594 ( .A(G57), .ZN(G237) );
  NAND2_X1 U595 ( .A1(G132), .A2(G82), .ZN(n542) );
  XNOR2_X1 U596 ( .A(n542), .B(KEYINPUT22), .ZN(n543) );
  XNOR2_X1 U597 ( .A(n543), .B(KEYINPUT94), .ZN(n544) );
  NOR2_X1 U598 ( .A1(G218), .A2(n544), .ZN(n545) );
  NAND2_X1 U599 ( .A1(G96), .A2(n545), .ZN(n836) );
  NAND2_X1 U600 ( .A1(n836), .A2(G2106), .ZN(n549) );
  NAND2_X1 U601 ( .A1(G120), .A2(G69), .ZN(n546) );
  NOR2_X1 U602 ( .A1(G237), .A2(n546), .ZN(n547) );
  NAND2_X1 U603 ( .A1(G108), .A2(n547), .ZN(n835) );
  NAND2_X1 U604 ( .A1(G567), .A2(n835), .ZN(n548) );
  AND2_X1 U605 ( .A1(n549), .A2(n548), .ZN(G319) );
  XOR2_X1 U606 ( .A(G2443), .B(G2446), .Z(n551) );
  XNOR2_X1 U607 ( .A(G2427), .B(G2451), .ZN(n550) );
  XNOR2_X1 U608 ( .A(n551), .B(n550), .ZN(n557) );
  XOR2_X1 U609 ( .A(G2430), .B(G2454), .Z(n553) );
  XNOR2_X1 U610 ( .A(G1341), .B(G1348), .ZN(n552) );
  XNOR2_X1 U611 ( .A(n553), .B(n552), .ZN(n555) );
  XOR2_X1 U612 ( .A(G2435), .B(G2438), .Z(n554) );
  XNOR2_X1 U613 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U614 ( .A(n557), .B(n556), .Z(n558) );
  AND2_X1 U615 ( .A1(G14), .A2(n558), .ZN(G401) );
  NAND2_X1 U616 ( .A1(G123), .A2(n859), .ZN(n559) );
  XNOR2_X1 U617 ( .A(n559), .B(KEYINPUT18), .ZN(n561) );
  NAND2_X1 U618 ( .A1(G111), .A2(n858), .ZN(n560) );
  NAND2_X1 U619 ( .A1(n561), .A2(n560), .ZN(n565) );
  NAND2_X1 U620 ( .A1(G135), .A2(n862), .ZN(n563) );
  NAND2_X1 U621 ( .A1(G99), .A2(n863), .ZN(n562) );
  NAND2_X1 U622 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U623 ( .A1(n565), .A2(n564), .ZN(n917) );
  XNOR2_X1 U624 ( .A(n917), .B(G2096), .ZN(n566) );
  XNOR2_X1 U625 ( .A(n566), .B(KEYINPUT81), .ZN(n567) );
  OR2_X1 U626 ( .A1(G2100), .A2(n567), .ZN(G156) );
  NAND2_X1 U627 ( .A1(G64), .A2(n649), .ZN(n569) );
  NAND2_X1 U628 ( .A1(G52), .A2(n656), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n569), .A2(n568), .ZN(n574) );
  NAND2_X1 U630 ( .A1(G90), .A2(n652), .ZN(n571) );
  NAND2_X1 U631 ( .A1(G77), .A2(n648), .ZN(n570) );
  NAND2_X1 U632 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U633 ( .A(KEYINPUT9), .B(n572), .Z(n573) );
  NOR2_X1 U634 ( .A1(n574), .A2(n573), .ZN(G171) );
  INV_X1 U635 ( .A(G171), .ZN(G301) );
  NAND2_X1 U636 ( .A1(G88), .A2(n652), .ZN(n576) );
  NAND2_X1 U637 ( .A1(G75), .A2(n648), .ZN(n575) );
  NAND2_X1 U638 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U639 ( .A(KEYINPUT85), .B(n577), .ZN(n582) );
  NAND2_X1 U640 ( .A1(G62), .A2(n649), .ZN(n579) );
  NAND2_X1 U641 ( .A1(G50), .A2(n656), .ZN(n578) );
  NAND2_X1 U642 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U643 ( .A(KEYINPUT84), .B(n580), .Z(n581) );
  NAND2_X1 U644 ( .A1(n582), .A2(n581), .ZN(G303) );
  XOR2_X1 U645 ( .A(G168), .B(KEYINPUT8), .Z(n583) );
  XNOR2_X1 U646 ( .A(KEYINPUT78), .B(n583), .ZN(G286) );
  NAND2_X1 U647 ( .A1(G94), .A2(G452), .ZN(n584) );
  XNOR2_X1 U648 ( .A(n584), .B(KEYINPUT71), .ZN(G173) );
  NAND2_X1 U649 ( .A1(G7), .A2(G661), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n585), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U651 ( .A(G223), .B(KEYINPUT73), .ZN(n831) );
  NAND2_X1 U652 ( .A1(n831), .A2(G567), .ZN(n586) );
  XOR2_X1 U653 ( .A(KEYINPUT11), .B(n586), .Z(G234) );
  NAND2_X1 U654 ( .A1(G56), .A2(n649), .ZN(n587) );
  XOR2_X1 U655 ( .A(KEYINPUT14), .B(n587), .Z(n593) );
  NAND2_X1 U656 ( .A1(n652), .A2(G81), .ZN(n588) );
  XNOR2_X1 U657 ( .A(n588), .B(KEYINPUT12), .ZN(n590) );
  NAND2_X1 U658 ( .A1(G68), .A2(n648), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U660 ( .A(KEYINPUT13), .B(n591), .Z(n592) );
  NOR2_X1 U661 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U662 ( .A1(n656), .A2(G43), .ZN(n594) );
  NAND2_X1 U663 ( .A1(n595), .A2(n594), .ZN(n932) );
  INV_X1 U664 ( .A(G860), .ZN(n632) );
  NOR2_X1 U665 ( .A1(n932), .A2(n632), .ZN(n596) );
  XOR2_X1 U666 ( .A(KEYINPUT74), .B(n596), .Z(G153) );
  NAND2_X1 U667 ( .A1(G868), .A2(G301), .ZN(n606) );
  NAND2_X1 U668 ( .A1(n656), .A2(G54), .ZN(n603) );
  NAND2_X1 U669 ( .A1(G92), .A2(n652), .ZN(n598) );
  NAND2_X1 U670 ( .A1(G66), .A2(n649), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n598), .A2(n597), .ZN(n601) );
  NAND2_X1 U672 ( .A1(G79), .A2(n648), .ZN(n599) );
  XNOR2_X1 U673 ( .A(KEYINPUT75), .B(n599), .ZN(n600) );
  NOR2_X1 U674 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n603), .A2(n602), .ZN(n604) );
  INV_X1 U676 ( .A(n933), .ZN(n729) );
  INV_X1 U677 ( .A(G868), .ZN(n614) );
  NAND2_X1 U678 ( .A1(n729), .A2(n614), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n606), .A2(n605), .ZN(G284) );
  NAND2_X1 U680 ( .A1(G91), .A2(n652), .ZN(n608) );
  NAND2_X1 U681 ( .A1(G65), .A2(n649), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U683 ( .A1(G78), .A2(n648), .ZN(n610) );
  NAND2_X1 U684 ( .A1(G53), .A2(n656), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U686 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U687 ( .A(KEYINPUT72), .B(n613), .ZN(n943) );
  INV_X1 U688 ( .A(n943), .ZN(G299) );
  NAND2_X1 U689 ( .A1(G868), .A2(G286), .ZN(n616) );
  NAND2_X1 U690 ( .A1(G299), .A2(n614), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(G297) );
  NAND2_X1 U692 ( .A1(n632), .A2(G559), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n617), .A2(n933), .ZN(n618) );
  XNOR2_X1 U694 ( .A(n618), .B(KEYINPUT79), .ZN(n619) );
  XOR2_X1 U695 ( .A(KEYINPUT16), .B(n619), .Z(G148) );
  NAND2_X1 U696 ( .A1(n933), .A2(G868), .ZN(n620) );
  XNOR2_X1 U697 ( .A(KEYINPUT80), .B(n620), .ZN(n621) );
  NOR2_X1 U698 ( .A1(G559), .A2(n621), .ZN(n623) );
  NOR2_X1 U699 ( .A1(G868), .A2(n932), .ZN(n622) );
  NOR2_X1 U700 ( .A1(n623), .A2(n622), .ZN(G282) );
  NAND2_X1 U701 ( .A1(G93), .A2(n652), .ZN(n625) );
  NAND2_X1 U702 ( .A1(G80), .A2(n648), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n630) );
  NAND2_X1 U704 ( .A1(n649), .A2(G67), .ZN(n626) );
  XNOR2_X1 U705 ( .A(n626), .B(KEYINPUT82), .ZN(n628) );
  NAND2_X1 U706 ( .A1(G55), .A2(n656), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n671) );
  NAND2_X1 U709 ( .A1(G559), .A2(n933), .ZN(n631) );
  XOR2_X1 U710 ( .A(n932), .B(n631), .Z(n667) );
  NAND2_X1 U711 ( .A1(n632), .A2(n667), .ZN(n633) );
  XOR2_X1 U712 ( .A(n671), .B(n633), .Z(G145) );
  NAND2_X1 U713 ( .A1(G86), .A2(n652), .ZN(n635) );
  NAND2_X1 U714 ( .A1(G61), .A2(n649), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n648), .A2(G73), .ZN(n636) );
  XOR2_X1 U717 ( .A(KEYINPUT2), .B(n636), .Z(n637) );
  NOR2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U719 ( .A(KEYINPUT83), .B(n639), .Z(n641) );
  NAND2_X1 U720 ( .A1(n656), .A2(G48), .ZN(n640) );
  NAND2_X1 U721 ( .A1(n641), .A2(n640), .ZN(G305) );
  NAND2_X1 U722 ( .A1(G49), .A2(n656), .ZN(n643) );
  NAND2_X1 U723 ( .A1(G74), .A2(G651), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U725 ( .A1(n649), .A2(n644), .ZN(n647) );
  NAND2_X1 U726 ( .A1(n645), .A2(G87), .ZN(n646) );
  NAND2_X1 U727 ( .A1(n647), .A2(n646), .ZN(G288) );
  NAND2_X1 U728 ( .A1(G72), .A2(n648), .ZN(n651) );
  NAND2_X1 U729 ( .A1(G60), .A2(n649), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(n655) );
  NAND2_X1 U731 ( .A1(n652), .A2(G85), .ZN(n653) );
  XOR2_X1 U732 ( .A(KEYINPUT70), .B(n653), .Z(n654) );
  NOR2_X1 U733 ( .A1(n655), .A2(n654), .ZN(n658) );
  NAND2_X1 U734 ( .A1(n656), .A2(G47), .ZN(n657) );
  NAND2_X1 U735 ( .A1(n658), .A2(n657), .ZN(G290) );
  XOR2_X1 U736 ( .A(G303), .B(G305), .Z(n666) );
  XOR2_X1 U737 ( .A(KEYINPUT88), .B(KEYINPUT86), .Z(n659) );
  XNOR2_X1 U738 ( .A(G288), .B(n659), .ZN(n660) );
  XOR2_X1 U739 ( .A(n660), .B(KEYINPUT19), .Z(n662) );
  XOR2_X1 U740 ( .A(n943), .B(KEYINPUT87), .Z(n661) );
  XNOR2_X1 U741 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U742 ( .A(n671), .B(n663), .ZN(n664) );
  XNOR2_X1 U743 ( .A(n664), .B(G290), .ZN(n665) );
  XNOR2_X1 U744 ( .A(n666), .B(n665), .ZN(n877) );
  XNOR2_X1 U745 ( .A(n877), .B(n667), .ZN(n668) );
  XNOR2_X1 U746 ( .A(n668), .B(KEYINPUT89), .ZN(n669) );
  NAND2_X1 U747 ( .A1(n669), .A2(G868), .ZN(n670) );
  XOR2_X1 U748 ( .A(KEYINPUT90), .B(n670), .Z(n673) );
  NOR2_X1 U749 ( .A1(n671), .A2(G868), .ZN(n672) );
  NOR2_X1 U750 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U751 ( .A(KEYINPUT91), .B(n674), .ZN(G295) );
  NAND2_X1 U752 ( .A1(G2078), .A2(G2084), .ZN(n676) );
  XOR2_X1 U753 ( .A(KEYINPUT92), .B(KEYINPUT20), .Z(n675) );
  XNOR2_X1 U754 ( .A(n676), .B(n675), .ZN(n677) );
  NAND2_X1 U755 ( .A1(G2090), .A2(n677), .ZN(n678) );
  XNOR2_X1 U756 ( .A(KEYINPUT21), .B(n678), .ZN(n679) );
  NAND2_X1 U757 ( .A1(n679), .A2(G2072), .ZN(n680) );
  XOR2_X1 U758 ( .A(KEYINPUT93), .B(n680), .Z(G158) );
  NAND2_X1 U759 ( .A1(G661), .A2(G483), .ZN(n681) );
  XNOR2_X1 U760 ( .A(KEYINPUT95), .B(n681), .ZN(n682) );
  NAND2_X1 U761 ( .A1(n682), .A2(G319), .ZN(n683) );
  XOR2_X1 U762 ( .A(KEYINPUT96), .B(n683), .Z(n834) );
  NAND2_X1 U763 ( .A1(G36), .A2(n834), .ZN(G176) );
  NAND2_X1 U764 ( .A1(G138), .A2(n862), .ZN(n685) );
  NAND2_X1 U765 ( .A1(G102), .A2(n863), .ZN(n684) );
  NAND2_X1 U766 ( .A1(n685), .A2(n684), .ZN(n689) );
  NAND2_X1 U767 ( .A1(n858), .A2(G114), .ZN(n687) );
  NAND2_X1 U768 ( .A1(G126), .A2(n859), .ZN(n686) );
  NAND2_X1 U769 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U770 ( .A1(n689), .A2(n688), .ZN(G164) );
  XOR2_X1 U771 ( .A(KEYINPUT99), .B(G1991), .Z(n988) );
  NAND2_X1 U772 ( .A1(n858), .A2(G107), .ZN(n691) );
  NAND2_X1 U773 ( .A1(G119), .A2(n859), .ZN(n690) );
  NAND2_X1 U774 ( .A1(n691), .A2(n690), .ZN(n694) );
  NAND2_X1 U775 ( .A1(n862), .A2(G131), .ZN(n692) );
  XOR2_X1 U776 ( .A(KEYINPUT98), .B(n692), .Z(n693) );
  NOR2_X1 U777 ( .A1(n694), .A2(n693), .ZN(n696) );
  NAND2_X1 U778 ( .A1(n863), .A2(G95), .ZN(n695) );
  NAND2_X1 U779 ( .A1(n696), .A2(n695), .ZN(n846) );
  NAND2_X1 U780 ( .A1(n988), .A2(n846), .ZN(n697) );
  XNOR2_X1 U781 ( .A(n697), .B(KEYINPUT100), .ZN(n708) );
  NAND2_X1 U782 ( .A1(G105), .A2(n863), .ZN(n698) );
  XNOR2_X1 U783 ( .A(n698), .B(KEYINPUT38), .ZN(n705) );
  NAND2_X1 U784 ( .A1(n858), .A2(G117), .ZN(n700) );
  NAND2_X1 U785 ( .A1(G129), .A2(n859), .ZN(n699) );
  NAND2_X1 U786 ( .A1(n700), .A2(n699), .ZN(n703) );
  NAND2_X1 U787 ( .A1(G141), .A2(n862), .ZN(n701) );
  XNOR2_X1 U788 ( .A(KEYINPUT101), .B(n701), .ZN(n702) );
  NOR2_X1 U789 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U790 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U791 ( .A(KEYINPUT102), .B(n706), .ZN(n872) );
  NAND2_X1 U792 ( .A1(n872), .A2(G1996), .ZN(n707) );
  NAND2_X1 U793 ( .A1(n708), .A2(n707), .ZN(n923) );
  NOR2_X1 U794 ( .A1(G164), .A2(G1384), .ZN(n714) );
  NAND2_X1 U795 ( .A1(G160), .A2(G40), .ZN(n711) );
  NOR2_X1 U796 ( .A1(n714), .A2(n711), .ZN(n826) );
  NAND2_X1 U797 ( .A1(n923), .A2(n826), .ZN(n709) );
  XOR2_X1 U798 ( .A(n709), .B(KEYINPUT103), .Z(n810) );
  XNOR2_X1 U799 ( .A(G1986), .B(G290), .ZN(n937) );
  NAND2_X1 U800 ( .A1(n826), .A2(n937), .ZN(n710) );
  NAND2_X1 U801 ( .A1(n810), .A2(n710), .ZN(n798) );
  XOR2_X1 U802 ( .A(G2078), .B(KEYINPUT25), .Z(n983) );
  NAND2_X2 U803 ( .A1(n716), .A2(n714), .ZN(n755) );
  NOR2_X1 U804 ( .A1(n983), .A2(n755), .ZN(n713) );
  NOR2_X1 U805 ( .A1(n733), .A2(G1961), .ZN(n712) );
  NOR2_X1 U806 ( .A1(n713), .A2(n712), .ZN(n751) );
  OR2_X1 U807 ( .A1(n751), .A2(G301), .ZN(n746) );
  AND2_X1 U808 ( .A1(n727), .A2(n933), .ZN(n719) );
  AND2_X1 U809 ( .A1(G1996), .A2(n714), .ZN(n715) );
  NAND2_X1 U810 ( .A1(n716), .A2(n715), .ZN(n718) );
  NAND2_X1 U811 ( .A1(n719), .A2(n728), .ZN(n721) );
  INV_X1 U812 ( .A(KEYINPUT105), .ZN(n720) );
  XNOR2_X1 U813 ( .A(n721), .B(n720), .ZN(n726) );
  NAND2_X1 U814 ( .A1(n755), .A2(G1348), .ZN(n722) );
  XNOR2_X1 U815 ( .A(n722), .B(KEYINPUT106), .ZN(n724) );
  NAND2_X1 U816 ( .A1(n733), .A2(G2067), .ZN(n723) );
  NAND2_X1 U817 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U818 ( .A1(n726), .A2(n725), .ZN(n732) );
  NAND2_X1 U819 ( .A1(n728), .A2(n727), .ZN(n730) );
  NAND2_X1 U820 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U821 ( .A1(n732), .A2(n731), .ZN(n739) );
  NAND2_X1 U822 ( .A1(n733), .A2(G2072), .ZN(n734) );
  XNOR2_X1 U823 ( .A(KEYINPUT27), .B(n734), .ZN(n737) );
  NAND2_X1 U824 ( .A1(G1956), .A2(n755), .ZN(n735) );
  XOR2_X1 U825 ( .A(KEYINPUT104), .B(n735), .Z(n736) );
  NOR2_X1 U826 ( .A1(n737), .A2(n736), .ZN(n740) );
  NAND2_X1 U827 ( .A1(n740), .A2(n943), .ZN(n738) );
  NAND2_X1 U828 ( .A1(n739), .A2(n738), .ZN(n743) );
  NOR2_X1 U829 ( .A1(n740), .A2(n943), .ZN(n741) );
  XOR2_X1 U830 ( .A(n741), .B(KEYINPUT28), .Z(n742) );
  NAND2_X1 U831 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U832 ( .A(KEYINPUT29), .B(n744), .Z(n745) );
  NAND2_X1 U833 ( .A1(n746), .A2(n745), .ZN(n767) );
  NAND2_X2 U834 ( .A1(G8), .A2(n755), .ZN(n792) );
  NOR2_X1 U835 ( .A1(G1966), .A2(n792), .ZN(n770) );
  NOR2_X1 U836 ( .A1(G2084), .A2(n755), .ZN(n766) );
  NOR2_X1 U837 ( .A1(n770), .A2(n766), .ZN(n747) );
  NAND2_X1 U838 ( .A1(n747), .A2(G8), .ZN(n748) );
  XNOR2_X1 U839 ( .A(n748), .B(KEYINPUT30), .ZN(n749) );
  XNOR2_X1 U840 ( .A(n750), .B(KEYINPUT107), .ZN(n753) );
  NAND2_X1 U841 ( .A1(n751), .A2(G301), .ZN(n752) );
  NAND2_X1 U842 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U843 ( .A(KEYINPUT31), .B(n754), .ZN(n768) );
  NOR2_X1 U844 ( .A1(G1971), .A2(n792), .ZN(n757) );
  NOR2_X1 U845 ( .A1(G2090), .A2(n755), .ZN(n756) );
  NOR2_X1 U846 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U847 ( .A1(n758), .A2(G303), .ZN(n760) );
  AND2_X1 U848 ( .A1(n768), .A2(n760), .ZN(n759) );
  NAND2_X1 U849 ( .A1(n767), .A2(n759), .ZN(n763) );
  INV_X1 U850 ( .A(n760), .ZN(n761) );
  OR2_X1 U851 ( .A1(n761), .A2(G286), .ZN(n762) );
  AND2_X1 U852 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U853 ( .A1(n764), .A2(G8), .ZN(n765) );
  XNOR2_X1 U854 ( .A(n765), .B(KEYINPUT32), .ZN(n774) );
  NAND2_X1 U855 ( .A1(G8), .A2(n766), .ZN(n772) );
  AND2_X1 U856 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U857 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U858 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U859 ( .A1(n774), .A2(n773), .ZN(n788) );
  NOR2_X1 U860 ( .A1(G1976), .A2(G288), .ZN(n781) );
  NOR2_X1 U861 ( .A1(G1971), .A2(G303), .ZN(n775) );
  NOR2_X1 U862 ( .A1(n781), .A2(n775), .ZN(n950) );
  NAND2_X1 U863 ( .A1(n788), .A2(n950), .ZN(n778) );
  NAND2_X1 U864 ( .A1(G1976), .A2(G288), .ZN(n938) );
  INV_X1 U865 ( .A(n938), .ZN(n776) );
  NOR2_X1 U866 ( .A1(n792), .A2(n776), .ZN(n777) );
  AND2_X1 U867 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U868 ( .A1(KEYINPUT33), .A2(n779), .ZN(n780) );
  XNOR2_X1 U869 ( .A(n780), .B(KEYINPUT108), .ZN(n784) );
  NAND2_X1 U870 ( .A1(n781), .A2(KEYINPUT33), .ZN(n782) );
  NOR2_X1 U871 ( .A1(n792), .A2(n782), .ZN(n783) );
  NOR2_X1 U872 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U873 ( .A(G1981), .B(G305), .Z(n940) );
  NAND2_X1 U874 ( .A1(n785), .A2(n940), .ZN(n796) );
  NOR2_X1 U875 ( .A1(G2090), .A2(G303), .ZN(n786) );
  NAND2_X1 U876 ( .A1(G8), .A2(n786), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n789) );
  AND2_X1 U878 ( .A1(n789), .A2(n792), .ZN(n794) );
  NOR2_X1 U879 ( .A1(G1981), .A2(G305), .ZN(n790) );
  XOR2_X1 U880 ( .A(n790), .B(KEYINPUT24), .Z(n791) );
  NOR2_X1 U881 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n795) );
  AND2_X1 U883 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U884 ( .A1(n798), .A2(n797), .ZN(n809) );
  XNOR2_X1 U885 ( .A(G2067), .B(KEYINPUT37), .ZN(n823) );
  NAND2_X1 U886 ( .A1(G140), .A2(n862), .ZN(n800) );
  NAND2_X1 U887 ( .A1(G104), .A2(n863), .ZN(n799) );
  NAND2_X1 U888 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U889 ( .A(KEYINPUT34), .B(n801), .ZN(n806) );
  NAND2_X1 U890 ( .A1(n858), .A2(G116), .ZN(n803) );
  NAND2_X1 U891 ( .A1(G128), .A2(n859), .ZN(n802) );
  NAND2_X1 U892 ( .A1(n803), .A2(n802), .ZN(n804) );
  XOR2_X1 U893 ( .A(KEYINPUT35), .B(n804), .Z(n805) );
  NOR2_X1 U894 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U895 ( .A(KEYINPUT36), .B(n807), .ZN(n873) );
  NOR2_X1 U896 ( .A1(n823), .A2(n873), .ZN(n919) );
  NAND2_X1 U897 ( .A1(n919), .A2(n826), .ZN(n808) );
  XOR2_X1 U898 ( .A(KEYINPUT97), .B(n808), .Z(n821) );
  NAND2_X1 U899 ( .A1(n809), .A2(n821), .ZN(n829) );
  XOR2_X1 U900 ( .A(KEYINPUT113), .B(KEYINPUT39), .Z(n820) );
  NOR2_X1 U901 ( .A1(G1996), .A2(n872), .ZN(n914) );
  INV_X1 U902 ( .A(n810), .ZN(n816) );
  NOR2_X1 U903 ( .A1(n846), .A2(n988), .ZN(n811) );
  XNOR2_X1 U904 ( .A(n811), .B(KEYINPUT110), .ZN(n916) );
  NOR2_X1 U905 ( .A1(G1986), .A2(G290), .ZN(n812) );
  XOR2_X1 U906 ( .A(n812), .B(KEYINPUT109), .Z(n813) );
  NOR2_X1 U907 ( .A1(n916), .A2(n813), .ZN(n814) );
  XOR2_X1 U908 ( .A(KEYINPUT111), .B(n814), .Z(n815) );
  NOR2_X1 U909 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U910 ( .A(n817), .B(KEYINPUT112), .ZN(n818) );
  NOR2_X1 U911 ( .A1(n914), .A2(n818), .ZN(n819) );
  XNOR2_X1 U912 ( .A(n820), .B(n819), .ZN(n822) );
  NAND2_X1 U913 ( .A1(n822), .A2(n821), .ZN(n824) );
  NAND2_X1 U914 ( .A1(n823), .A2(n873), .ZN(n911) );
  NAND2_X1 U915 ( .A1(n824), .A2(n911), .ZN(n825) );
  NAND2_X1 U916 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U917 ( .A(n827), .B(KEYINPUT114), .ZN(n828) );
  NAND2_X1 U918 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U919 ( .A(n830), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n831), .ZN(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U922 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U924 ( .A1(n834), .A2(n833), .ZN(G188) );
  XNOR2_X1 U925 ( .A(G69), .B(KEYINPUT115), .ZN(G235) );
  INV_X1 U927 ( .A(G132), .ZN(G219) );
  INV_X1 U928 ( .A(G120), .ZN(G236) );
  INV_X1 U929 ( .A(G82), .ZN(G220) );
  NOR2_X1 U930 ( .A1(n836), .A2(n835), .ZN(G325) );
  INV_X1 U931 ( .A(G325), .ZN(G261) );
  NAND2_X1 U932 ( .A1(G112), .A2(n858), .ZN(n838) );
  NAND2_X1 U933 ( .A1(G100), .A2(n863), .ZN(n837) );
  NAND2_X1 U934 ( .A1(n838), .A2(n837), .ZN(n839) );
  XNOR2_X1 U935 ( .A(n839), .B(KEYINPUT117), .ZN(n841) );
  NAND2_X1 U936 ( .A1(G136), .A2(n862), .ZN(n840) );
  NAND2_X1 U937 ( .A1(n841), .A2(n840), .ZN(n844) );
  NAND2_X1 U938 ( .A1(n859), .A2(G124), .ZN(n842) );
  XOR2_X1 U939 ( .A(KEYINPUT44), .B(n842), .Z(n843) );
  NOR2_X1 U940 ( .A1(n844), .A2(n843), .ZN(G162) );
  XOR2_X1 U941 ( .A(G160), .B(n917), .Z(n845) );
  XNOR2_X1 U942 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U943 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n848) );
  XNOR2_X1 U944 ( .A(G164), .B(G162), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U946 ( .A(n850), .B(n849), .Z(n871) );
  NAND2_X1 U947 ( .A1(G139), .A2(n862), .ZN(n852) );
  NAND2_X1 U948 ( .A1(G103), .A2(n863), .ZN(n851) );
  NAND2_X1 U949 ( .A1(n852), .A2(n851), .ZN(n857) );
  NAND2_X1 U950 ( .A1(n858), .A2(G115), .ZN(n854) );
  NAND2_X1 U951 ( .A1(G127), .A2(n859), .ZN(n853) );
  NAND2_X1 U952 ( .A1(n854), .A2(n853), .ZN(n855) );
  XOR2_X1 U953 ( .A(KEYINPUT47), .B(n855), .Z(n856) );
  NOR2_X1 U954 ( .A1(n857), .A2(n856), .ZN(n906) );
  NAND2_X1 U955 ( .A1(n858), .A2(G118), .ZN(n861) );
  NAND2_X1 U956 ( .A1(G130), .A2(n859), .ZN(n860) );
  NAND2_X1 U957 ( .A1(n861), .A2(n860), .ZN(n868) );
  NAND2_X1 U958 ( .A1(G142), .A2(n862), .ZN(n865) );
  NAND2_X1 U959 ( .A1(G106), .A2(n863), .ZN(n864) );
  NAND2_X1 U960 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U961 ( .A(KEYINPUT45), .B(n866), .Z(n867) );
  NOR2_X1 U962 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U963 ( .A(n906), .B(n869), .ZN(n870) );
  XNOR2_X1 U964 ( .A(n871), .B(n870), .ZN(n875) );
  XOR2_X1 U965 ( .A(n873), .B(n872), .Z(n874) );
  XNOR2_X1 U966 ( .A(n875), .B(n874), .ZN(n876) );
  NOR2_X1 U967 ( .A1(G37), .A2(n876), .ZN(G395) );
  XNOR2_X1 U968 ( .A(n932), .B(n877), .ZN(n879) );
  XOR2_X1 U969 ( .A(G301), .B(n933), .Z(n878) );
  XNOR2_X1 U970 ( .A(n879), .B(n878), .ZN(n880) );
  XOR2_X1 U971 ( .A(n880), .B(G286), .Z(n881) );
  NOR2_X1 U972 ( .A1(G37), .A2(n881), .ZN(G397) );
  XNOR2_X1 U973 ( .A(G1956), .B(KEYINPUT41), .ZN(n891) );
  XOR2_X1 U974 ( .A(G1986), .B(G1976), .Z(n883) );
  XNOR2_X1 U975 ( .A(G1961), .B(G1971), .ZN(n882) );
  XNOR2_X1 U976 ( .A(n883), .B(n882), .ZN(n887) );
  XOR2_X1 U977 ( .A(G1991), .B(G1981), .Z(n885) );
  XNOR2_X1 U978 ( .A(G1966), .B(G1996), .ZN(n884) );
  XNOR2_X1 U979 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U980 ( .A(n887), .B(n886), .Z(n889) );
  XNOR2_X1 U981 ( .A(G2474), .B(KEYINPUT116), .ZN(n888) );
  XNOR2_X1 U982 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U983 ( .A(n891), .B(n890), .ZN(G229) );
  XOR2_X1 U984 ( .A(G2100), .B(G2096), .Z(n893) );
  XNOR2_X1 U985 ( .A(KEYINPUT42), .B(G2678), .ZN(n892) );
  XNOR2_X1 U986 ( .A(n893), .B(n892), .ZN(n897) );
  XOR2_X1 U987 ( .A(KEYINPUT43), .B(G2090), .Z(n895) );
  XNOR2_X1 U988 ( .A(G2072), .B(G2067), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U990 ( .A(n897), .B(n896), .Z(n899) );
  XNOR2_X1 U991 ( .A(G2078), .B(G2084), .ZN(n898) );
  XNOR2_X1 U992 ( .A(n899), .B(n898), .ZN(G227) );
  NOR2_X1 U993 ( .A1(G395), .A2(G397), .ZN(n900) );
  XNOR2_X1 U994 ( .A(n900), .B(KEYINPUT118), .ZN(n901) );
  NAND2_X1 U995 ( .A1(G319), .A2(n901), .ZN(n902) );
  NOR2_X1 U996 ( .A1(G401), .A2(n902), .ZN(n905) );
  NOR2_X1 U997 ( .A1(G229), .A2(G227), .ZN(n903) );
  XOR2_X1 U998 ( .A(KEYINPUT49), .B(n903), .Z(n904) );
  NAND2_X1 U999 ( .A1(n905), .A2(n904), .ZN(G225) );
  INV_X1 U1000 ( .A(G225), .ZN(G308) );
  INV_X1 U1001 ( .A(G303), .ZN(G166) );
  INV_X1 U1002 ( .A(G96), .ZN(G221) );
  INV_X1 U1003 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1004 ( .A(G2072), .B(n906), .Z(n908) );
  XOR2_X1 U1005 ( .A(G164), .B(G2078), .Z(n907) );
  NOR2_X1 U1006 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(KEYINPUT120), .B(n909), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n910), .B(KEYINPUT50), .ZN(n912) );
  NAND2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(n928) );
  XOR2_X1 U1010 ( .A(G2090), .B(G162), .Z(n913) );
  NOR2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(n915) );
  XOR2_X1 U1012 ( .A(KEYINPUT51), .B(n915), .Z(n925) );
  NOR2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(n921) );
  XOR2_X1 U1014 ( .A(G2084), .B(G160), .Z(n918) );
  NOR2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1016 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1017 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1018 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1019 ( .A(KEYINPUT119), .B(n926), .Z(n927) );
  NOR2_X1 U1020 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1021 ( .A(KEYINPUT52), .B(n929), .ZN(n930) );
  XNOR2_X1 U1022 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n999) );
  NAND2_X1 U1023 ( .A1(n930), .A2(n999), .ZN(n931) );
  NAND2_X1 U1024 ( .A1(n931), .A2(G29), .ZN(n1009) );
  XOR2_X1 U1025 ( .A(G16), .B(KEYINPUT56), .Z(n955) );
  XNOR2_X1 U1026 ( .A(G1341), .B(n932), .ZN(n953) );
  XNOR2_X1 U1027 ( .A(G1348), .B(n933), .ZN(n935) );
  NAND2_X1 U1028 ( .A1(G1971), .A2(G303), .ZN(n934) );
  NAND2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1030 ( .A1(n937), .A2(n936), .ZN(n939) );
  NAND2_X1 U1031 ( .A1(n939), .A2(n938), .ZN(n949) );
  XNOR2_X1 U1032 ( .A(G1966), .B(G168), .ZN(n941) );
  NAND2_X1 U1033 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1034 ( .A(n942), .B(KEYINPUT57), .ZN(n947) );
  XOR2_X1 U1035 ( .A(G171), .B(G1961), .Z(n945) );
  XOR2_X1 U1036 ( .A(n943), .B(G1956), .Z(n944) );
  NOR2_X1 U1037 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1038 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1039 ( .A1(n949), .A2(n948), .ZN(n951) );
  NAND2_X1 U1040 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1041 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1042 ( .A1(n955), .A2(n954), .ZN(n1006) );
  XOR2_X1 U1043 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n965) );
  XNOR2_X1 U1044 ( .A(G1956), .B(G20), .ZN(n957) );
  XNOR2_X1 U1045 ( .A(G19), .B(G1341), .ZN(n956) );
  NOR2_X1 U1046 ( .A1(n957), .A2(n956), .ZN(n963) );
  XOR2_X1 U1047 ( .A(KEYINPUT124), .B(G4), .Z(n959) );
  XNOR2_X1 U1048 ( .A(G1348), .B(KEYINPUT59), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(n959), .B(n958), .ZN(n961) );
  XNOR2_X1 U1050 ( .A(G1981), .B(G6), .ZN(n960) );
  NOR2_X1 U1051 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1052 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1053 ( .A(n965), .B(n964), .ZN(n978) );
  XNOR2_X1 U1054 ( .A(KEYINPUT123), .B(G1961), .ZN(n966) );
  XNOR2_X1 U1055 ( .A(n966), .B(G5), .ZN(n976) );
  XNOR2_X1 U1056 ( .A(G1971), .B(G22), .ZN(n968) );
  XNOR2_X1 U1057 ( .A(G23), .B(G1976), .ZN(n967) );
  NOR2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1059 ( .A(KEYINPUT126), .B(n969), .Z(n971) );
  XNOR2_X1 U1060 ( .A(G1986), .B(G24), .ZN(n970) );
  NOR2_X1 U1061 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1062 ( .A(KEYINPUT58), .B(n972), .Z(n974) );
  XNOR2_X1 U1063 ( .A(G1966), .B(G21), .ZN(n973) );
  NOR2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1065 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1066 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1067 ( .A(KEYINPUT61), .B(n979), .Z(n980) );
  NOR2_X1 U1068 ( .A1(G16), .A2(n980), .ZN(n1003) );
  XNOR2_X1 U1069 ( .A(G1996), .B(G32), .ZN(n982) );
  XNOR2_X1 U1070 ( .A(G26), .B(G2067), .ZN(n981) );
  NOR2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n987) );
  XNOR2_X1 U1072 ( .A(n983), .B(G27), .ZN(n985) );
  XNOR2_X1 U1073 ( .A(G2072), .B(G33), .ZN(n984) );
  NOR2_X1 U1074 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1075 ( .A1(n987), .A2(n986), .ZN(n992) );
  XOR2_X1 U1076 ( .A(n988), .B(G25), .Z(n989) );
  NAND2_X1 U1077 ( .A1(n989), .A2(G28), .ZN(n990) );
  XNOR2_X1 U1078 ( .A(KEYINPUT122), .B(n990), .ZN(n991) );
  NOR2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1080 ( .A(KEYINPUT53), .B(n993), .Z(n996) );
  XOR2_X1 U1081 ( .A(KEYINPUT54), .B(G34), .Z(n994) );
  XNOR2_X1 U1082 ( .A(G2084), .B(n994), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n998) );
  XNOR2_X1 U1084 ( .A(G35), .B(G2090), .ZN(n997) );
  NOR2_X1 U1085 ( .A1(n998), .A2(n997), .ZN(n1000) );
  XNOR2_X1 U1086 ( .A(n1000), .B(n999), .ZN(n1001) );
  NOR2_X1 U1087 ( .A1(G29), .A2(n1001), .ZN(n1002) );
  NOR2_X1 U1088 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1089 ( .A1(G11), .A2(n1004), .ZN(n1005) );
  NOR2_X1 U1090 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1091 ( .A(KEYINPUT127), .B(n1007), .Z(n1008) );
  NAND2_X1 U1092 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1093 ( .A(KEYINPUT62), .B(n1010), .ZN(G150) );
  INV_X1 U1094 ( .A(G150), .ZN(G311) );
endmodule

