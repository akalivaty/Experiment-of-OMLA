//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 1 0 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028;
  INV_X1    g000(.A(KEYINPUT96), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(KEYINPUT1), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n189), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT68), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n189), .A2(new_n191), .A3(new_n193), .A4(KEYINPUT68), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n198), .B1(new_n192), .B2(G146), .ZN(new_n199));
  NOR3_X1   g013(.A1(new_n190), .A2(KEYINPUT64), .A3(G143), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n191), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n188), .B1(new_n191), .B2(KEYINPUT1), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n196), .A2(new_n197), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G107), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT75), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT75), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G107), .ZN(new_n208));
  INV_X1    g022(.A(G104), .ZN(new_n209));
  AND3_X1   g023(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT78), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(new_n209), .B2(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n205), .A2(KEYINPUT78), .A3(G104), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(G101), .B1(new_n210), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(G107), .B1(new_n209), .B2(KEYINPUT3), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n209), .A2(KEYINPUT3), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n209), .A2(KEYINPUT3), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n207), .A2(G107), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n205), .A2(KEYINPUT75), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G101), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n218), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT80), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n215), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n225), .B1(new_n215), .B2(new_n224), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n204), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n191), .A2(new_n193), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  OR3_X1    g044(.A1(new_n230), .A2(new_n202), .A3(KEYINPUT79), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n196), .A2(new_n197), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT79), .B1(new_n230), .B2(new_n202), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n215), .A2(new_n224), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n228), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT11), .ZN(new_n239));
  INV_X1    g053(.A(G134), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(G137), .ZN(new_n241));
  INV_X1    g055(.A(G137), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT11), .A3(G134), .ZN(new_n243));
  INV_X1    g057(.A(G131), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n240), .A2(G137), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n241), .A2(new_n243), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT65), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n246), .B(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n241), .A2(new_n243), .A3(new_n245), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT66), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n241), .A2(new_n243), .A3(new_n251), .A4(new_n245), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(G131), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n248), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT12), .B1(new_n238), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT12), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n248), .A2(new_n253), .ZN(new_n257));
  AOI211_X1 g071(.A(new_n256), .B(new_n257), .C1(new_n228), .C2(new_n237), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT83), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n218), .A2(new_n222), .ZN(new_n260));
  XOR2_X1   g074(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(G101), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G104), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n265), .B1(new_n206), .B2(new_n208), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n216), .A2(new_n217), .ZN(new_n267));
  OAI21_X1  g081(.A(G101), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n224), .A2(new_n268), .A3(KEYINPUT4), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT76), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT76), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n224), .A2(new_n268), .A3(new_n271), .A4(KEYINPUT4), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n263), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(KEYINPUT0), .A2(G128), .ZN(new_n274));
  OR2_X1    g088(.A1(KEYINPUT0), .A2(G128), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n201), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  OR2_X1    g090(.A1(new_n229), .A2(new_n274), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT10), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n273), .A2(new_n278), .B1(new_n279), .B2(new_n237), .ZN(new_n280));
  INV_X1    g094(.A(new_n214), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n223), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n266), .A2(new_n267), .A3(G101), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT80), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n201), .A2(new_n203), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n279), .B1(new_n232), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n215), .A2(new_n224), .A3(new_n225), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT81), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n285), .A2(new_n287), .A3(KEYINPUT81), .A4(new_n288), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n280), .A2(new_n293), .A3(new_n257), .ZN(new_n294));
  INV_X1    g108(.A(G953), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G227), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n296), .B(KEYINPUT74), .ZN(new_n297));
  XNOR2_X1  g111(.A(G110), .B(G140), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n297), .B(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n232), .A2(new_n286), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n300), .B1(new_n285), .B2(new_n288), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n232), .A2(new_n233), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n235), .B1(new_n302), .B2(new_n231), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n254), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n256), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT83), .ZN(new_n306));
  OAI211_X1 g120(.A(KEYINPUT12), .B(new_n254), .C1(new_n301), .C2(new_n303), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n259), .A2(new_n294), .A3(new_n299), .A4(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT84), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n280), .A2(new_n293), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n254), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n294), .ZN(new_n314));
  INV_X1    g128(.A(new_n299), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n294), .A2(new_n299), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n317), .A2(KEYINPUT84), .A3(new_n259), .A4(new_n308), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n311), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G469), .ZN(new_n320));
  INV_X1    g134(.A(G902), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(G469), .A2(G902), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n317), .A2(KEYINPUT82), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n294), .A2(new_n299), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT82), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n324), .A2(new_n313), .A3(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n294), .B1(new_n258), .B2(new_n255), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n315), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(G469), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n322), .A2(new_n323), .A3(new_n331), .ZN(new_n332));
  XOR2_X1   g146(.A(KEYINPUT9), .B(G234), .Z(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(G221), .B1(new_n334), .B2(G902), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n295), .A2(G952), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n337), .B1(G234), .B2(G237), .ZN(new_n338));
  XOR2_X1   g152(.A(KEYINPUT21), .B(G898), .Z(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  AOI211_X1 g154(.A(new_n321), .B(new_n295), .C1(G234), .C2(G237), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n338), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(G237), .A2(G953), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(G143), .A3(G214), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(G143), .B1(new_n344), .B2(G214), .ZN(new_n347));
  OAI21_X1  g161(.A(G131), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n347), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n244), .A3(new_n345), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT17), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n348), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT91), .ZN(new_n353));
  XNOR2_X1  g167(.A(G125), .B(G140), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT16), .ZN(new_n355));
  INV_X1    g169(.A(G140), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G125), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n357), .A2(KEYINPUT16), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n355), .A2(G146), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(G146), .B1(new_n355), .B2(new_n358), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n349), .A2(new_n345), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(KEYINPUT17), .A3(G131), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT91), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n348), .A2(new_n350), .A3(new_n365), .A4(new_n351), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n353), .A2(new_n362), .A3(new_n364), .A4(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(G113), .B(G122), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(new_n209), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n363), .A2(KEYINPUT18), .A3(G131), .ZN(new_n370));
  INV_X1    g184(.A(G125), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G140), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n357), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G146), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n354), .A2(new_n190), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT90), .ZN(new_n376));
  OR2_X1    g190(.A1(new_n374), .A2(KEYINPUT90), .ZN(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT18), .A2(G131), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n349), .A2(new_n345), .A3(new_n378), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n370), .A2(new_n376), .A3(new_n377), .A4(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n367), .A2(new_n369), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n369), .B1(new_n367), .B2(new_n380), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n321), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G475), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n354), .B(KEYINPUT19), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n190), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n348), .A2(new_n350), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(new_n359), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n380), .ZN(new_n390));
  INV_X1    g204(.A(new_n369), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(G475), .B1(new_n381), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n321), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(KEYINPUT20), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n397), .B1(new_n393), .B2(new_n321), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n343), .B(new_n385), .C1(new_n395), .C2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G478), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(KEYINPUT15), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT95), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n333), .A2(G217), .A3(new_n295), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT92), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n188), .B2(G143), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n192), .A2(KEYINPUT92), .A3(G128), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT93), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n408), .B1(new_n188), .B2(G143), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n192), .A2(KEYINPUT93), .A3(G128), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n406), .B(new_n407), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n409), .A2(new_n410), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n411), .B(G134), .C1(new_n412), .C2(KEYINPUT13), .ZN(new_n413));
  OR2_X1    g227(.A1(new_n409), .A2(new_n410), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n406), .A2(new_n407), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT13), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n414), .B(new_n415), .C1(new_n416), .C2(new_n240), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n206), .A2(new_n208), .ZN(new_n418));
  XNOR2_X1  g232(.A(G116), .B(G122), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n418), .B(new_n419), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n413), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT14), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G122), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(G116), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n205), .B1(new_n425), .B2(KEYINPUT14), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n423), .A2(new_n426), .B1(new_n418), .B2(new_n419), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n240), .B1(new_n414), .B2(new_n415), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n411), .A2(G134), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT94), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n427), .B(KEYINPUT94), .C1(new_n428), .C2(new_n429), .ZN(new_n433));
  AOI211_X1 g247(.A(new_n404), .B(new_n421), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n404), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n433), .ZN(new_n436));
  INV_X1    g250(.A(new_n421), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n403), .B1(new_n439), .B2(G902), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n436), .A2(new_n437), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n404), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n436), .A2(new_n437), .A3(new_n435), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(KEYINPUT95), .A3(new_n321), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n402), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n439), .A2(G902), .A3(new_n401), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n399), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(G214), .B1(G237), .B2(G902), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n270), .A2(new_n272), .ZN(new_n450));
  XOR2_X1   g264(.A(KEYINPUT2), .B(G113), .Z(new_n451));
  XNOR2_X1  g265(.A(G116), .B(G119), .ZN(new_n452));
  OR2_X1    g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n452), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT69), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n453), .A2(KEYINPUT69), .A3(new_n454), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n450), .A2(new_n262), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT85), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n452), .A2(KEYINPUT5), .ZN(new_n462));
  INV_X1    g276(.A(G119), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(G116), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n462), .B(G113), .C1(KEYINPUT5), .C2(new_n464), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n285), .A2(new_n288), .A3(new_n454), .A4(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT85), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n273), .A2(new_n467), .A3(new_n459), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n461), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(G110), .B(G122), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n461), .A2(new_n470), .A3(new_n466), .A4(new_n468), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(KEYINPUT6), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n371), .B1(new_n276), .B2(new_n277), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT86), .B1(new_n300), .B2(G125), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT86), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n204), .A2(new_n477), .A3(new_n371), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n475), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G224), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(G953), .ZN(new_n481));
  XOR2_X1   g295(.A(new_n479), .B(new_n481), .Z(new_n482));
  INV_X1    g296(.A(KEYINPUT6), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n469), .A2(new_n483), .A3(new_n471), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n474), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(G210), .B1(G237), .B2(G902), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n476), .A2(new_n478), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT87), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT87), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n476), .A2(new_n489), .A3(new_n478), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  XOR2_X1   g305(.A(KEYINPUT88), .B(KEYINPUT7), .Z(new_n492));
  OAI22_X1  g306(.A1(new_n491), .A2(new_n475), .B1(new_n481), .B2(new_n492), .ZN(new_n493));
  XOR2_X1   g307(.A(new_n470), .B(KEYINPUT8), .Z(new_n494));
  NAND2_X1  g308(.A1(new_n465), .A2(new_n454), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n235), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n494), .B1(new_n466), .B2(new_n496), .ZN(new_n497));
  AOI211_X1 g311(.A(new_n481), .B(new_n475), .C1(new_n476), .C2(new_n478), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n497), .B1(new_n498), .B2(KEYINPUT7), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n493), .A2(new_n473), .A3(new_n499), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n500), .A2(new_n321), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n485), .A2(new_n486), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n486), .B1(new_n485), .B2(new_n501), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n448), .B(new_n449), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n187), .B1(new_n336), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n504), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n506), .A2(KEYINPUT96), .A3(new_n335), .A4(new_n332), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT32), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n344), .A2(G210), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(new_n223), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n511));
  XOR2_X1   g325(.A(new_n510), .B(new_n511), .Z(new_n512));
  NAND2_X1  g326(.A1(new_n254), .A2(new_n278), .ZN(new_n513));
  OR2_X1    g327(.A1(new_n246), .A2(new_n247), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n246), .A2(new_n247), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n242), .A2(G134), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n245), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n514), .A2(new_n515), .B1(G131), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n300), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n453), .A2(KEYINPUT69), .A3(new_n454), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT69), .B1(new_n453), .B2(new_n454), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n513), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT70), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT28), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n524), .B1(new_n523), .B2(new_n525), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT67), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n204), .B1(new_n518), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n517), .A2(G131), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n248), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT67), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n522), .B1(new_n535), .B2(new_n513), .ZN(new_n536));
  INV_X1    g350(.A(new_n523), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT28), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n512), .B1(new_n529), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT30), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n540), .B1(new_n513), .B2(new_n519), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n531), .A2(new_n534), .B1(new_n254), .B2(new_n278), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n541), .B1(new_n542), .B2(new_n540), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n523), .B(new_n512), .C1(new_n543), .C2(new_n522), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT31), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n300), .B1(new_n533), .B2(KEYINPUT67), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n518), .A2(new_n530), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n540), .B(new_n513), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n541), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n537), .B1(new_n551), .B2(new_n459), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(KEYINPUT31), .A3(new_n512), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n539), .B1(new_n546), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(G472), .A2(G902), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n508), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n512), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n513), .B1(new_n547), .B2(new_n548), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n459), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n525), .B1(new_n560), .B2(new_n523), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n523), .A2(new_n525), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT70), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n526), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n558), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT31), .B1(new_n552), .B2(new_n512), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n522), .B1(new_n549), .B2(new_n550), .ZN(new_n567));
  NOR4_X1   g381(.A1(new_n567), .A2(new_n545), .A3(new_n537), .A4(new_n558), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n565), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(KEYINPUT32), .A3(new_n555), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n512), .B1(new_n561), .B2(new_n564), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n552), .A2(new_n558), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT29), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n513), .A2(new_n519), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n459), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n575), .A2(new_n523), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n526), .B(new_n563), .C1(new_n576), .C2(new_n525), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n512), .A2(KEYINPUT29), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n321), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(G472), .B1(new_n573), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n557), .A2(new_n570), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(G217), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n582), .B1(G234), .B2(new_n321), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT23), .B1(new_n188), .B2(G119), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n188), .A2(G119), .ZN(new_n585));
  MUX2_X1   g399(.A(KEYINPUT23), .B(new_n584), .S(new_n585), .Z(new_n586));
  XNOR2_X1  g400(.A(G119), .B(G128), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT24), .B(G110), .Z(new_n588));
  OAI22_X1  g402(.A1(new_n586), .A2(G110), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n589), .A2(new_n359), .A3(new_n375), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n586), .A2(G110), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n588), .A2(new_n587), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n591), .B(new_n592), .C1(new_n360), .C2(new_n361), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n295), .A2(G221), .A3(G234), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT71), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT22), .B(G137), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n594), .B(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT25), .B1(new_n600), .B2(new_n321), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n594), .A2(new_n599), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n598), .B1(new_n590), .B2(new_n593), .ZN(new_n603));
  OAI211_X1 g417(.A(KEYINPUT25), .B(new_n321), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n583), .B1(new_n601), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT72), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI211_X1 g422(.A(KEYINPUT72), .B(new_n583), .C1(new_n601), .C2(new_n605), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n583), .A2(G902), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT73), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n610), .B1(new_n600), .B2(new_n613), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n581), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n505), .A2(new_n507), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(G101), .ZN(G3));
  INV_X1    g431(.A(new_n614), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n336), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(G472), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n569), .B2(new_n321), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n555), .B2(new_n569), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n502), .A2(new_n503), .ZN(new_n625));
  INV_X1    g439(.A(new_n449), .ZN(new_n626));
  AOI21_X1  g440(.A(KEYINPUT95), .B1(new_n444), .B2(new_n321), .ZN(new_n627));
  AOI211_X1 g441(.A(new_n403), .B(G902), .C1(new_n442), .C2(new_n443), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n400), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n442), .A2(KEYINPUT33), .A3(new_n443), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT33), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n631), .B1(new_n434), .B2(new_n438), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n630), .A2(new_n632), .A3(G478), .A4(new_n321), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n385), .B1(new_n395), .B2(new_n398), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR4_X1   g450(.A1(new_n625), .A2(new_n626), .A3(new_n342), .A4(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n624), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT34), .B(G104), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT97), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n638), .B(new_n640), .ZN(G6));
  NAND2_X1  g455(.A1(new_n485), .A2(new_n501), .ZN(new_n642));
  INV_X1    g456(.A(new_n486), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n485), .A2(new_n486), .A3(new_n501), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n646), .A2(new_n449), .A3(new_n343), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n446), .A2(new_n447), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n394), .B(new_n396), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n385), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n624), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  NOR2_X1   g468(.A1(new_n598), .A2(KEYINPUT36), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n594), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n613), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n608), .A2(new_n609), .A3(new_n657), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n622), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n505), .A2(new_n507), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT37), .B(G110), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  AND2_X1   g476(.A1(new_n332), .A2(new_n335), .ZN(new_n663));
  INV_X1    g477(.A(new_n338), .ZN(new_n664));
  INV_X1    g478(.A(new_n341), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n664), .B1(new_n665), .B2(G900), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n649), .A2(new_n385), .A3(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n648), .A2(new_n667), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n449), .B(new_n658), .C1(new_n502), .C2(new_n503), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n663), .A2(new_n581), .A3(new_n668), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  XNOR2_X1  g486(.A(new_n666), .B(KEYINPUT39), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n663), .A2(new_n673), .ZN(new_n674));
  OR2_X1    g488(.A1(new_n674), .A2(KEYINPUT40), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT38), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n676), .B1(new_n502), .B2(new_n503), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n644), .A2(KEYINPUT38), .A3(new_n645), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n635), .B(new_n449), .C1(new_n446), .C2(new_n447), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n512), .B1(new_n567), .B2(new_n537), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT98), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n576), .A2(new_n558), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n321), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n683), .B1(new_n682), .B2(new_n684), .ZN(new_n687));
  OAI21_X1  g501(.A(G472), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n557), .A2(new_n688), .A3(new_n570), .ZN(new_n689));
  INV_X1    g503(.A(new_n658), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n674), .A2(KEYINPUT40), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n675), .A2(new_n681), .A3(new_n691), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G143), .ZN(G45));
  AOI21_X1  g508(.A(G478), .B1(new_n440), .B2(new_n445), .ZN(new_n695));
  INV_X1    g509(.A(new_n633), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n635), .B(new_n666), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT99), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n634), .A2(KEYINPUT99), .A3(new_n635), .A4(new_n666), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n663), .A2(new_n581), .A3(new_n670), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  INV_X1    g518(.A(KEYINPUT101), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT100), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n320), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n319), .A2(new_n321), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n708), .B1(new_n319), .B2(new_n321), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n705), .B1(new_n711), .B2(new_n335), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n319), .A2(new_n321), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n707), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n319), .A2(new_n321), .A3(new_n708), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n714), .A2(new_n705), .A3(new_n715), .A4(new_n335), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT102), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n718), .A2(new_n719), .A3(new_n615), .A4(new_n637), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n714), .A2(new_n335), .A3(new_n715), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT101), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n722), .A2(new_n637), .A3(new_n615), .A4(new_n716), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(KEYINPUT102), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT41), .B(G113), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G15));
  NAND3_X1  g541(.A1(new_n718), .A2(new_n615), .A3(new_n651), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G116), .ZN(G18));
  AND2_X1   g543(.A1(new_n581), .A2(new_n448), .ZN(new_n730));
  AND4_X1   g544(.A1(new_n670), .A2(new_n722), .A3(new_n716), .A4(new_n730), .ZN(new_n731));
  XOR2_X1   g545(.A(KEYINPUT103), .B(G119), .Z(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G21));
  INV_X1    g547(.A(new_n680), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n646), .A2(new_n343), .A3(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n577), .A2(new_n558), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n737), .B1(new_n566), .B2(new_n568), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n555), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n546), .A2(new_n553), .ZN(new_n740));
  AOI21_X1  g554(.A(G902), .B1(new_n740), .B2(new_n565), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n739), .B1(new_n741), .B2(new_n620), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n618), .A2(new_n742), .ZN(new_n743));
  AND4_X1   g557(.A1(new_n716), .A2(new_n722), .A3(new_n736), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n424), .ZN(G24));
  NOR2_X1   g559(.A1(new_n625), .A2(new_n626), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n739), .B(new_n658), .C1(new_n741), .C2(new_n620), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n701), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n722), .A2(new_n746), .A3(new_n748), .A4(new_n716), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G125), .ZN(G27));
  INV_X1    g564(.A(KEYINPUT42), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n330), .A2(KEYINPUT104), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n330), .A2(KEYINPUT104), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n328), .B(G469), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n322), .A2(new_n754), .A3(new_n323), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n755), .A2(new_n335), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n644), .A2(new_n449), .A3(new_n645), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT105), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n644), .A2(KEYINPUT105), .A3(new_n449), .A4(new_n645), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n756), .A2(new_n615), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n751), .B1(new_n761), .B2(new_n701), .ZN(new_n762));
  AND4_X1   g576(.A1(new_n335), .A2(new_n759), .A3(new_n755), .A4(new_n760), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n763), .A2(KEYINPUT42), .A3(new_n615), .A4(new_n702), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G131), .ZN(G33));
  AOI21_X1  g580(.A(KEYINPUT105), .B1(new_n625), .B2(new_n449), .ZN(new_n767));
  INV_X1    g581(.A(new_n760), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n769), .A2(new_n615), .A3(new_n668), .A4(new_n756), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G134), .ZN(G36));
  OAI211_X1 g585(.A(new_n328), .B(KEYINPUT45), .C1(new_n752), .C2(new_n753), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n328), .A2(new_n330), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n772), .B(G469), .C1(new_n773), .C2(KEYINPUT45), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(KEYINPUT46), .A3(new_n323), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n322), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT46), .B1(new_n774), .B2(new_n323), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n335), .A3(new_n673), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  INV_X1    g594(.A(new_n635), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n634), .A2(new_n781), .ZN(new_n782));
  XOR2_X1   g596(.A(new_n782), .B(KEYINPUT43), .Z(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  OR3_X1    g598(.A1(new_n784), .A2(new_n622), .A3(new_n690), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n779), .B1(new_n780), .B2(new_n785), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n786), .B(new_n769), .C1(new_n780), .C2(new_n785), .ZN(new_n787));
  XNOR2_X1  g601(.A(KEYINPUT106), .B(G137), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(G39));
  NAND2_X1  g603(.A1(new_n778), .A2(new_n335), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT47), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(KEYINPUT107), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(KEYINPUT107), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n792), .B1(new_n790), .B2(new_n794), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n793), .A2(new_n795), .A3(new_n581), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(new_n618), .A3(new_n702), .A4(new_n769), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  OR2_X1    g612(.A1(G952), .A2(G953), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n449), .B1(new_n677), .B2(new_n678), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n722), .A2(new_n716), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT115), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n783), .A2(new_n338), .A3(new_n743), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n722), .A2(new_n800), .A3(new_n804), .A4(new_n716), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n802), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT117), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n718), .A2(new_n338), .A3(new_n769), .A4(new_n783), .ZN(new_n811));
  OAI21_X1  g625(.A(KEYINPUT118), .B1(new_n811), .B2(new_n747), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n759), .A2(new_n760), .ZN(new_n813));
  NOR4_X1   g627(.A1(new_n712), .A2(new_n813), .A3(new_n717), .A4(new_n664), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n815));
  INV_X1    g629(.A(new_n747), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n814), .A2(new_n815), .A3(new_n816), .A4(new_n783), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n809), .B1(new_n806), .B2(KEYINPUT117), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n810), .B(new_n818), .C1(new_n820), .C2(new_n808), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n718), .A2(new_n338), .A3(new_n769), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n822), .A2(new_n618), .A3(new_n689), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n634), .A2(new_n635), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT119), .B1(new_n821), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n808), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n828), .A2(new_n819), .B1(new_n817), .B2(new_n812), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(new_n825), .A3(new_n830), .A4(new_n810), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n833));
  INV_X1    g647(.A(new_n711), .ZN(new_n834));
  OAI22_X1  g648(.A1(new_n793), .A2(new_n795), .B1(new_n335), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n803), .A2(new_n769), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n833), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT120), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n832), .A2(new_n840), .A3(new_n837), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n625), .A2(new_n680), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n756), .A2(new_n691), .A3(new_n666), .A4(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n749), .A3(new_n671), .A4(new_n703), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n846), .B(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT112), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT53), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI211_X1 g664(.A(new_n731), .B(new_n744), .C1(new_n720), .C2(new_n724), .ZN(new_n851));
  INV_X1    g665(.A(new_n616), .ZN(new_n852));
  OR3_X1    g666(.A1(new_n446), .A2(KEYINPUT109), .A3(new_n447), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT109), .B1(new_n446), .B2(new_n447), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n853), .A2(new_n781), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n647), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n619), .A2(new_n856), .A3(new_n622), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n660), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n852), .B1(new_n858), .B2(KEYINPUT110), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT110), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n660), .A2(new_n860), .A3(new_n857), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n861), .A2(new_n638), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n851), .A2(new_n728), .A3(new_n859), .A4(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n690), .A2(new_n667), .ZN(new_n864));
  AND4_X1   g678(.A1(new_n335), .A2(new_n332), .A3(new_n581), .A4(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT111), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n853), .A2(new_n854), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n769), .A2(new_n865), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n759), .A2(new_n760), .A3(new_n867), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n332), .A2(new_n581), .A3(new_n864), .A4(new_n335), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT111), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n868), .A2(new_n770), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n762), .B2(new_n764), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n749), .A2(new_n671), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n847), .A3(new_n703), .A4(new_n845), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n846), .A2(KEYINPUT52), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n763), .A2(new_n748), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n873), .A2(new_n875), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n850), .B1(new_n863), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n875), .A2(new_n876), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n880), .B1(new_n881), .B2(KEYINPUT112), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n858), .A2(KEYINPUT110), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n883), .A2(new_n616), .A3(new_n638), .A4(new_n861), .ZN(new_n884));
  INV_X1    g698(.A(new_n731), .ZN(new_n885));
  INV_X1    g699(.A(new_n744), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n725), .A2(new_n728), .A3(new_n885), .A4(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n868), .A2(new_n770), .A3(new_n871), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n889), .A2(new_n765), .A3(new_n877), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n881), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n882), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n843), .B1(new_n879), .B2(new_n892), .ZN(new_n893));
  XOR2_X1   g707(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n894));
  OAI21_X1  g708(.A(KEYINPUT53), .B1(new_n863), .B2(new_n878), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n888), .A2(new_n891), .A3(new_n880), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n829), .A2(new_n825), .A3(new_n810), .ZN(new_n899));
  OR3_X1    g713(.A1(new_n834), .A2(KEYINPUT114), .A3(new_n335), .ZN(new_n900));
  OAI21_X1  g714(.A(KEYINPUT114), .B1(new_n834), .B2(new_n335), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n900), .B(new_n901), .C1(new_n793), .C2(new_n795), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n902), .A2(new_n836), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n833), .B1(new_n899), .B2(new_n903), .ZN(new_n904));
  NOR4_X1   g718(.A1(new_n822), .A2(new_n618), .A3(new_n636), .A4(new_n689), .ZN(new_n905));
  INV_X1    g719(.A(new_n615), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n811), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n907), .B(new_n908), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n909), .A2(KEYINPUT48), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(KEYINPUT48), .ZN(new_n911));
  AOI211_X1 g725(.A(new_n337), .B(new_n905), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n803), .A2(new_n746), .A3(new_n718), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n898), .A2(new_n904), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n799), .B1(new_n842), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n782), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n916), .A2(new_n614), .A3(new_n335), .A4(new_n449), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT108), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n919), .A2(new_n920), .A3(new_n689), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n711), .B(KEYINPUT49), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n921), .A2(new_n679), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n915), .A2(new_n923), .ZN(G75));
  NAND2_X1  g738(.A1(new_n895), .A2(new_n896), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n925), .A2(new_n321), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(G210), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT56), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n474), .A2(new_n484), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(new_n482), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT55), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n927), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n931), .B1(new_n927), .B2(new_n928), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n295), .A2(G952), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(G51));
  XOR2_X1   g749(.A(new_n323), .B(KEYINPUT57), .Z(new_n936));
  AND3_X1   g750(.A1(new_n895), .A2(new_n894), .A3(new_n896), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n936), .B1(new_n937), .B2(new_n897), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(KEYINPUT122), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n940), .B(new_n936), .C1(new_n937), .C2(new_n897), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n939), .A2(new_n319), .A3(new_n941), .ZN(new_n942));
  OR3_X1    g756(.A1(new_n925), .A2(new_n321), .A3(new_n774), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n934), .B1(new_n942), .B2(new_n943), .ZN(G54));
  NAND3_X1  g758(.A1(new_n926), .A2(KEYINPUT58), .A3(G475), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n945), .A2(new_n392), .A3(new_n381), .ZN(new_n946));
  INV_X1    g760(.A(new_n934), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n381), .A2(new_n392), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n926), .A2(KEYINPUT58), .A3(G475), .A4(new_n948), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(G60));
  AND2_X1   g764(.A1(new_n630), .A2(new_n632), .ZN(new_n951));
  NAND2_X1  g765(.A1(G478), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT59), .Z(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n951), .B(new_n954), .C1(new_n937), .C2(new_n897), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n898), .A2(new_n953), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n947), .B(new_n955), .C1(new_n956), .C2(new_n951), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(G63));
  NAND2_X1  g772(.A1(G217), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT60), .Z(new_n960));
  NAND3_X1  g774(.A1(new_n895), .A2(new_n896), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n600), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n888), .A2(new_n891), .A3(new_n880), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n880), .B1(new_n888), .B2(new_n891), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n966), .A2(KEYINPUT123), .A3(new_n656), .A4(new_n960), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n895), .A2(new_n896), .A3(new_n656), .A4(new_n960), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT123), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n934), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT124), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n967), .B2(new_n970), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n963), .B(new_n971), .C1(new_n973), .C2(KEYINPUT61), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n968), .A2(new_n969), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n968), .A2(new_n969), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n947), .B(new_n963), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n978));
  OAI21_X1  g792(.A(KEYINPUT124), .B1(new_n975), .B2(new_n976), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n974), .A2(new_n980), .ZN(G66));
  XNOR2_X1  g795(.A(new_n863), .B(KEYINPUT125), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n295), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT126), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n982), .A2(KEYINPUT126), .A3(new_n295), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(G953), .B1(new_n340), .B2(new_n480), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n929), .B1(G898), .B2(new_n295), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n990), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n987), .A2(new_n992), .A3(new_n988), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n991), .A2(new_n993), .ZN(G69));
  XNOR2_X1  g808(.A(new_n551), .B(new_n386), .ZN(new_n995));
  NAND2_X1  g809(.A1(G900), .A2(G953), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n787), .A2(new_n765), .ZN(new_n997));
  NOR4_X1   g811(.A1(new_n779), .A2(new_n625), .A3(new_n906), .A4(new_n680), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n874), .A2(new_n703), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n997), .A2(new_n797), .A3(new_n770), .A4(new_n1000), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n995), .B(new_n996), .C1(new_n1001), .C2(G953), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n855), .A2(new_n636), .ZN(new_n1003));
  NOR4_X1   g817(.A1(new_n674), .A2(new_n906), .A3(new_n813), .A4(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(new_n999), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n693), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT62), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1005), .A2(KEYINPUT62), .A3(new_n693), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1004), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n797), .A2(new_n1010), .A3(new_n787), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n1011), .A2(new_n295), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n995), .B(KEYINPUT127), .Z(new_n1013));
  OAI21_X1  g827(.A(new_n1002), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n295), .B1(G227), .B2(G900), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1015), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n1002), .B(new_n1017), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1016), .A2(new_n1018), .ZN(G72));
  NAND2_X1  g833(.A1(G472), .A2(G902), .ZN(new_n1020));
  XOR2_X1   g834(.A(new_n1020), .B(KEYINPUT63), .Z(new_n1021));
  OAI21_X1  g835(.A(new_n1021), .B1(new_n1001), .B2(new_n982), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1022), .A2(new_n558), .A3(new_n552), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1021), .B1(new_n1011), .B2(new_n982), .ZN(new_n1024));
  INV_X1    g838(.A(new_n682), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n879), .A2(new_n892), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n1027), .A2(new_n572), .A3(new_n682), .A4(new_n1021), .ZN(new_n1028));
  AND4_X1   g842(.A1(new_n947), .A2(new_n1023), .A3(new_n1026), .A4(new_n1028), .ZN(G57));
endmodule


