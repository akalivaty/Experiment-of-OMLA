//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999;
  OR2_X1    g000(.A1(KEYINPUT71), .A2(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT71), .A2(G953), .ZN(new_n188));
  AND2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(G210), .A3(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT27), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G101), .ZN(new_n193));
  XOR2_X1   g007(.A(new_n192), .B(new_n193), .Z(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G116), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G119), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT68), .B1(new_n198), .B2(G116), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT68), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(new_n196), .A3(G119), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n197), .B1(new_n199), .B2(new_n201), .ZN(new_n202));
  XOR2_X1   g016(.A(KEYINPUT2), .B(G113), .Z(new_n203));
  OR2_X1    g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n203), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT1), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n208), .A2(new_n210), .A3(new_n211), .A4(G128), .ZN(new_n212));
  AOI21_X1  g026(.A(G128), .B1(new_n208), .B2(new_n210), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n209), .A2(KEYINPUT1), .A3(G146), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT67), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT67), .ZN(new_n217));
  XNOR2_X1  g031(.A(G143), .B(G146), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n217), .B(new_n214), .C1(new_n218), .C2(G128), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT11), .ZN(new_n221));
  INV_X1    g035(.A(G134), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n221), .B1(new_n222), .B2(G137), .ZN(new_n223));
  INV_X1    g037(.A(G137), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(KEYINPUT11), .A3(G134), .ZN(new_n225));
  INV_X1    g039(.A(G131), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n222), .A2(G137), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n223), .A2(new_n225), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n222), .A2(G137), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n224), .A2(G134), .ZN(new_n230));
  OAI21_X1  g044(.A(G131), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n228), .A2(new_n231), .A3(KEYINPUT70), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n212), .A2(new_n220), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n223), .A2(new_n225), .A3(new_n227), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G131), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n240), .A3(new_n228), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(KEYINPUT66), .A3(G131), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n244));
  OAI211_X1 g058(.A(KEYINPUT0), .B(G128), .C1(new_n218), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n208), .A2(new_n210), .ZN(new_n246));
  NAND2_X1  g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(KEYINPUT65), .A3(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n249));
  NOR3_X1   g063(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(new_n208), .B2(new_n210), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n245), .A2(new_n248), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n237), .B1(new_n243), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n249), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n246), .A2(KEYINPUT65), .A3(new_n247), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n247), .B1(new_n246), .B2(KEYINPUT65), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n257), .A2(KEYINPUT69), .A3(new_n241), .A4(new_n242), .ZN(new_n258));
  AOI211_X1 g072(.A(new_n206), .B(new_n236), .C1(new_n253), .C2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n206), .ZN(new_n260));
  INV_X1    g074(.A(new_n212), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n261), .B1(new_n216), .B2(new_n219), .ZN(new_n262));
  OR2_X1    g076(.A1(new_n262), .A2(new_n232), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n257), .A2(new_n242), .A3(new_n241), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n260), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT28), .B1(new_n259), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n236), .A2(new_n206), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT28), .B1(new_n267), .B2(new_n264), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n195), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT30), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n263), .A2(new_n271), .A3(new_n264), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n236), .B1(new_n253), .B2(new_n258), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n272), .B1(new_n273), .B2(new_n271), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n206), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n259), .A2(new_n194), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT31), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT31), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n270), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(G472), .A2(G902), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT32), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n265), .B1(new_n273), .B2(new_n260), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT28), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n194), .B1(new_n287), .B2(new_n268), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n275), .A2(KEYINPUT31), .A3(new_n276), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT31), .B1(new_n275), .B2(new_n276), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT32), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n292), .A3(new_n282), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n273), .A2(new_n260), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n294), .B(KEYINPUT28), .C1(new_n295), .C2(new_n259), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n253), .A2(new_n258), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n206), .B1(new_n297), .B2(new_n236), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n273), .A2(new_n260), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n286), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n269), .A2(KEYINPUT72), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n296), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT29), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n194), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G902), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n269), .B(new_n195), .C1(new_n285), .C2(new_n286), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n259), .B1(new_n274), .B2(new_n206), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n307), .B(new_n303), .C1(new_n308), .C2(new_n195), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n305), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n284), .A2(new_n293), .B1(G472), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G217), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(G234), .B2(new_n306), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(G125), .B(G140), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT16), .ZN(new_n316));
  INV_X1    g130(.A(G125), .ZN(new_n317));
  OR3_X1    g131(.A1(new_n317), .A2(KEYINPUT16), .A3(G140), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n207), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n316), .A2(G146), .A3(new_n318), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G110), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n324), .B1(new_n198), .B2(G128), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n198), .A2(G128), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n324), .A2(new_n198), .A3(G128), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT24), .B(G110), .ZN(new_n330));
  OR3_X1    g144(.A1(new_n198), .A2(KEYINPUT73), .A3(G128), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT73), .B1(new_n198), .B2(G128), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n332), .A3(new_n326), .ZN(new_n333));
  OAI221_X1 g147(.A(new_n322), .B1(new_n323), .B2(new_n329), .C1(new_n330), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n315), .A2(new_n207), .ZN(new_n335));
  XOR2_X1   g149(.A(KEYINPUT74), .B(G110), .Z(new_n336));
  AND2_X1   g150(.A1(new_n329), .A2(new_n336), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n333), .A2(new_n330), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n321), .B(new_n335), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT22), .B(G137), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n334), .A2(new_n339), .A3(new_n343), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n306), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT25), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n345), .A2(KEYINPUT25), .A3(new_n306), .A4(new_n346), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n314), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n345), .A2(new_n346), .ZN(new_n352));
  NOR3_X1   g166(.A1(new_n352), .A2(G902), .A3(new_n313), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n311), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n187), .A2(G214), .A3(new_n190), .A4(new_n188), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n357), .A2(new_n209), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n209), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(KEYINPUT18), .A3(G131), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n315), .B(new_n207), .ZN(new_n362));
  NAND2_X1  g176(.A1(KEYINPUT18), .A2(G131), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n358), .A2(new_n359), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n361), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(G113), .B(G122), .ZN(new_n366));
  INV_X1    g180(.A(G104), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n366), .B(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(KEYINPUT90), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n226), .B1(new_n358), .B2(new_n359), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT17), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(new_n320), .A3(new_n321), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n358), .A2(new_n226), .A3(new_n359), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n374), .A2(new_n370), .A3(KEYINPUT17), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n365), .B(new_n369), .C1(new_n372), .C2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n365), .ZN(new_n377));
  INV_X1    g191(.A(new_n372), .ZN(new_n378));
  INV_X1    g192(.A(new_n375), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n376), .B1(new_n380), .B2(new_n368), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n306), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G475), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT20), .ZN(new_n384));
  NOR2_X1   g198(.A1(G475), .A2(G902), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT89), .B1(new_n374), .B2(new_n370), .ZN(new_n386));
  INV_X1    g200(.A(new_n370), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT89), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(new_n373), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n315), .B(KEYINPUT19), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n207), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n386), .A2(new_n389), .A3(new_n321), .A4(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n368), .B1(new_n392), .B2(new_n365), .ZN(new_n393));
  INV_X1    g207(.A(new_n376), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n384), .B(new_n385), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n391), .A2(new_n321), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n387), .A2(new_n373), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n397), .B1(new_n398), .B2(KEYINPUT89), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n377), .B1(new_n399), .B2(new_n389), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n376), .B1(new_n400), .B2(new_n368), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n384), .B1(new_n401), .B2(new_n385), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n383), .B1(new_n396), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G952), .ZN(new_n404));
  AOI211_X1 g218(.A(G953), .B(new_n404), .C1(G234), .C2(G237), .ZN(new_n405));
  AOI211_X1 g219(.A(new_n306), .B(new_n189), .C1(G234), .C2(G237), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT21), .B(G898), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT14), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT91), .ZN(new_n411));
  INV_X1    g225(.A(G122), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n411), .B1(new_n412), .B2(G116), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n196), .A2(KEYINPUT91), .A3(G122), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n410), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT95), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n196), .A2(G122), .ZN(new_n417));
  OR3_X1    g231(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n416), .B1(new_n415), .B2(new_n417), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n413), .A2(new_n410), .A3(new_n414), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G107), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n413), .A2(new_n414), .ZN(new_n423));
  INV_X1    g237(.A(G107), .ZN(new_n424));
  INV_X1    g238(.A(new_n417), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(KEYINPUT94), .ZN(new_n428));
  XNOR2_X1  g242(.A(G128), .B(G143), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(G134), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT94), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  NOR3_X1   g246(.A1(new_n428), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n422), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT9), .B(G234), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n435), .A2(new_n312), .A3(G953), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n429), .A2(KEYINPUT13), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n209), .A2(G128), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n437), .B(G134), .C1(KEYINPUT13), .C2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT93), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n439), .A2(new_n440), .B1(new_n222), .B2(new_n429), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT92), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n424), .B1(new_n423), .B2(new_n425), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n443), .B1(new_n427), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n444), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(KEYINPUT92), .A3(new_n426), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n441), .A2(new_n442), .A3(new_n445), .A4(new_n447), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n434), .A2(new_n436), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n436), .B1(new_n434), .B2(new_n448), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n306), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT96), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g267(.A(KEYINPUT96), .B(new_n306), .C1(new_n449), .C2(new_n450), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G478), .ZN(new_n456));
  OR2_X1    g270(.A1(new_n456), .A2(KEYINPUT15), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n434), .A2(new_n448), .ZN(new_n458));
  INV_X1    g272(.A(new_n436), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n434), .A2(new_n436), .A3(new_n448), .ZN(new_n461));
  AOI21_X1  g275(.A(G902), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT97), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n457), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n455), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n457), .B1(new_n451), .B2(new_n463), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n409), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n189), .A2(G227), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(KEYINPUT76), .ZN(new_n470));
  XNOR2_X1  g284(.A(G110), .B(G140), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n470), .B(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT77), .B(G104), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT3), .B1(new_n473), .B2(G107), .ZN(new_n474));
  AOI21_X1  g288(.A(G101), .B1(new_n473), .B2(G107), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT3), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(new_n424), .A3(G104), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n474), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n367), .A2(KEYINPUT77), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT77), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(G104), .ZN(new_n481));
  AOI21_X1  g295(.A(G107), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n424), .A2(G104), .ZN(new_n483));
  OAI21_X1  g297(.A(G101), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n262), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n212), .B(new_n214), .C1(G128), .C2(new_n218), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n478), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n243), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT12), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n489), .B(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT10), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n262), .A2(new_n492), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n478), .A2(new_n484), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n479), .A2(new_n481), .A3(G107), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n496), .B(new_n477), .C1(new_n482), .C2(new_n476), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G101), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(KEYINPUT4), .A3(new_n478), .ZN(new_n499));
  INV_X1    g313(.A(G101), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n499), .A2(new_n257), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT78), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n488), .A2(new_n504), .A3(new_n492), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n504), .B1(new_n488), .B2(new_n492), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n495), .B(new_n503), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n243), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n472), .B1(new_n491), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n508), .ZN(new_n511));
  INV_X1    g325(.A(new_n472), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n512), .B1(new_n507), .B2(new_n508), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n511), .B1(new_n513), .B2(KEYINPUT79), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT79), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n488), .A2(new_n492), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT78), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n488), .A2(new_n504), .A3(new_n492), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n519), .A2(new_n243), .A3(new_n495), .A4(new_n503), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n515), .B1(new_n520), .B2(new_n512), .ZN(new_n521));
  OAI211_X1 g335(.A(G469), .B(new_n510), .C1(new_n514), .C2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(G469), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n513), .A2(new_n491), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n512), .B1(new_n511), .B2(new_n520), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n523), .B(new_n306), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(G469), .A2(G902), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n522), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(G221), .B1(new_n435), .B2(G902), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(KEYINPUT75), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n468), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT88), .ZN(new_n533));
  OAI21_X1  g347(.A(G210), .B1(G237), .B2(G902), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(KEYINPUT86), .ZN(new_n535));
  NAND2_X1  g349(.A1(KEYINPUT84), .A2(KEYINPUT7), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n262), .A2(G125), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n252), .A2(new_n317), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G224), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT7), .B1(new_n540), .B2(G953), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n257), .A2(G125), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(G125), .B2(new_n262), .ZN(new_n544));
  INV_X1    g358(.A(new_n541), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n536), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n204), .A2(new_n205), .B1(new_n497), .B2(new_n501), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n499), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n202), .A2(KEYINPUT5), .ZN(new_n549));
  INV_X1    g363(.A(G113), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT5), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n550), .B1(new_n197), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n549), .A2(new_n552), .B1(new_n202), .B2(new_n203), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n494), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(G110), .B(G122), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n548), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n552), .B(KEYINPUT83), .ZN(new_n557));
  INV_X1    g371(.A(new_n549), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n205), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n494), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n555), .B(KEYINPUT8), .Z(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(new_n485), .B2(new_n553), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n542), .A2(new_n546), .A3(new_n556), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n306), .ZN(new_n565));
  INV_X1    g379(.A(new_n555), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT81), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(KEYINPUT82), .A3(KEYINPUT6), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n568), .B1(KEYINPUT82), .B2(KEYINPUT6), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT80), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n548), .A2(new_n554), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n570), .B1(new_n548), .B2(new_n554), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n566), .B(new_n569), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n548), .A2(new_n554), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT80), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n548), .A2(new_n554), .A3(new_n570), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n555), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n556), .A2(new_n567), .A3(KEYINPUT6), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n573), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n540), .A2(G953), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n544), .B(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n565), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT85), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n535), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n566), .B1(new_n571), .B2(new_n572), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n556), .A2(new_n567), .A3(KEYINPUT6), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n581), .B1(new_n588), .B2(new_n573), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n589), .A2(KEYINPUT85), .A3(new_n565), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT87), .B1(new_n585), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n583), .A2(new_n584), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT85), .B1(new_n589), .B2(new_n565), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT87), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n592), .A2(new_n593), .A3(new_n594), .A4(new_n535), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n535), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n583), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(G214), .B1(G237), .B2(G902), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n533), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI211_X1 g415(.A(new_n565), .B(new_n535), .C1(new_n579), .C2(new_n582), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(new_n591), .B2(new_n595), .ZN(new_n603));
  INV_X1    g417(.A(new_n600), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n603), .A2(KEYINPUT88), .A3(new_n604), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n356), .B(new_n532), .C1(new_n601), .C2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  INV_X1    g421(.A(new_n408), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n579), .A2(new_n582), .ZN(new_n609));
  INV_X1    g423(.A(new_n565), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n597), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n600), .B1(new_n611), .B2(new_n602), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT98), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(new_n459), .B2(KEYINPUT99), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n617), .B1(new_n449), .B2(new_n450), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n460), .A2(new_n461), .A3(new_n616), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n618), .A2(new_n619), .A3(G478), .A4(new_n306), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n614), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n393), .A2(new_n394), .ZN(new_n622));
  INV_X1    g436(.A(new_n385), .ZN(new_n623));
  OAI21_X1  g437(.A(KEYINPUT20), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n624), .A2(new_n395), .B1(G475), .B2(new_n382), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n535), .B1(new_n589), .B2(new_n565), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n598), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT98), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(new_n629), .A3(new_n600), .ZN(new_n630));
  AND4_X1   g444(.A1(new_n608), .A2(new_n613), .A3(new_n626), .A4(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n291), .A2(new_n306), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n633), .A2(G472), .B1(new_n282), .B2(new_n291), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n528), .A2(new_n530), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n634), .A2(new_n635), .A3(new_n354), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(new_n367), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  NOR2_X1   g454(.A1(new_n467), .A2(new_n403), .ZN(new_n641));
  AND4_X1   g455(.A1(new_n608), .A2(new_n613), .A3(new_n630), .A4(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n636), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT35), .B(G107), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  INV_X1    g460(.A(new_n634), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n344), .A2(KEYINPUT36), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n340), .B(new_n648), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n649), .A2(new_n306), .A3(new_n314), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n351), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n532), .B(new_n652), .C1(new_n601), .C2(new_n605), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  NOR3_X1   g469(.A1(new_n311), .A2(new_n531), .A3(new_n651), .ZN(new_n656));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n405), .B1(new_n406), .B2(new_n657), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n467), .A2(new_n403), .A3(new_n658), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n613), .A2(new_n630), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G128), .ZN(G30));
  XOR2_X1   g476(.A(new_n658), .B(KEYINPUT39), .Z(new_n663));
  NAND2_X1  g477(.A1(new_n635), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT103), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n603), .B(KEYINPUT38), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n467), .A2(new_n625), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n669), .A2(new_n600), .A3(new_n651), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n308), .A2(new_n194), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n298), .A2(new_n299), .A3(new_n194), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n306), .ZN(new_n674));
  OAI21_X1  g488(.A(G472), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT101), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI211_X1 g491(.A(KEYINPUT101), .B(G472), .C1(new_n672), .C2(new_n674), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n291), .A2(new_n292), .A3(new_n282), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n292), .B1(new_n291), .B2(new_n282), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n679), .B(KEYINPUT102), .C1(new_n680), .C2(new_n681), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n667), .A2(new_n671), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(new_n209), .ZN(G45));
  NAND2_X1  g503(.A1(new_n614), .A2(new_n620), .ZN(new_n690));
  INV_X1    g504(.A(new_n658), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n403), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n613), .A2(new_n630), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT105), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n613), .A2(new_n696), .A3(new_n630), .A4(new_n693), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n695), .A2(new_n656), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  NOR2_X1   g513(.A1(new_n524), .A2(new_n525), .ZN(new_n700));
  OAI21_X1  g514(.A(G469), .B1(new_n700), .B2(G902), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n530), .A3(new_n526), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n311), .A2(new_n355), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n631), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT41), .B(G113), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G15));
  NAND2_X1  g520(.A1(new_n642), .A2(new_n703), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G116), .ZN(G18));
  INV_X1    g522(.A(new_n702), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n613), .A2(new_n630), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n311), .A2(new_n651), .ZN(new_n711));
  INV_X1    g525(.A(new_n468), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT106), .B(G119), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G21));
  AND3_X1   g529(.A1(new_n613), .A2(new_n669), .A3(new_n630), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n302), .A2(new_n195), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n279), .A2(new_n280), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n283), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n701), .A2(new_n608), .A3(new_n530), .A4(new_n526), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT107), .B(G472), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n291), .B2(new_n306), .ZN(new_n723));
  NOR4_X1   g537(.A1(new_n719), .A2(new_n720), .A3(new_n723), .A4(new_n355), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n716), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  NOR4_X1   g540(.A1(new_n719), .A2(new_n692), .A3(new_n723), .A4(new_n651), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n710), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G125), .ZN(G27));
  AOI211_X1 g543(.A(new_n604), .B(new_n602), .C1(new_n591), .C2(new_n595), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n635), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n692), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(KEYINPUT108), .B1(new_n680), .B2(new_n681), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n310), .A2(G472), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n284), .A2(new_n737), .A3(new_n293), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n739), .A2(new_n740), .A3(new_n354), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n740), .B1(new_n739), .B2(new_n354), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n732), .B(new_n734), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n730), .A2(new_n356), .A3(new_n635), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n733), .B1(new_n745), .B2(new_n692), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n226), .ZN(G33));
  NAND4_X1  g563(.A1(new_n730), .A2(new_n356), .A3(new_n635), .A4(new_n659), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G134), .ZN(G36));
  NAND2_X1  g565(.A1(new_n603), .A2(new_n600), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n625), .A2(new_n690), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n753), .A2(KEYINPUT43), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(KEYINPUT43), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n756), .A2(new_n634), .A3(new_n651), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n752), .B1(new_n757), .B2(KEYINPUT44), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(KEYINPUT44), .B2(new_n757), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n510), .B1(new_n514), .B2(new_n521), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n523), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n760), .A2(new_n761), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n527), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n767), .A2(KEYINPUT111), .A3(KEYINPUT46), .A4(new_n527), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n766), .B1(new_n762), .B2(new_n763), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n762), .A2(new_n763), .ZN(new_n773));
  OAI211_X1 g587(.A(KEYINPUT46), .B(new_n527), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n770), .A2(new_n526), .A3(new_n771), .A4(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n530), .A3(new_n663), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n759), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(new_n224), .ZN(G39));
  NAND2_X1  g594(.A1(new_n777), .A2(new_n530), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n777), .A2(KEYINPUT47), .A3(new_n530), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n692), .A2(new_n354), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n785), .A2(new_n311), .A3(new_n730), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  NAND2_X1  g602(.A1(new_n701), .A2(new_n526), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n789), .A2(new_n530), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n783), .A2(new_n784), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n754), .A2(new_n405), .A3(new_n755), .ZN(new_n792));
  INV_X1    g606(.A(new_n719), .ZN(new_n793));
  INV_X1    g607(.A(new_n723), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(new_n354), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n730), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n791), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n668), .A2(new_n604), .A3(new_n709), .A4(new_n796), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT50), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n752), .A2(new_n702), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n354), .A2(new_n405), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n687), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT118), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n687), .A2(new_n803), .A3(new_n807), .A4(new_n804), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n806), .A2(new_n625), .A3(new_n621), .A4(new_n808), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n752), .A2(new_n792), .A3(new_n702), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n719), .A2(new_n651), .A3(new_n723), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT117), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n802), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT51), .B1(new_n799), .B2(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n802), .A2(new_n813), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n791), .A2(new_n798), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n816), .A2(new_n817), .A3(new_n818), .A4(new_n809), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n810), .B1(new_n741), .B2(new_n742), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT48), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n806), .A2(new_n626), .A3(new_n808), .ZN(new_n823));
  AOI211_X1 g637(.A(new_n404), .B(G953), .C1(new_n796), .C2(new_n710), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n820), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT119), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n820), .A2(new_n828), .A3(new_n825), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n351), .A2(new_n650), .A3(new_n658), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n528), .A2(new_n831), .A3(new_n530), .ZN(new_n832));
  AND4_X1   g646(.A1(new_n630), .A2(new_n613), .A3(new_n832), .A4(new_n669), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n686), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n698), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n661), .A2(new_n728), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT52), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n656), .A2(new_n660), .B1(new_n710), .B2(new_n727), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n838), .A2(new_n839), .A3(new_n698), .A4(new_n834), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT113), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n641), .A2(new_n626), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n636), .A2(new_n843), .A3(new_n408), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n844), .B1(new_n601), .B2(new_n605), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n606), .A2(new_n653), .A3(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n704), .A2(new_n707), .A3(new_n713), .A4(new_n725), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT112), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n613), .A2(new_n630), .A3(new_n709), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n850), .A2(new_n468), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n851), .A2(new_n711), .B1(new_n716), .B2(new_n724), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(KEYINPUT112), .A3(new_n704), .A4(new_n707), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n846), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n467), .A2(new_n625), .A3(new_n691), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n727), .B1(new_n711), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n750), .B1(new_n856), .B2(new_n731), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n857), .B1(new_n743), .B2(new_n746), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT113), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n837), .A2(new_n859), .A3(new_n840), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n842), .A2(new_n854), .A3(new_n858), .A4(new_n860), .ZN(new_n861));
  XNOR2_X1  g675(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n849), .A2(new_n853), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n606), .A2(new_n653), .A3(new_n845), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(new_n858), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n841), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(KEYINPUT53), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT54), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n847), .A2(KEYINPUT116), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n847), .A2(KEYINPUT116), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(KEYINPUT53), .A3(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n858), .ZN(new_n873));
  NOR4_X1   g687(.A1(new_n872), .A2(new_n873), .A3(new_n841), .A4(new_n846), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT115), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n861), .A2(new_n876), .A3(new_n862), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n876), .B1(new_n861), .B2(new_n862), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n869), .B1(new_n879), .B2(KEYINPUT54), .ZN(new_n880));
  OAI22_X1  g694(.A1(new_n830), .A2(new_n880), .B1(G952), .B2(G953), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n789), .A2(KEYINPUT49), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n789), .A2(KEYINPUT49), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n354), .A2(new_n600), .A3(new_n530), .ZN(new_n884));
  NOR4_X1   g698(.A1(new_n882), .A2(new_n883), .A3(new_n753), .A4(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n668), .A2(new_n687), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n881), .A2(new_n886), .ZN(G75));
  NAND3_X1  g701(.A1(new_n879), .A2(G902), .A3(new_n535), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n579), .B(new_n582), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT55), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n890), .A2(KEYINPUT56), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n189), .A2(G952), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT121), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n888), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n879), .A2(KEYINPUT120), .A3(G902), .A4(new_n535), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n895), .B1(new_n900), .B2(new_n890), .ZN(G51));
  XOR2_X1   g715(.A(new_n527), .B(KEYINPUT57), .Z(new_n902));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n837), .A2(new_n859), .A3(new_n840), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n859), .B1(new_n837), .B2(new_n840), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n866), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n862), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT115), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n861), .A2(new_n876), .A3(new_n862), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n903), .B1(new_n910), .B2(new_n875), .ZN(new_n911));
  AOI211_X1 g725(.A(KEYINPUT54), .B(new_n874), .C1(new_n908), .C2(new_n909), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n902), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n700), .B(KEYINPUT122), .Z(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n874), .B1(new_n908), .B2(new_n909), .ZN(new_n916));
  OR3_X1    g730(.A1(new_n916), .A2(new_n306), .A3(new_n767), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n893), .B1(new_n915), .B2(new_n917), .ZN(G54));
  NAND4_X1  g732(.A1(new_n879), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n919), .A2(new_n622), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(new_n622), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n920), .A2(new_n921), .A3(new_n893), .ZN(G60));
  AND2_X1   g736(.A1(new_n618), .A2(new_n619), .ZN(new_n923));
  NAND2_X1  g737(.A1(G478), .A2(G902), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT59), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n923), .B1(new_n880), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n923), .A2(new_n925), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n916), .A2(new_n903), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n879), .A2(KEYINPUT54), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n894), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n926), .A2(new_n930), .A3(new_n931), .ZN(G63));
  XNOR2_X1  g746(.A(new_n352), .B(KEYINPUT124), .ZN(new_n933));
  NAND2_X1  g747(.A1(G217), .A2(G902), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT60), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n933), .B1(new_n916), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n935), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n879), .A2(new_n649), .A3(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n936), .A2(new_n938), .A3(KEYINPUT61), .A4(new_n894), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n936), .A2(new_n894), .A3(new_n938), .ZN(new_n940));
  XNOR2_X1  g754(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(G66));
  INV_X1    g756(.A(new_n189), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n854), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT125), .ZN(new_n945));
  OAI21_X1  g759(.A(G953), .B1(new_n407), .B2(new_n540), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n588), .B(new_n573), .C1(G898), .C2(new_n189), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(G69));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n950));
  INV_X1    g764(.A(new_n779), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n665), .A2(new_n752), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n952), .B(new_n356), .C1(new_n626), .C2(new_n641), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n838), .A2(new_n698), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n688), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n688), .A2(new_n955), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n954), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n943), .B1(new_n961), .B2(new_n787), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n274), .B(new_n390), .Z(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n950), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n954), .ZN(new_n966));
  INV_X1    g780(.A(new_n960), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n966), .B(new_n787), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n189), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n970), .A2(KEYINPUT126), .A3(new_n963), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n963), .B1(G900), .B2(new_n943), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n716), .B1(new_n741), .B2(new_n742), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n778), .A2(new_n973), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n779), .A2(new_n974), .A3(new_n955), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n750), .B1(new_n744), .B2(new_n747), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n976), .A2(KEYINPUT127), .ZN(new_n977));
  INV_X1    g791(.A(new_n750), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n748), .A2(KEYINPUT127), .A3(new_n978), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n787), .B(new_n975), .C1(new_n977), .C2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n972), .B1(new_n980), .B2(new_n943), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n965), .A2(new_n971), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n983), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n965), .A2(new_n971), .A3(new_n981), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n984), .A2(new_n986), .ZN(G72));
  INV_X1    g801(.A(new_n672), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n961), .A2(new_n787), .A3(new_n854), .ZN(new_n989));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT63), .Z(new_n991));
  AOI21_X1  g805(.A(new_n988), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n863), .A2(new_n868), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n277), .B1(new_n195), .B2(new_n308), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n993), .A2(new_n991), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n308), .A2(new_n194), .ZN(new_n996));
  INV_X1    g810(.A(new_n854), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n980), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n996), .B1(new_n998), .B2(new_n991), .ZN(new_n999));
  NOR4_X1   g813(.A1(new_n992), .A2(new_n995), .A3(new_n999), .A4(new_n893), .ZN(G57));
endmodule


