//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n207));
  INV_X1    g0007(.A(G226), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n207), .B1(new_n202), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n206), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT1), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n206), .A2(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(KEYINPUT0), .ZN(new_n219));
  INV_X1    g0019(.A(new_n201), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G50), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(new_n218), .A2(new_n219), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n226), .B1(new_n219), .B2(new_n218), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n216), .A2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  INV_X1    g0036(.A(G107), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n237), .A2(G97), .ZN(new_n238));
  INV_X1    g0038(.A(G97), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n239), .A2(G107), .ZN(new_n240));
  AND2_X1   g0040(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  NOR2_X1   g0047(.A1(KEYINPUT64), .A2(G41), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT64), .A2(G41), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G45), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  AND2_X1   g0054(.A1(new_n254), .A2(G274), .ZN(new_n255));
  AND2_X1   g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  AOI21_X1  g0058(.A(G1), .B1(new_n258), .B2(new_n252), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n260), .A2(G244), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G33), .ZN(new_n265));
  AND3_X1   g0065(.A1(new_n263), .A2(new_n265), .A3(G1698), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n263), .A2(new_n265), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n266), .A2(G238), .B1(G107), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G232), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n268), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  AOI211_X1 g0073(.A(new_n256), .B(new_n261), .C1(new_n273), .C2(new_n257), .ZN(new_n274));
  INV_X1    g0074(.A(G179), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n274), .A2(G169), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n254), .A2(G13), .A3(G20), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G77), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n223), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n284), .B1(G1), .B2(new_n224), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n281), .B1(new_n285), .B2(new_n280), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT66), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n287), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(new_n288), .B2(new_n290), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n224), .A2(G33), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT15), .B(G87), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n292), .B1(new_n224), .B2(new_n280), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n286), .B1(new_n295), .B2(new_n283), .ZN(new_n296));
  OR3_X1    g0096(.A1(new_n276), .A2(new_n277), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n274), .A2(G190), .ZN(new_n298));
  INV_X1    g0098(.A(G200), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n298), .B(new_n296), .C1(new_n299), .C2(new_n274), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g0101(.A(new_n301), .B(KEYINPUT67), .Z(new_n302));
  AOI21_X1  g0102(.A(new_n256), .B1(G238), .B2(new_n260), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n266), .A2(G232), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G97), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n304), .B(new_n305), .C1(new_n208), .C2(new_n272), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n257), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(KEYINPUT13), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT13), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n310), .B1(new_n303), .B2(new_n307), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G190), .ZN(new_n313));
  INV_X1    g0113(.A(G68), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G20), .ZN(new_n315));
  OAI221_X1 g0115(.A(new_n315), .B1(new_n293), .B2(new_n280), .C1(new_n290), .C2(new_n202), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n283), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT69), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT11), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n317), .A2(KEYINPUT69), .ZN(new_n322));
  OR3_X1    g0122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n321), .B1(new_n320), .B2(new_n322), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n278), .A2(G68), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT12), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n285), .A2(new_n314), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n323), .A2(new_n324), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(G200), .B1(new_n309), .B2(new_n311), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n313), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(G169), .B1(new_n309), .B2(new_n311), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT14), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT14), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n335), .B(G169), .C1(new_n309), .C2(new_n311), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n312), .A2(G179), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n334), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n332), .B1(new_n338), .B2(new_n329), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n270), .A2(G226), .A3(G1698), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n270), .A2(G223), .A3(new_n271), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n341), .B(new_n342), .C1(new_n262), .C2(new_n209), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n257), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n253), .A2(new_n255), .B1(new_n260), .B2(G232), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n299), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n344), .A2(new_n345), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n346), .B1(G190), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G58), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n349), .A2(new_n314), .ZN(new_n350));
  OAI21_X1  g0150(.A(G20), .B1(new_n350), .B2(new_n201), .ZN(new_n351));
  INV_X1    g0151(.A(G159), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n351), .B1(new_n352), .B2(new_n290), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT7), .B1(new_n267), .B2(new_n224), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n314), .B1(new_n354), .B2(KEYINPUT70), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT7), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n270), .B2(G20), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n267), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT70), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n353), .B1(new_n355), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n284), .B1(new_n361), .B2(KEYINPUT16), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT16), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n314), .B1(new_n357), .B2(new_n358), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n363), .B1(new_n364), .B2(new_n353), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n287), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n367), .A2(new_n279), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n285), .B2(new_n367), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n348), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT17), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n369), .B1(new_n362), .B2(new_n365), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT17), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n374), .A3(new_n348), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n366), .A2(new_n370), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n344), .A2(G179), .A3(new_n345), .ZN(new_n378));
  INV_X1    g0178(.A(G169), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n344), .B2(new_n345), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT18), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n377), .A2(new_n381), .A3(KEYINPUT18), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n376), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n266), .A2(G223), .B1(G77), .B2(new_n267), .ZN(new_n386));
  INV_X1    g0186(.A(G222), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(new_n272), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n257), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n256), .B1(G226), .B2(new_n260), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G190), .ZN(new_n392));
  MUX2_X1   g0192(.A(new_n278), .B(new_n285), .S(G50), .Z(new_n393));
  NAND2_X1  g0193(.A1(new_n203), .A2(G20), .ZN(new_n394));
  INV_X1    g0194(.A(G150), .ZN(new_n395));
  OAI221_X1 g0195(.A(new_n394), .B1(new_n395), .B2(new_n290), .C1(new_n287), .C2(new_n293), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n283), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT9), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n398), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT9), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n392), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n391), .A2(new_n299), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n392), .A2(KEYINPUT68), .A3(new_n400), .A4(new_n402), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT10), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n406), .B(new_n407), .C1(new_n403), .C2(new_n404), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n391), .A2(KEYINPUT65), .A3(new_n275), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT65), .ZN(new_n412));
  INV_X1    g0212(.A(new_n391), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n412), .B1(new_n413), .B2(G179), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n401), .B1(new_n413), .B2(new_n379), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n411), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n409), .A2(new_n410), .A3(new_n416), .ZN(new_n417));
  NOR4_X1   g0217(.A1(new_n302), .A2(new_n340), .A3(new_n385), .A4(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n263), .A2(new_n265), .A3(G250), .A4(new_n271), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n263), .A2(new_n265), .A3(G257), .A4(G1698), .ZN(new_n420));
  INV_X1    g0220(.A(G294), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n419), .B(new_n420), .C1(new_n262), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n257), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT5), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n249), .A2(new_n424), .A3(new_n250), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n254), .B(G45), .C1(new_n424), .C2(G41), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(new_n427), .A3(G274), .ZN(new_n428));
  INV_X1    g0228(.A(new_n257), .ZN(new_n429));
  INV_X1    g0229(.A(new_n250), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n430), .A2(new_n248), .A3(KEYINPUT5), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n429), .B(G264), .C1(new_n431), .C2(new_n426), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n423), .A2(new_n428), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(G200), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n423), .A2(G190), .A3(new_n428), .A4(new_n432), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n279), .A2(KEYINPUT25), .A3(new_n237), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT25), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n278), .B2(G107), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(KEYINPUT81), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT81), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(new_n438), .C1(new_n278), .C2(G107), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n254), .A2(G33), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n284), .A2(KEYINPUT72), .A3(new_n278), .A4(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n278), .A2(new_n444), .A3(new_n223), .A4(new_n282), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT72), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n237), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n443), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT23), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n224), .B2(G107), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n237), .A2(KEYINPUT23), .A3(G20), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G116), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n262), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n224), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n263), .A2(new_n265), .A3(new_n224), .A4(G87), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT22), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT22), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n270), .A2(new_n461), .A3(new_n224), .A4(G87), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n458), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n283), .B1(new_n463), .B2(KEYINPUT24), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n460), .A2(new_n462), .ZN(new_n465));
  INV_X1    g0265(.A(new_n458), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n465), .A2(KEYINPUT24), .A3(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n450), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n436), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n422), .A2(new_n257), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n432), .A2(new_n428), .ZN(new_n471));
  OAI21_X1  g0271(.A(G169), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n423), .A2(G179), .A3(new_n428), .A4(new_n432), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n465), .A2(new_n466), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT24), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n463), .A2(KEYINPUT24), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n477), .A2(new_n283), .A3(new_n478), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n474), .A2(KEYINPUT82), .B1(new_n479), .B2(new_n450), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT82), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n472), .A2(new_n481), .A3(new_n473), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n469), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT71), .ZN(new_n484));
  NOR4_X1   g0284(.A1(new_n484), .A2(new_n280), .A3(G20), .A4(G33), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT71), .B1(new_n289), .B2(G77), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT6), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n238), .A2(new_n240), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n237), .A2(KEYINPUT6), .A3(G97), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n487), .B1(new_n491), .B2(new_n224), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n237), .B1(new_n357), .B2(new_n358), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n283), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n278), .A2(G97), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n445), .A2(new_n448), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(G97), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n263), .A2(new_n265), .A3(G250), .A4(G1698), .ZN(new_n499));
  NOR2_X1   g0299(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n500), .B1(G33), .B2(G283), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n263), .A2(new_n265), .A3(G244), .A4(new_n271), .ZN(new_n502));
  NAND2_X1  g0302(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n499), .B(new_n501), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n502), .A2(new_n503), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n257), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n257), .B1(new_n425), .B2(new_n427), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G257), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(new_n428), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n498), .B1(G200), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n506), .A2(new_n508), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n511), .A2(G190), .A3(new_n428), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(new_n275), .A3(new_n428), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n509), .A2(new_n379), .B1(new_n494), .B2(new_n497), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n510), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT76), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n496), .A2(G87), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT19), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n224), .B1(new_n305), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n209), .A2(new_n239), .A3(new_n237), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n263), .A2(new_n265), .A3(new_n224), .A4(G68), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n518), .B1(new_n293), .B2(new_n239), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n283), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n294), .A2(new_n279), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n525), .A2(KEYINPUT75), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT75), .B1(new_n525), .B2(new_n526), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n517), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n270), .A2(G244), .A3(G1698), .ZN(new_n530));
  INV_X1    g0330(.A(new_n456), .ZN(new_n531));
  INV_X1    g0331(.A(G238), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n530), .B(new_n531), .C1(new_n272), .C2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n257), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n254), .A2(G45), .A3(G274), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT74), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OR2_X1    g0337(.A1(new_n535), .A2(new_n536), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n210), .B1(new_n254), .B2(G45), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n537), .A2(new_n538), .B1(new_n429), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n299), .B1(new_n534), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n516), .B1(new_n529), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n528), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n525), .A2(KEYINPUT75), .A3(new_n526), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n534), .A2(new_n540), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G200), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n545), .A2(KEYINPUT76), .A3(new_n547), .A4(new_n517), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n534), .A2(new_n540), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G190), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n542), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n546), .A2(G179), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(new_n379), .B2(new_n546), .ZN(new_n553));
  INV_X1    g0353(.A(new_n496), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n545), .B1(new_n294), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n483), .A2(new_n515), .A3(new_n551), .A4(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT21), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n507), .A2(G270), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n428), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n263), .A2(new_n265), .A3(G257), .A4(new_n271), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT77), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT77), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n270), .A2(new_n563), .A3(G257), .A4(new_n271), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n264), .A2(G33), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n567));
  OAI21_X1  g0367(.A(G303), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n263), .A2(new_n265), .A3(G264), .A4(G1698), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n429), .B1(new_n571), .B2(KEYINPUT78), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n568), .A2(new_n569), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n562), .B2(new_n564), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT78), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n560), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n282), .A2(new_n223), .B1(G20), .B2(new_n455), .ZN(new_n578));
  AOI21_X1  g0378(.A(G20), .B1(G33), .B2(G283), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(G33), .B2(new_n239), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT20), .ZN(new_n582));
  OAI21_X1  g0382(.A(KEYINPUT79), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n582), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT79), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n578), .A2(new_n580), .A3(new_n585), .A4(KEYINPUT20), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  MUX2_X1   g0387(.A(new_n278), .B(new_n446), .S(G116), .Z(new_n588));
  AOI21_X1  g0388(.A(new_n379), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n558), .B1(new_n577), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n560), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n257), .B1(new_n574), .B2(new_n575), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n571), .A2(KEYINPUT78), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(KEYINPUT21), .A3(new_n589), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n587), .A2(new_n588), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n577), .A2(G179), .A3(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n591), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT80), .ZN(new_n600));
  OAI211_X1 g0400(.A(G190), .B(new_n592), .C1(new_n593), .C2(new_n594), .ZN(new_n601));
  INV_X1    g0401(.A(new_n597), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n601), .B(new_n602), .C1(new_n577), .C2(new_n299), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n599), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n603), .A2(new_n598), .A3(new_n596), .A4(new_n591), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT80), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n557), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n418), .A2(new_n607), .ZN(G372));
  NAND2_X1  g0408(.A1(new_n551), .A2(new_n556), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n514), .A2(new_n513), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT26), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OR2_X1    g0411(.A1(new_n436), .A2(new_n468), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n509), .A2(G200), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n512), .A2(new_n494), .A3(new_n497), .A4(new_n613), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n612), .A2(new_n614), .A3(new_n610), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n545), .A2(new_n547), .A3(new_n517), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT83), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n529), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n619), .A2(KEYINPUT83), .A3(new_n547), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n620), .A3(new_n550), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n474), .A2(new_n468), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n591), .A2(new_n596), .A3(new_n598), .A4(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n615), .A2(new_n556), .A3(new_n621), .A4(new_n623), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n556), .B(KEYINPUT84), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT26), .ZN(new_n626));
  INV_X1    g0426(.A(new_n610), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n621), .A2(new_n626), .A3(new_n556), .A4(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n611), .A2(new_n624), .A3(new_n625), .A4(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n418), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n384), .A2(new_n382), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n338), .A2(new_n329), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n297), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n372), .A2(new_n375), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(new_n332), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n631), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n409), .A2(new_n410), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n416), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n630), .A2(new_n638), .ZN(G369));
  XOR2_X1   g0439(.A(KEYINPUT85), .B(KEYINPUT27), .Z(new_n640));
  INV_X1    g0440(.A(G13), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n641), .A2(G1), .A3(G20), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n640), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G213), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(G343), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n602), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n600), .B1(new_n599), .B2(new_n603), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n605), .A2(KEYINPUT80), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n599), .A2(new_n650), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n468), .A2(new_n647), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n483), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n474), .A2(KEYINPUT82), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n659), .A2(new_n482), .A3(new_n468), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n658), .B1(new_n660), .B2(new_n648), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n656), .A2(KEYINPUT86), .A3(G330), .A4(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n649), .B1(new_n604), .B2(new_n606), .ZN(new_n663));
  OAI211_X1 g0463(.A(G330), .B(new_n661), .C1(new_n663), .C2(new_n654), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT86), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n591), .A2(new_n596), .A3(new_n598), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n483), .A2(new_n668), .A3(new_n648), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n474), .A2(new_n468), .A3(new_n648), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n669), .A2(KEYINPUT87), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(KEYINPUT87), .B1(new_n669), .B2(new_n670), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n667), .A2(new_n673), .ZN(G399));
  INV_X1    g0474(.A(new_n251), .ZN(new_n675));
  INV_X1    g0475(.A(new_n217), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n520), .A2(G116), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G1), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n221), .B2(new_n678), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT28), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n660), .A2(new_n610), .A3(new_n612), .A4(new_n614), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n609), .A2(new_n683), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n684), .B(new_n648), .C1(new_n651), .C2(new_n652), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT30), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n577), .A2(G179), .ZN(new_n687));
  INV_X1    g0487(.A(new_n433), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n511), .A2(new_n549), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n686), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n511), .A2(new_n549), .A3(new_n688), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n691), .A2(KEYINPUT30), .A3(G179), .A4(new_n577), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n549), .A2(new_n688), .A3(G179), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(new_n595), .A3(new_n509), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n690), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n647), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n696), .A2(KEYINPUT31), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n685), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n696), .A2(KEYINPUT31), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n698), .A2(G330), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT88), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n699), .B1(new_n685), .B2(new_n697), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT88), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(new_n704), .A3(G330), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n629), .A2(new_n648), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n621), .A2(new_n556), .A3(new_n627), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT26), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n660), .A2(new_n598), .A3(new_n596), .A4(new_n591), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n615), .A2(new_n710), .A3(new_n556), .A4(new_n621), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n551), .A2(new_n626), .A3(new_n556), .A4(new_n627), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n709), .A2(new_n711), .A3(new_n625), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n648), .ZN(new_n714));
  MUX2_X1   g0514(.A(new_n707), .B(new_n714), .S(KEYINPUT29), .Z(new_n715));
  NOR2_X1   g0515(.A1(new_n706), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n682), .B1(new_n716), .B2(G1), .ZN(G364));
  INV_X1    g0517(.A(new_n656), .ZN(new_n718));
  INV_X1    g0518(.A(G330), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n641), .A2(G20), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n254), .B1(new_n721), .B2(G45), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n678), .A2(KEYINPUT89), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT89), .ZN(new_n724));
  INV_X1    g0524(.A(new_n722), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n724), .B1(new_n677), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n720), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(G330), .B2(new_n656), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n224), .A2(G190), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n731), .A2(new_n275), .A3(G200), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT91), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G107), .ZN(new_n738));
  INV_X1    g0538(.A(G190), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n224), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n275), .A2(new_n299), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n275), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n743), .A2(new_n202), .B1(new_n745), .B2(new_n349), .ZN(new_n746));
  NOR4_X1   g0546(.A1(new_n224), .A2(new_n739), .A3(new_n299), .A4(G179), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n741), .A2(new_n731), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n748), .A2(new_n209), .B1(new_n749), .B2(new_n314), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G179), .A2(G200), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n224), .B1(new_n752), .B2(G190), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n239), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n744), .A2(new_n731), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n267), .B(new_n754), .C1(G77), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n731), .A2(new_n752), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n352), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT32), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n738), .A2(new_n751), .A3(new_n756), .A4(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n757), .ZN(new_n761));
  AOI22_X1  g0561(.A1(G329), .A2(new_n761), .B1(new_n755), .B2(G311), .ZN(new_n762));
  XOR2_X1   g0562(.A(KEYINPUT33), .B(G317), .Z(new_n763));
  OAI21_X1  g0563(.A(new_n762), .B1(new_n749), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n745), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n270), .B(new_n764), .C1(G322), .C2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G283), .ZN(new_n767));
  INV_X1    g0567(.A(G303), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n748), .A2(KEYINPUT94), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n748), .A2(KEYINPUT94), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n766), .B1(new_n767), .B2(new_n736), .C1(new_n768), .C2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(KEYINPUT92), .B(G326), .ZN(new_n773));
  INV_X1    g0573(.A(new_n753), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n742), .A2(new_n773), .B1(new_n774), .B2(G294), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT93), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n760), .B1(new_n772), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n223), .B1(G20), .B2(new_n379), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n676), .A2(new_n267), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT90), .Z(new_n781));
  AOI22_X1  g0581(.A1(new_n781), .A2(G355), .B1(new_n455), .B2(new_n676), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n246), .A2(new_n252), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n676), .A2(new_n270), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(G45), .B2(new_n221), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n782), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G13), .A2(G33), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(G20), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n778), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n727), .B1(new_n786), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n789), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n779), .B(new_n791), .C1(new_n656), .C2(new_n792), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n730), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(G396));
  INV_X1    g0595(.A(new_n706), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n297), .A2(new_n647), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n300), .B1(new_n296), .B2(new_n648), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n797), .B1(new_n297), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n707), .B(new_n799), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n801), .A2(KEYINPUT96), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(KEYINPUT96), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n796), .A2(new_n800), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n802), .A2(new_n727), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n778), .A2(new_n787), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n728), .B1(G77), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n771), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G107), .ZN(new_n810));
  INV_X1    g0610(.A(new_n755), .ZN(new_n811));
  INV_X1    g0611(.A(G311), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n811), .A2(new_n455), .B1(new_n757), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(KEYINPUT95), .B(G283), .Z(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n815), .A2(new_n749), .B1(new_n421), .B2(new_n745), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n270), .B(new_n754), .C1(G303), .C2(new_n742), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n737), .A2(G87), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n810), .A2(new_n817), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n742), .A2(G137), .B1(new_n755), .B2(G159), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n765), .A2(G143), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n821), .B(new_n822), .C1(new_n395), .C2(new_n749), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT34), .Z(new_n824));
  INV_X1    g0624(.A(G132), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n270), .B1(new_n757), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(G58), .B2(new_n774), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n827), .B1(new_n314), .B2(new_n736), .C1(new_n771), .C2(new_n202), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n820), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n808), .B1(new_n829), .B2(new_n778), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n799), .B2(new_n788), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n805), .A2(new_n831), .ZN(G384));
  INV_X1    g0632(.A(new_n491), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n833), .A2(KEYINPUT35), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n834), .A2(G116), .A3(new_n225), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(KEYINPUT35), .B2(new_n833), .ZN(new_n836));
  XOR2_X1   g0636(.A(KEYINPUT97), .B(KEYINPUT36), .Z(new_n837));
  OAI21_X1  g0637(.A(G77), .B1(new_n349), .B2(new_n314), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n221), .A2(new_n838), .B1(G50), .B2(new_n314), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n254), .A2(G13), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n836), .A2(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n696), .A2(KEYINPUT31), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n607), .B2(new_n648), .ZN(new_n843));
  OAI21_X1  g0643(.A(KEYINPUT100), .B1(new_n843), .B2(new_n699), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT100), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n698), .A2(new_n845), .A3(new_n700), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT99), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n632), .B2(new_n648), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n333), .A2(KEYINPUT14), .B1(new_n312), .B2(G179), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n330), .B1(new_n849), .B2(new_n336), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n850), .A2(KEYINPUT99), .A3(new_n647), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n329), .A2(new_n647), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n339), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n844), .A2(new_n846), .A3(new_n799), .A4(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n645), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n377), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n377), .A2(new_n381), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n860), .A2(new_n858), .A3(new_n371), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT37), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n860), .A2(new_n858), .A3(new_n863), .A4(new_n371), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n385), .A2(new_n859), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n865), .A2(KEYINPUT38), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n378), .A2(new_n380), .A3(new_n857), .ZN(new_n867));
  OR2_X1    g0667(.A1(new_n361), .A2(KEYINPUT16), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n369), .B1(new_n868), .B2(new_n362), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n371), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n864), .ZN(new_n872));
  INV_X1    g0672(.A(new_n382), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n873), .A2(new_n383), .B1(new_n372), .B2(new_n375), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n869), .A2(new_n645), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n872), .B(KEYINPUT38), .C1(new_n874), .C2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n866), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT40), .B1(new_n856), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n845), .B1(new_n698), .B2(new_n700), .ZN(new_n881));
  AOI211_X1 g0681(.A(KEYINPUT100), .B(new_n699), .C1(new_n685), .C2(new_n697), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n385), .A2(new_n875), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT38), .B1(new_n884), .B2(new_n872), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT40), .B1(new_n886), .B2(new_n877), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n883), .A2(new_n799), .A3(new_n855), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n880), .A2(new_n888), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n883), .A2(new_n418), .ZN(new_n890));
  OAI21_X1  g0690(.A(G330), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n892), .A2(KEYINPUT101), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n892), .A2(KEYINPUT101), .ZN(new_n894));
  AOI211_X1 g0694(.A(new_n893), .B(new_n894), .C1(new_n889), .C2(new_n890), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT39), .B1(new_n878), .B2(new_n885), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n877), .B(new_n897), .C1(new_n865), .C2(KEYINPUT38), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n632), .A2(new_n647), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n629), .A2(new_n799), .A3(new_n648), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n797), .B(KEYINPUT98), .Z(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n904), .B(new_n855), .C1(new_n878), .C2(new_n885), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n631), .A2(new_n645), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n901), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n638), .B1(new_n715), .B2(new_n418), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n907), .B(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n895), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n254), .B2(new_n721), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n895), .A2(new_n909), .ZN(new_n912));
  OAI221_X1 g0712(.A(new_n841), .B1(new_n836), .B2(new_n837), .C1(new_n911), .C2(new_n912), .ZN(G367));
  NAND2_X1  g0713(.A1(new_n529), .A2(new_n647), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n625), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n621), .A2(new_n556), .A3(new_n914), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n915), .B1(KEYINPUT102), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(KEYINPUT102), .B2(new_n916), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n918), .A2(new_n792), .ZN(new_n919));
  INV_X1    g0719(.A(new_n784), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n235), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n790), .B1(new_n217), .B2(new_n294), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n728), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI22_X1  g0723(.A1(G107), .A2(new_n774), .B1(new_n755), .B2(new_n814), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n924), .A2(KEYINPUT106), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT46), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n771), .A2(new_n926), .A3(new_n455), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n925), .B1(new_n928), .B2(KEYINPUT107), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n737), .A2(G97), .ZN(new_n930));
  INV_X1    g0730(.A(G317), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n745), .A2(new_n768), .B1(new_n757), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n926), .B1(new_n748), .B2(new_n455), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n933), .B(new_n267), .C1(new_n421), .C2(new_n749), .ZN(new_n934));
  AOI211_X1 g0734(.A(new_n932), .B(new_n934), .C1(G311), .C2(new_n742), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT107), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n927), .A2(new_n936), .B1(KEYINPUT106), .B2(new_n924), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n929), .A2(new_n930), .A3(new_n935), .A4(new_n937), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n765), .A2(G150), .B1(new_n742), .B2(G143), .ZN(new_n939));
  INV_X1    g0739(.A(G137), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n939), .B1(new_n940), .B2(new_n757), .C1(new_n352), .C2(new_n749), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n753), .A2(new_n314), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n748), .A2(new_n349), .B1(new_n811), .B2(new_n202), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n270), .B1(new_n736), .B2(new_n280), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n944), .B1(KEYINPUT108), .B2(new_n945), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n945), .A2(KEYINPUT108), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n938), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT47), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n778), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n948), .B2(new_n949), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n923), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n919), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n498), .A2(new_n647), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n515), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n627), .A2(new_n647), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  XOR2_X1   g0758(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n959));
  OAI211_X1 g0759(.A(new_n958), .B(new_n959), .C1(new_n671), .C2(new_n672), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n958), .B1(new_n671), .B2(new_n672), .ZN(new_n961));
  INV_X1    g0761(.A(new_n959), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n958), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT44), .B1(new_n673), .B2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT44), .ZN(new_n966));
  NOR4_X1   g0766(.A1(new_n671), .A2(new_n672), .A3(new_n966), .A4(new_n958), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n960), .B(new_n963), .C1(new_n965), .C2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT105), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n968), .A2(new_n667), .A3(new_n969), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n671), .A2(new_n672), .A3(new_n958), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT44), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n662), .A2(new_n666), .A3(new_n969), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n963), .A2(new_n960), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n970), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n599), .A2(new_n647), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n669), .B1(new_n661), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n720), .B(new_n978), .Z(new_n979));
  OAI21_X1  g0779(.A(new_n716), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n677), .B(KEYINPUT41), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n725), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n977), .A2(new_n515), .A3(new_n483), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n983), .A2(KEYINPUT42), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n610), .B1(new_n956), .B2(new_n660), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n983), .A2(KEYINPUT42), .B1(new_n986), .B2(new_n648), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n918), .A2(KEYINPUT43), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n662), .A2(new_n666), .A3(new_n958), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(KEYINPUT103), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT103), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n662), .A2(new_n666), .A3(new_n993), .A4(new_n958), .ZN(new_n994));
  AND3_X1   g0794(.A1(new_n991), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n992), .B1(new_n991), .B2(new_n994), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n989), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n991), .A2(new_n994), .ZN(new_n998));
  INV_X1    g0798(.A(new_n992), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n991), .A2(new_n992), .A3(new_n994), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1000), .A2(new_n988), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n954), .B1(new_n982), .B2(new_n1003), .ZN(G387));
  OAI21_X1  g0804(.A(new_n784), .B1(new_n232), .B2(new_n252), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n781), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1005), .B1(new_n679), .B2(new_n1006), .ZN(new_n1007));
  OR3_X1    g0807(.A1(new_n287), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1008));
  OAI21_X1  g0808(.A(KEYINPUT50), .B1(new_n287), .B2(G50), .ZN(new_n1009));
  AOI21_X1  g0809(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1008), .A2(new_n679), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n1007), .A2(new_n1011), .B1(new_n237), .B2(new_n676), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n790), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n728), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n743), .A2(new_n352), .B1(new_n748), .B2(new_n280), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n267), .B(new_n1015), .C1(G68), .C2(new_n755), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n753), .A2(new_n294), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n202), .A2(new_n745), .B1(new_n749), .B2(new_n287), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G150), .B2(new_n761), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1016), .A2(new_n930), .A3(new_n1017), .A4(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n270), .B1(new_n761), .B2(new_n773), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G294), .A2(new_n747), .B1(new_n774), .B2(new_n814), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n742), .A2(G322), .B1(new_n755), .B2(G303), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n812), .B2(new_n749), .C1(new_n931), .C2(new_n745), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT48), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1022), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT109), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n1025), .B2(new_n1024), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1021), .B1(new_n455), .B2(new_n736), .C1(new_n1028), .C2(KEYINPUT49), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1028), .A2(KEYINPUT49), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1020), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1014), .B1(new_n1031), .B2(new_n778), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n661), .B2(new_n792), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1033), .A2(KEYINPUT110), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(KEYINPUT110), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n720), .B(new_n978), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n1034), .A2(new_n1035), .B1(new_n725), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n716), .A2(new_n1036), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n677), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n716), .A2(new_n1036), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1037), .B1(new_n1039), .B2(new_n1040), .ZN(G393));
  OR2_X1    g0841(.A1(new_n968), .A2(new_n667), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n968), .A2(new_n667), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n1038), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n716), .A2(new_n1036), .A3(new_n970), .A4(new_n975), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1045), .A2(new_n677), .A3(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1042), .A2(new_n725), .A3(new_n1043), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n243), .A2(new_n920), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n790), .B1(new_n239), .B2(new_n217), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n728), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n267), .B1(new_n748), .B2(new_n815), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G322), .A2(new_n761), .B1(new_n755), .B2(G294), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n768), .B2(new_n749), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1052), .B(new_n1054), .C1(G116), .C2(new_n774), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n743), .A2(new_n931), .B1(new_n745), .B2(new_n812), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT52), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1055), .A2(new_n738), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n267), .B1(new_n761), .B2(G143), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n819), .B(new_n1061), .C1(new_n314), .C2(new_n748), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT112), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n743), .A2(new_n395), .B1(new_n745), .B2(new_n352), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n811), .A2(new_n287), .B1(new_n202), .B2(new_n749), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(G77), .B2(new_n774), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1066), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1060), .B1(new_n1063), .B2(new_n1070), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1071), .A2(KEYINPUT113), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n951), .B1(new_n1071), .B2(KEYINPUT113), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1051), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n792), .B2(new_n958), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1048), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1047), .A2(new_n1076), .ZN(G390));
  NAND3_X1  g0877(.A1(new_n883), .A2(G330), .A3(new_n418), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n908), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n799), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n702), .B2(new_n705), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n1081), .A2(new_n855), .B1(new_n719), .B2(new_n856), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n904), .ZN(new_n1083));
  NOR4_X1   g0883(.A1(new_n843), .A2(KEYINPUT88), .A3(new_n719), .A4(new_n699), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n704), .B1(new_n703), .B2(G330), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n799), .B(new_n855), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n844), .A2(new_n846), .A3(G330), .A4(new_n799), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n848), .A2(new_n851), .B1(new_n339), .B2(new_n853), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n713), .A2(new_n648), .A3(new_n799), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n903), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1086), .A2(new_n1089), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1079), .B1(new_n1083), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1088), .B1(new_n1090), .B2(new_n903), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT114), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n632), .B2(new_n647), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n900), .A2(KEYINPUT114), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1097), .B(new_n1098), .C1(new_n866), .C2(new_n878), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n1095), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n900), .B1(new_n904), .B2(new_n855), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1100), .B(new_n1086), .C1(new_n899), .C2(new_n1101), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n1101), .A2(new_n899), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n856), .A2(new_n719), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n677), .B1(new_n1094), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1079), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n904), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n856), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(G330), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n799), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n1088), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1110), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1093), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1109), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1117), .A2(new_n1106), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n1108), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n727), .B1(new_n287), .B2(new_n806), .ZN(new_n1120));
  NOR3_X1   g0920(.A1(new_n748), .A2(KEYINPUT53), .A3(new_n395), .ZN(new_n1121));
  OAI21_X1  g0921(.A(KEYINPUT53), .B1(new_n748), .B2(new_n395), .ZN(new_n1122));
  XOR2_X1   g0922(.A(KEYINPUT54), .B(G143), .Z(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1122), .B(new_n270), .C1(new_n811), .C2(new_n1124), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1121), .B(new_n1125), .C1(G159), .C2(new_n774), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n825), .A2(new_n745), .B1(new_n749), .B2(new_n940), .ZN(new_n1127));
  INV_X1    g0927(.A(G128), .ZN(new_n1128));
  INV_X1    g0928(.A(G125), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n743), .A2(new_n1128), .B1(new_n757), .B2(new_n1129), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1127), .B(new_n1130), .C1(new_n737), .C2(G50), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n743), .A2(new_n767), .B1(new_n811), .B2(new_n239), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n749), .A2(new_n237), .B1(new_n757), .B2(new_n421), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n267), .B1(new_n753), .B2(new_n280), .C1(new_n455), .C2(new_n745), .ZN(new_n1134));
  NOR3_X1   g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n809), .A2(G87), .B1(G68), .B2(new_n737), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1126), .A2(new_n1131), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1120), .B1(new_n951), .B2(new_n1137), .C1(new_n899), .C2(new_n788), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1102), .A2(new_n1105), .A3(new_n725), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(KEYINPUT115), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT115), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1102), .A2(new_n1105), .A3(new_n1142), .A4(new_n725), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1139), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1119), .A2(new_n1144), .ZN(G378));
  AOI21_X1  g0945(.A(new_n1091), .B1(new_n1081), .B2(new_n855), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n904), .A2(new_n1082), .B1(new_n1146), .B2(new_n1089), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1109), .B1(new_n1147), .B2(new_n1106), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(KEYINPUT57), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT116), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n417), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n401), .A2(new_n645), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n409), .A2(KEYINPUT116), .A3(new_n410), .A4(new_n416), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1154), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1156), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1152), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n1155), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1154), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n1151), .A3(new_n1163), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n879), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n883), .A2(new_n799), .A3(new_n1166), .A4(new_n855), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1167), .A2(KEYINPUT40), .B1(new_n1111), .B2(new_n887), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1165), .B1(new_n1168), .B2(new_n719), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n907), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1165), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n889), .A2(G330), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1171), .B1(new_n889), .B2(G330), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n719), .B(new_n1165), .C1(new_n880), .C2(new_n888), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n907), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n678), .B1(new_n1150), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1148), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT117), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1173), .A2(new_n1176), .A3(KEYINPUT117), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1179), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1178), .B1(new_n1183), .B2(KEYINPUT57), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1165), .A2(new_n787), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n728), .B1(G50), .B2(new_n807), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n675), .A2(new_n270), .ZN(new_n1188));
  AOI211_X1 g0988(.A(G50), .B(new_n1188), .C1(new_n262), .C2(new_n258), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n765), .A2(G107), .B1(new_n742), .B2(G116), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1190), .B1(new_n767), .B2(new_n757), .C1(new_n736), .C2(new_n349), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1188), .B1(new_n748), .B2(new_n280), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n811), .A2(new_n294), .B1(new_n239), .B2(new_n749), .ZN(new_n1193));
  OR4_X1    g0993(.A1(new_n942), .A2(new_n1191), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT58), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1189), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n1128), .A2(new_n745), .B1(new_n749), .B2(new_n825), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n747), .A2(new_n1123), .B1(new_n755), .B2(G137), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n1129), .B2(new_n743), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1197), .B(new_n1199), .C1(G150), .C2(new_n774), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT59), .Z(new_n1201));
  AOI211_X1 g1001(.A(G33), .B(G41), .C1(new_n761), .C2(G124), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n736), .B2(new_n352), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1196), .B1(new_n1195), .B2(new_n1194), .C1(new_n1201), .C2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1187), .B1(new_n1204), .B2(new_n778), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1185), .A2(new_n725), .B1(new_n1186), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1184), .A2(new_n1206), .ZN(G375));
  INV_X1    g1007(.A(new_n1147), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1088), .A2(new_n787), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n270), .B1(new_n753), .B2(new_n202), .C1(new_n743), .C2(new_n825), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n1124), .A2(new_n749), .B1(new_n940), .B2(new_n745), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n811), .A2(new_n395), .B1(new_n757), .B2(new_n1128), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n809), .A2(G159), .B1(G58), .B2(new_n737), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n809), .A2(G97), .B1(G77), .B2(new_n737), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1017), .B(new_n267), .C1(new_n455), .C2(new_n749), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n743), .A2(new_n421), .B1(new_n745), .B2(new_n767), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n811), .A2(new_n237), .B1(new_n757), .B2(new_n768), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1213), .A2(new_n1214), .B1(new_n1215), .B2(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1220), .A2(new_n951), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n727), .B(new_n1221), .C1(new_n314), .C2(new_n806), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1208), .A2(new_n725), .B1(new_n1209), .B2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1083), .A2(new_n1079), .A3(new_n1093), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1117), .A2(new_n981), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1225), .ZN(G381));
  NOR2_X1   g1026(.A1(G375), .A2(G378), .ZN(new_n1227));
  INV_X1    g1027(.A(G384), .ZN(new_n1228));
  INV_X1    g1028(.A(G390), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1037), .B(new_n794), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1231));
  NOR4_X1   g1031(.A1(new_n1230), .A2(G387), .A3(G381), .A4(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1227), .A2(new_n1232), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT118), .ZN(G407));
  INV_X1    g1034(.A(G213), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n1227), .B2(new_n646), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1233), .A2(KEYINPUT118), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1233), .A2(KEYINPUT118), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1236), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT119), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(G407), .A2(KEYINPUT119), .A3(new_n1236), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(G409));
  INV_X1    g1043(.A(new_n954), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n980), .A2(new_n981), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n722), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n997), .A2(new_n1002), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1244), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(KEYINPUT123), .B1(new_n1248), .B2(G390), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(G393), .A2(G396), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1231), .ZN(new_n1251));
  OAI211_X1 g1051(.A(G390), .B(new_n954), .C1(new_n982), .C2(new_n1003), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1229), .A2(G387), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1249), .A2(new_n1251), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT123), .ZN(new_n1255));
  AND4_X1   g1055(.A1(new_n1255), .A2(new_n1253), .A3(new_n1252), .A4(new_n1251), .ZN(new_n1256));
  OR2_X1    g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  XOR2_X1   g1057(.A(new_n1257), .B(KEYINPUT126), .Z(new_n1258));
  AND2_X1   g1058(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n677), .B1(new_n1259), .B2(new_n1149), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1173), .A2(new_n1176), .A3(KEYINPUT117), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT117), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1148), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT57), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1260), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n725), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1186), .A2(new_n1205), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(G378), .B1(new_n1265), .B2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT60), .B1(new_n1147), .B2(new_n1079), .ZN(new_n1270));
  OAI21_X1  g1070(.A(KEYINPUT120), .B1(new_n1270), .B2(new_n1094), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1147), .A2(KEYINPUT60), .A3(new_n1079), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT121), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n678), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1147), .A2(KEYINPUT121), .A3(KEYINPUT60), .A4(new_n1079), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT60), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1224), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT120), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1277), .A2(new_n1278), .A3(new_n1117), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1271), .A2(new_n1274), .A3(new_n1275), .A4(new_n1279), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1280), .A2(G384), .A3(new_n1223), .ZN(new_n1281));
  AOI21_X1  g1081(.A(G384), .B1(new_n1280), .B2(new_n1223), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1144), .B(new_n1267), .C1(new_n1108), .C2(new_n1118), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n722), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n981), .B(new_n1148), .C1(new_n1261), .C2(new_n1262), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1286), .A2(new_n1287), .B1(G213), .B2(new_n646), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1269), .A2(new_n1283), .A3(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT122), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT62), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1269), .A2(new_n1283), .A3(KEYINPUT122), .A4(new_n1288), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1289), .A2(KEYINPUT62), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT61), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1282), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1280), .A2(G384), .A3(new_n1223), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n646), .A2(G213), .A3(G2897), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1297), .A2(new_n1298), .A3(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1299), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1302));
  INV_X1    g1102(.A(G378), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1303), .B1(new_n1184), .B2(new_n1206), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n646), .A2(G213), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1300), .B(new_n1302), .C1(new_n1304), .C2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1295), .A2(new_n1296), .A3(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1258), .B1(new_n1294), .B2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT125), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT63), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1307), .B1(G375), .B2(G378), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT122), .B1(new_n1313), .B2(new_n1283), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1293), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1312), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1296), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(KEYINPUT124), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT124), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1319), .B(new_n1296), .C1(new_n1254), .C2(new_n1256), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1269), .A2(new_n1283), .A3(KEYINPUT63), .A4(new_n1288), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1308), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1311), .B1(new_n1316), .B2(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(KEYINPUT63), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1326));
  NOR3_X1   g1126(.A1(new_n1326), .A2(KEYINPUT125), .A3(new_n1323), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1310), .B1(new_n1325), .B2(new_n1327), .ZN(G405));
  NOR2_X1   g1128(.A1(new_n1227), .A2(new_n1304), .ZN(new_n1329));
  OR2_X1    g1129(.A1(new_n1329), .A2(new_n1257), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1257), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT127), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1283), .A2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1332), .A2(new_n1334), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1330), .A2(new_n1333), .A3(new_n1283), .A4(new_n1331), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(G402));
endmodule


