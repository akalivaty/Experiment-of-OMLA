//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n202), .A2(new_n203), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n210), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n212), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n215), .B(new_n221), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n201), .A2(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n203), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n241), .B(new_n246), .ZN(G351));
  NAND3_X1  g0047(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G116), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n209), .A2(G33), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n248), .A2(new_n252), .A3(new_n219), .A4(new_n253), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n253), .A2(new_n219), .B1(G20), .B2(new_n250), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G283), .ZN(new_n256));
  INV_X1    g0056(.A(G97), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n256), .B(new_n210), .C1(G33), .C2(new_n257), .ZN(new_n258));
  AND3_X1   g0058(.A1(new_n255), .A2(KEYINPUT20), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(KEYINPUT20), .B1(new_n255), .B2(new_n258), .ZN(new_n260));
  OAI221_X1 g0060(.A(new_n251), .B1(new_n250), .B2(new_n254), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT21), .ZN(new_n262));
  INV_X1    g0062(.A(G169), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT78), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G1), .A3(G13), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G274), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(G1), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT5), .A2(G41), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(KEYINPUT5), .A2(G41), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n269), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n264), .B1(new_n267), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n209), .A2(G45), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT5), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n275), .B1(new_n278), .B2(new_n270), .ZN(new_n279));
  INV_X1    g0079(.A(G274), .ZN(new_n280));
  INV_X1    g0080(.A(new_n219), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n280), .B1(new_n281), .B2(new_n265), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n279), .A2(new_n282), .A3(KEYINPUT78), .ZN(new_n283));
  INV_X1    g0083(.A(new_n266), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n274), .A2(new_n283), .B1(new_n285), .B2(G270), .ZN(new_n286));
  INV_X1    g0086(.A(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT3), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G33), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n288), .A2(new_n290), .A3(G264), .A4(G1698), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n288), .A2(new_n290), .A3(G257), .A4(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G303), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT3), .B(G33), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n291), .B(new_n293), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n284), .ZN(new_n297));
  AOI211_X1 g0097(.A(new_n262), .B(new_n263), .C1(new_n286), .C2(new_n297), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n286), .A2(G179), .A3(new_n297), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n261), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n274), .A2(new_n283), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n285), .A2(G270), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n297), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n261), .B1(new_n303), .B2(G200), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n304), .B1(new_n305), .B2(new_n303), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n303), .A2(new_n261), .A3(G169), .ZN(new_n307));
  AND3_X1   g0107(.A1(new_n307), .A2(KEYINPUT81), .A3(new_n262), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT81), .B1(new_n307), .B2(new_n262), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n300), .B(new_n306), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n253), .A2(new_n219), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n248), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT64), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n249), .A2(new_n312), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT64), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n209), .A2(G20), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(G50), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n249), .A2(new_n201), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT8), .B(G58), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n210), .A2(G33), .ZN(new_n324));
  INV_X1    g0124(.A(G150), .ZN(new_n325));
  NOR2_X1   g0125(.A1(G20), .A2(G33), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n323), .A2(new_n324), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(G20), .B2(new_n204), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n321), .B(new_n322), .C1(new_n313), .C2(new_n329), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT9), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n295), .A2(G222), .A3(new_n292), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n295), .A2(G223), .A3(G1698), .ZN(new_n333));
  INV_X1    g0133(.A(G77), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n332), .B(new_n333), .C1(new_n334), .C2(new_n295), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n284), .ZN(new_n336));
  AOI21_X1  g0136(.A(G1), .B1(new_n277), .B2(new_n268), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(new_n266), .A3(G274), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n284), .A2(new_n337), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n339), .B1(G226), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n342), .A2(new_n305), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(G200), .B2(new_n342), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n331), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT10), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT10), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n331), .A2(new_n347), .A3(new_n344), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n342), .A2(new_n263), .ZN(new_n349));
  AND2_X1   g0149(.A1(KEYINPUT65), .A2(G179), .ZN(new_n350));
  NOR2_X1   g0150(.A1(KEYINPUT65), .A2(G179), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n330), .B(new_n349), .C1(new_n353), .C2(new_n342), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT66), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n354), .A2(new_n355), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n346), .A2(new_n348), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n288), .A2(new_n290), .A3(G226), .A4(G1698), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n288), .A2(new_n290), .A3(G223), .A4(new_n292), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G33), .A2(G87), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n284), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n266), .A2(G232), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n338), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  AND3_X1   g0167(.A1(new_n363), .A2(new_n353), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n263), .B1(new_n363), .B2(new_n367), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT73), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n363), .A2(new_n367), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G169), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n366), .B1(new_n284), .B2(new_n362), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n353), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT73), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n288), .A2(new_n290), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT7), .B1(new_n377), .B2(new_n210), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT7), .ZN(new_n379));
  AOI211_X1 g0179(.A(new_n379), .B(G20), .C1(new_n288), .C2(new_n290), .ZN(new_n380));
  OAI21_X1  g0180(.A(G68), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT16), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G58), .A2(G68), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT72), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT72), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(G58), .A3(G68), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n386), .A3(new_n216), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n387), .A2(G20), .B1(G159), .B2(new_n326), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n381), .A2(new_n382), .A3(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n379), .B1(new_n295), .B2(G20), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n289), .A2(G33), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n287), .A2(KEYINPUT3), .ZN(new_n392));
  OAI211_X1 g0192(.A(KEYINPUT7), .B(new_n210), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n203), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n387), .A2(G20), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n326), .A2(G159), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT16), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n313), .B1(new_n389), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT8), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G58), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n319), .A2(new_n403), .A3(new_n320), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n403), .A2(new_n248), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  OAI22_X1  g0207(.A1(new_n371), .A2(new_n376), .B1(new_n399), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT18), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n389), .A2(new_n398), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n312), .ZN(new_n411));
  INV_X1    g0211(.A(new_n407), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n370), .B1(new_n368), .B2(new_n369), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n373), .A2(KEYINPUT73), .A3(new_n375), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT18), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n413), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n363), .A2(G190), .A3(new_n367), .ZN(new_n419));
  INV_X1    g0219(.A(G200), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n419), .B1(new_n420), .B2(new_n374), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n411), .A2(new_n412), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT17), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n399), .A2(new_n407), .A3(new_n421), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT17), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n409), .A2(new_n418), .A3(new_n425), .A4(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n320), .A2(G77), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n314), .A2(new_n430), .B1(G77), .B2(new_n248), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT68), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n403), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n323), .A2(KEYINPUT68), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n327), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  XNOR2_X1  g0235(.A(KEYINPUT15), .B(G87), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n436), .A2(new_n324), .B1(new_n210), .B2(new_n334), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n312), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT69), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g0240(.A(KEYINPUT69), .B(new_n312), .C1(new_n435), .C2(new_n437), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n431), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n295), .A2(G232), .A3(new_n292), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n295), .A2(G238), .A3(G1698), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n377), .A2(G107), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n284), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n339), .B1(G244), .B2(new_n340), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT67), .ZN(new_n450));
  AOI21_X1  g0250(.A(KEYINPUT67), .B1(new_n448), .B2(new_n449), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n352), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n448), .A2(new_n449), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT67), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT67), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n263), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n443), .A2(new_n452), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(G190), .B1(new_n450), .B2(new_n451), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n455), .A2(G200), .A3(new_n456), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n460), .A3(new_n442), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g0262(.A(new_n462), .B(KEYINPUT70), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n295), .A2(G232), .A3(G1698), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G97), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n288), .A2(new_n290), .A3(G226), .A4(new_n292), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n284), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT13), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n340), .A2(G238), .B1(new_n282), .B2(new_n337), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n469), .B1(new_n468), .B2(new_n470), .ZN(new_n472));
  OAI21_X1  g0272(.A(G200), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI22_X1  g0273(.A1(new_n324), .A2(new_n334), .B1(new_n210), .B2(G68), .ZN(new_n474));
  OAI22_X1  g0274(.A1(new_n474), .A2(KEYINPUT71), .B1(new_n201), .B2(new_n327), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n474), .A2(KEYINPUT71), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n312), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT11), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT12), .B1(new_n248), .B2(G68), .ZN(new_n480));
  OR3_X1    g0280(.A1(new_n248), .A2(KEYINPUT12), .A3(G68), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n203), .B1(new_n209), .B2(G20), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n480), .A2(new_n481), .B1(new_n316), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n477), .B2(new_n478), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n468), .A2(new_n470), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT13), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n487), .A2(G190), .A3(new_n488), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n473), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(G169), .B1(new_n471), .B2(new_n472), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT14), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n487), .A2(G179), .A3(new_n488), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT14), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n494), .B(G169), .C1(new_n471), .C2(new_n472), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n492), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n485), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n490), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n358), .A2(new_n429), .A3(new_n463), .A4(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  AND2_X1   g0300(.A1(G97), .A2(G107), .ZN(new_n501));
  OAI22_X1  g0301(.A1(new_n501), .A2(new_n206), .B1(KEYINPUT74), .B2(KEYINPUT6), .ZN(new_n502));
  NOR2_X1   g0302(.A1(KEYINPUT74), .A2(KEYINPUT6), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(KEYINPUT6), .B2(new_n257), .ZN(new_n504));
  XNOR2_X1  g0304(.A(G97), .B(G107), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n502), .B(G20), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n326), .A2(G77), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(G107), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n509), .B1(new_n390), .B2(new_n393), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n312), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n254), .A2(new_n257), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT75), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n248), .B2(G97), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n249), .A2(KEYINPUT75), .A3(new_n257), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(KEYINPUT76), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n511), .A2(new_n516), .A3(KEYINPUT76), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n288), .A2(new_n290), .A3(G250), .A4(G1698), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n288), .A2(new_n290), .A3(G244), .A4(new_n292), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT4), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n256), .B(new_n520), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT77), .B1(new_n521), .B2(new_n522), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n521), .A2(KEYINPUT77), .A3(new_n522), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n266), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n285), .A2(G257), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n301), .A2(new_n528), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n527), .A2(G190), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n521), .A2(new_n522), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT77), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OR2_X1    g0333(.A1(new_n521), .A2(new_n522), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n520), .A2(new_n256), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n533), .A2(new_n534), .A3(new_n526), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n284), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n301), .A2(new_n528), .ZN(new_n538));
  AOI21_X1  g0338(.A(G200), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n518), .B(new_n519), .C1(new_n530), .C2(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(G169), .B1(new_n527), .B2(new_n529), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n537), .A2(new_n538), .A3(new_n353), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n511), .A2(new_n516), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT19), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n210), .B1(new_n465), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(G87), .B2(new_n207), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n288), .A2(new_n290), .A3(new_n210), .A4(G68), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n546), .B1(new_n324), .B2(new_n257), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n551), .A2(new_n312), .B1(new_n249), .B2(new_n436), .ZN(new_n552));
  INV_X1    g0352(.A(G87), .ZN(new_n553));
  OR3_X1    g0353(.A1(new_n254), .A2(KEYINPUT80), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT80), .B1(new_n254), .B2(new_n553), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n288), .A2(new_n290), .A3(G244), .A4(G1698), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n288), .A2(new_n290), .A3(G238), .A4(new_n292), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n558), .B(new_n559), .C1(new_n287), .C2(new_n250), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n284), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n282), .A2(new_n269), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT79), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n275), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n209), .A2(KEYINPUT79), .A3(G45), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n564), .A2(G250), .A3(new_n266), .A4(new_n565), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G200), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n561), .A2(new_n567), .A3(G190), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n557), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n552), .B1(new_n254), .B2(new_n436), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n568), .A2(new_n263), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n561), .A2(new_n567), .A3(new_n352), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n540), .A2(new_n545), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n295), .A2(new_n210), .A3(G87), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT22), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT22), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n295), .A2(new_n580), .A3(new_n210), .A4(G87), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT24), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n287), .A2(new_n250), .A3(G20), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n210), .A2(G107), .ZN(new_n585));
  OR2_X1    g0385(.A1(new_n585), .A2(KEYINPUT23), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(KEYINPUT23), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n584), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n582), .A2(new_n583), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n583), .B1(new_n582), .B2(new_n588), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n312), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(G13), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n593), .A2(G1), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n585), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT82), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT25), .ZN(new_n597));
  OR2_X1    g0397(.A1(new_n596), .A2(KEYINPUT25), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(KEYINPUT25), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n598), .A2(new_n594), .A3(new_n585), .A4(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n597), .B(new_n600), .C1(new_n509), .C2(new_n254), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT83), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n285), .A2(new_n603), .A3(G264), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n273), .A2(G264), .A3(new_n266), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT83), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n295), .A2(G257), .A3(G1698), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n295), .A2(G250), .A3(new_n292), .ZN(new_n608));
  NAND2_X1  g0408(.A1(G33), .A2(G294), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n604), .A2(new_n606), .B1(new_n610), .B2(new_n284), .ZN(new_n611));
  AOI21_X1  g0411(.A(G200), .B1(new_n611), .B2(new_n301), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n284), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n613), .A2(new_n301), .A3(new_n605), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n614), .A2(G190), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n592), .B(new_n602), .C1(new_n612), .C2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(G169), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n604), .A2(new_n606), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n618), .A2(G179), .A3(new_n301), .A4(new_n613), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n582), .A2(new_n588), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT24), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n313), .B1(new_n622), .B2(new_n589), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n620), .B1(new_n623), .B2(new_n601), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n616), .A2(new_n624), .ZN(new_n625));
  AND4_X1   g0425(.A1(new_n311), .A2(new_n500), .A3(new_n577), .A4(new_n625), .ZN(G372));
  NAND2_X1  g0426(.A1(new_n357), .A2(new_n356), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n346), .A2(new_n348), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n409), .A2(new_n418), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n495), .A2(new_n493), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n487), .A2(new_n488), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n494), .B1(new_n632), .B2(G169), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n497), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n490), .B2(new_n458), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n425), .A2(new_n427), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n630), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n627), .B1(new_n629), .B2(new_n637), .ZN(new_n638));
  XOR2_X1   g0438(.A(new_n638), .B(KEYINPUT86), .Z(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NOR3_X1   g0440(.A1(new_n527), .A2(new_n529), .A3(new_n352), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n263), .B1(new_n537), .B2(new_n538), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n511), .A2(new_n516), .A3(KEYINPUT76), .ZN(new_n643));
  OAI22_X1  g0443(.A1(new_n641), .A2(new_n642), .B1(new_n643), .B2(new_n517), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n571), .A2(new_n575), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT84), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n541), .A2(new_n542), .B1(new_n511), .B2(new_n516), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n576), .A2(new_n648), .A3(KEYINPUT26), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT85), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT84), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n651), .B(new_n640), .C1(new_n644), .C2(new_n645), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT85), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n576), .A2(new_n648), .A3(new_n653), .A4(KEYINPUT26), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n647), .A2(new_n650), .A3(new_n652), .A4(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n575), .ZN(new_n656));
  AND4_X1   g0456(.A1(new_n545), .A2(new_n540), .A3(new_n576), .A4(new_n616), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n624), .B(new_n300), .C1(new_n309), .C2(new_n308), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n500), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n639), .A2(new_n661), .ZN(G369));
  OAI21_X1  g0462(.A(new_n300), .B1(new_n308), .B2(new_n309), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n594), .A2(new_n210), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n664), .A2(KEYINPUT87), .A3(KEYINPUT27), .ZN(new_n665));
  AOI21_X1  g0465(.A(KEYINPUT87), .B1(new_n664), .B2(KEYINPUT27), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(G213), .B1(new_n664), .B2(KEYINPUT27), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n261), .ZN(new_n673));
  MUX2_X1   g0473(.A(new_n663), .B(new_n311), .S(new_n673), .Z(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n672), .B1(new_n623), .B2(new_n601), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n625), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n672), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n678), .B1(new_n624), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n663), .A2(new_n679), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n625), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n624), .A2(new_n672), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n681), .A2(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n658), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n540), .A2(new_n545), .A3(new_n576), .A4(new_n616), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT26), .B1(new_n644), .B2(new_n645), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n576), .A2(new_n648), .A3(new_n640), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(new_n575), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n679), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT89), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI211_X1 g0496(.A(KEYINPUT89), .B(new_n679), .C1(new_n690), .C2(new_n693), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(KEYINPUT29), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n672), .B1(new_n655), .B2(new_n659), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n577), .A2(new_n311), .A3(new_n625), .A4(new_n679), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n297), .A2(new_n301), .A3(new_n302), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n561), .A2(new_n567), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n705), .A2(G179), .A3(new_n706), .A4(new_n611), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n537), .A2(new_n538), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n704), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n706), .A2(new_n611), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n527), .A2(new_n529), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n710), .A2(new_n711), .A3(KEYINPUT30), .A4(new_n299), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n706), .A2(new_n353), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n611), .A2(new_n301), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n713), .A2(new_n708), .A3(new_n303), .A4(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n709), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n672), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT31), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n703), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G330), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT88), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n721), .A2(KEYINPUT88), .A3(G330), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n702), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT90), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n702), .A2(KEYINPUT90), .A3(new_n726), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n729), .A2(new_n209), .A3(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n213), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G41), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(G1), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n217), .B2(new_n734), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n731), .A2(new_n738), .ZN(G364));
  NOR2_X1   g0539(.A1(new_n674), .A2(G330), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT91), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n593), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n209), .B1(new_n742), .B2(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n733), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n741), .A2(new_n675), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n219), .B1(G20), .B2(new_n263), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n210), .A2(new_n420), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n353), .A2(G190), .A3(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n353), .A2(new_n305), .A3(new_n749), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(KEYINPUT33), .B(G317), .ZN(new_n754));
  AOI22_X1  g0554(.A1(G326), .A2(new_n751), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G311), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n210), .A2(G190), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n353), .A2(new_n420), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n210), .A2(new_n305), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n420), .A2(G179), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT93), .Z(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n755), .B1(new_n756), .B2(new_n758), .C1(new_n294), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n757), .A2(new_n760), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G179), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n757), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(G283), .A2(new_n766), .B1(new_n769), .B2(G329), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT94), .Z(new_n771));
  NAND2_X1  g0571(.A1(new_n767), .A2(G190), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G294), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n353), .A2(new_n420), .A3(new_n759), .ZN(new_n776));
  INV_X1    g0576(.A(G322), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n377), .B1(new_n774), .B2(new_n775), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n764), .A2(new_n771), .A3(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n758), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G68), .A2(new_n753), .B1(new_n780), .B2(G77), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n201), .B2(new_n750), .ZN(new_n782));
  INV_X1    g0582(.A(G159), .ZN(new_n783));
  OR3_X1    g0583(.A1(new_n768), .A2(KEYINPUT32), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(KEYINPUT32), .B1(new_n768), .B2(new_n783), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n784), .B(new_n785), .C1(new_n257), .C2(new_n774), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n776), .A2(new_n202), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n295), .B1(new_n765), .B2(new_n509), .C1(new_n553), .C2(new_n761), .ZN(new_n788));
  NOR4_X1   g0588(.A1(new_n782), .A2(new_n786), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n748), .B1(new_n779), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n213), .A2(G355), .A3(new_n295), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n732), .A2(new_n295), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(G45), .B2(new_n217), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n246), .A2(new_n268), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n791), .B1(G116), .B2(new_n213), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G13), .A2(G33), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n748), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT92), .Z(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n746), .B1(new_n795), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n790), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT95), .ZN(new_n804));
  INV_X1    g0604(.A(new_n798), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n674), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n747), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G396));
  NAND4_X1  g0608(.A1(new_n443), .A2(new_n679), .A3(new_n452), .A4(new_n457), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n443), .A2(new_n672), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n461), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n810), .B1(new_n458), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n700), .B(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n745), .B1(new_n814), .B2(new_n726), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n726), .B2(new_n814), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n748), .A2(new_n796), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n746), .B1(new_n334), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n776), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G294), .A2(new_n819), .B1(new_n780), .B2(G116), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n294), .B2(new_n750), .ZN(new_n821));
  INV_X1    g0621(.A(G283), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n763), .A2(new_n509), .B1(new_n822), .B2(new_n752), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n774), .A2(new_n257), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n377), .B1(new_n768), .B2(new_n756), .C1(new_n553), .C2(new_n765), .ZN(new_n825));
  NOR4_X1   g0625(.A1(new_n821), .A2(new_n823), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G137), .A2(new_n751), .B1(new_n753), .B2(G150), .ZN(new_n827));
  INV_X1    g0627(.A(G143), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n827), .B1(new_n828), .B2(new_n776), .C1(new_n783), .C2(new_n758), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT34), .Z(new_n830));
  AOI21_X1  g0630(.A(new_n377), .B1(new_n769), .B2(G132), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n765), .A2(new_n203), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n762), .B2(G50), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT96), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n831), .B1(new_n202), .B2(new_n774), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n830), .B1(KEYINPUT97), .B2(new_n837), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n837), .A2(KEYINPUT97), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n826), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n748), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n818), .B1(new_n797), .B2(new_n813), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n816), .A2(new_n842), .ZN(G384));
  NOR2_X1   g0643(.A1(new_n742), .A2(new_n209), .ZN(new_n844));
  INV_X1    g0644(.A(G330), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n812), .A2(new_n458), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n809), .ZN(new_n847));
  INV_X1    g0647(.A(new_n490), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n497), .A2(new_n672), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n634), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n497), .B(new_n672), .C1(new_n496), .C2(new_n490), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n847), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n721), .A2(new_n852), .A3(KEYINPUT40), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT100), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n669), .B1(new_n399), .B2(new_n407), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n408), .A2(new_n423), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n854), .B1(new_n856), .B2(KEYINPUT37), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n426), .B1(new_n413), .B2(new_n416), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT101), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g0661(.A(KEYINPUT101), .B(new_n669), .C1(new_n399), .C2(new_n407), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n858), .A2(new_n859), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n857), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n855), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n428), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n856), .A2(new_n854), .A3(KEYINPUT37), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n864), .A2(KEYINPUT38), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n861), .A2(new_n862), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n408), .A2(new_n423), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT37), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n871), .A2(new_n863), .B1(new_n428), .B2(new_n869), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n868), .B1(KEYINPUT38), .B2(new_n872), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n853), .A2(new_n873), .A3(KEYINPUT103), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT103), .B1(new_n853), .B2(new_n873), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT40), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n850), .A2(new_n851), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n813), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n719), .A2(new_n720), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n879), .B1(new_n703), .B2(new_n880), .ZN(new_n881));
  AND4_X1   g0681(.A1(KEYINPUT38), .A2(new_n864), .A3(new_n867), .A4(new_n866), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n859), .B1(new_n858), .B2(new_n855), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n854), .A2(new_n883), .B1(new_n428), .B2(new_n865), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT38), .B1(new_n884), .B2(new_n864), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n881), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n876), .B1(new_n877), .B2(new_n886), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT104), .Z(new_n888));
  AOI21_X1  g0688(.A(new_n499), .B1(new_n703), .B2(new_n880), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n845), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n889), .B2(new_n888), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n810), .B1(new_n700), .B2(new_n813), .ZN(new_n892));
  INV_X1    g0692(.A(new_n878), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT99), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n866), .A2(new_n867), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n857), .A2(new_n863), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n868), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT99), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n672), .B(new_n847), .C1(new_n655), .C2(new_n659), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n900), .B(new_n878), .C1(new_n901), .C2(new_n810), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n894), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT39), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n872), .A2(KEYINPUT38), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n904), .B1(new_n882), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n898), .A2(KEYINPUT39), .A3(new_n868), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n496), .A2(new_n497), .A3(new_n679), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n630), .A2(new_n670), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n903), .A2(KEYINPUT102), .A3(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT102), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n910), .A2(new_n911), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n894), .A2(new_n899), .A3(new_n902), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n699), .A2(new_n500), .A3(new_n701), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n639), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n918), .B(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n844), .B1(new_n891), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n891), .B2(new_n921), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT35), .ZN(new_n925));
  OAI211_X1 g0725(.A(G116), .B(new_n220), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n925), .B2(new_n924), .ZN(new_n927));
  XNOR2_X1  g0727(.A(KEYINPUT98), .B(KEYINPUT36), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n927), .B(new_n928), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n218), .A2(G77), .A3(new_n386), .A4(new_n384), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n242), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(G1), .A3(new_n593), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n923), .A2(new_n929), .A3(new_n932), .ZN(G367));
  NAND3_X1  g0733(.A1(new_n762), .A2(KEYINPUT46), .A3(G116), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT107), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n775), .A2(new_n752), .B1(new_n750), .B2(new_n756), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n822), .A2(new_n758), .B1(new_n776), .B2(new_n294), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n934), .A2(new_n935), .ZN(new_n940));
  INV_X1    g0740(.A(new_n761), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT46), .B1(new_n941), .B2(G116), .ZN(new_n942));
  INV_X1    g0742(.A(G317), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n377), .B1(new_n768), .B2(new_n943), .C1(new_n257), .C2(new_n765), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n942), .B(new_n944), .C1(G107), .C2(new_n773), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n936), .A2(new_n939), .A3(new_n940), .A4(new_n945), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n201), .A2(new_n758), .B1(new_n752), .B2(new_n783), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(KEYINPUT108), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n295), .B1(new_n761), .B2(new_n202), .ZN(new_n949));
  INV_X1    g0749(.A(G137), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n765), .A2(new_n334), .B1(new_n768), .B2(new_n950), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n949), .B(new_n951), .C1(G68), .C2(new_n773), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n947), .A2(KEYINPUT108), .ZN(new_n953));
  AOI22_X1  g0753(.A1(G143), .A2(new_n751), .B1(new_n819), .B2(G150), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n946), .B1(new_n948), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT47), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n748), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n576), .B1(new_n557), .B2(new_n679), .ZN(new_n959));
  OR3_X1    g0759(.A1(new_n575), .A2(new_n679), .A3(new_n557), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n798), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n213), .A2(new_n436), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n800), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n792), .A2(new_n237), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n746), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n958), .A2(new_n963), .A3(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n730), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT90), .B1(new_n702), .B2(new_n726), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n518), .A2(new_n519), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n672), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(new_n540), .A3(new_n545), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n971), .A2(new_n543), .A3(new_n672), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n685), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT44), .ZN(new_n978));
  XOR2_X1   g0778(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n979));
  NAND3_X1  g0779(.A1(new_n686), .A2(new_n975), .A3(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n979), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n685), .B2(new_n976), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n676), .B(new_n680), .C1(new_n978), .C2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT44), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n977), .B(new_n985), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n986), .A2(new_n681), .A3(new_n980), .A4(new_n982), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n683), .B1(new_n680), .B2(new_n682), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(KEYINPUT106), .B2(new_n675), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n675), .A2(KEYINPUT106), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n990), .B(new_n991), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n969), .A2(new_n970), .B1(new_n988), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n733), .B(KEYINPUT41), .Z(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n744), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n976), .A2(new_n683), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT42), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n545), .B1(new_n976), .B2(new_n624), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n679), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT43), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n962), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1001), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n681), .A2(new_n976), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n998), .A2(new_n1002), .A3(new_n962), .A4(new_n1000), .ZN(new_n1007));
  AND3_X1   g0807(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1006), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n968), .B1(new_n996), .B2(new_n1011), .ZN(G387));
  INV_X1    g0812(.A(new_n992), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n969), .B2(new_n970), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n729), .A2(new_n730), .A3(new_n992), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1014), .A2(new_n733), .A3(new_n1015), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n756), .A2(new_n752), .B1(new_n750), .B2(new_n777), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1017), .A2(KEYINPUT111), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(KEYINPUT111), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G317), .A2(new_n819), .B1(new_n780), .B2(G303), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT48), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n941), .A2(G294), .B1(new_n773), .B2(G283), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT49), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n765), .A2(new_n250), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n295), .B(new_n1030), .C1(G326), .C2(new_n769), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n941), .A2(G77), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n325), .B2(new_n768), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n774), .A2(new_n436), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n295), .B1(new_n765), .B2(new_n257), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n403), .A2(new_n753), .B1(new_n780), .B2(G68), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G50), .A2(new_n819), .B1(new_n751), .B2(G159), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n841), .B1(new_n1032), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n433), .A2(new_n434), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n201), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT50), .Z(new_n1044));
  INV_X1    g0844(.A(KEYINPUT110), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n735), .A2(KEYINPUT109), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n735), .A2(KEYINPUT109), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n268), .B1(new_n203), .B2(new_n334), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1044), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1049), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1051), .A2(KEYINPUT110), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n792), .B1(new_n268), .B2(new_n234), .C1(new_n1050), .C2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n213), .A2(new_n295), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1053), .B1(G107), .B2(new_n213), .C1(new_n735), .C2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n746), .B1(new_n1055), .B2(new_n801), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n680), .B2(new_n805), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n992), .A2(new_n743), .B1(new_n1041), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1016), .A2(new_n1059), .ZN(G393));
  AOI21_X1  g0860(.A(new_n992), .B1(new_n729), .B2(new_n730), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n988), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n734), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1014), .A2(new_n988), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1062), .A2(new_n744), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n801), .B1(new_n257), .B2(new_n213), .ZN(new_n1067));
  NOR3_X1   g0867(.A1(new_n241), .A2(new_n732), .A3(new_n295), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n745), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n325), .A2(new_n750), .B1(new_n776), .B2(new_n783), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT51), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n295), .B1(new_n765), .B2(new_n553), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n761), .A2(new_n203), .B1(new_n768), .B2(new_n828), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1072), .B(new_n1073), .C1(G77), .C2(new_n773), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n1042), .A2(new_n780), .B1(new_n753), .B2(G50), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1071), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G283), .A2(new_n941), .B1(new_n769), .B2(G322), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1077), .B(new_n377), .C1(new_n509), .C2(new_n765), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT112), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n753), .A2(G303), .B1(G116), .B2(new_n773), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1079), .B(new_n1080), .C1(new_n775), .C2(new_n758), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n756), .A2(new_n776), .B1(new_n750), .B2(new_n943), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT52), .Z(new_n1083));
  OAI21_X1  g0883(.A(new_n1076), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1069), .B1(new_n1084), .B2(new_n748), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n975), .B2(new_n805), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1066), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1065), .A2(new_n1088), .ZN(G390));
  NOR2_X1   g0889(.A1(new_n722), .A2(new_n879), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n696), .A2(new_n697), .A3(new_n809), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1091), .A2(new_n846), .A3(new_n878), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n873), .A2(new_n908), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n878), .B1(new_n901), .B2(new_n810), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1095), .A2(new_n908), .B1(new_n906), .B2(new_n907), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1090), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n724), .A2(new_n725), .A3(new_n813), .A4(new_n878), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n892), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n909), .B1(new_n1100), .B2(new_n878), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n906), .A2(new_n907), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1098), .B(new_n1099), .C1(new_n1101), .C2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1097), .A2(new_n744), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT114), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1105), .B(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1097), .A2(new_n1104), .ZN(new_n1108));
  OR3_X1    g0908(.A1(new_n722), .A2(new_n499), .A3(KEYINPUT113), .ZN(new_n1109));
  OAI21_X1  g0909(.A(KEYINPUT113), .B1(new_n722), .B2(new_n499), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n919), .A2(new_n1111), .A3(new_n639), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1091), .A2(new_n846), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n893), .B1(new_n722), .B2(new_n847), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1098), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n724), .A2(new_n725), .A3(new_n813), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1090), .B1(new_n1117), .B2(new_n893), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1116), .B1(new_n1118), .B2(new_n892), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1113), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1108), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1097), .A2(new_n1113), .A3(new_n1104), .A4(new_n1119), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1121), .A2(new_n733), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n817), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n745), .B1(new_n403), .B2(new_n1124), .ZN(new_n1125));
  XOR2_X1   g0925(.A(new_n1125), .B(KEYINPUT115), .Z(new_n1126));
  AOI22_X1  g0926(.A1(G116), .A2(new_n819), .B1(new_n780), .B2(G97), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n295), .B(new_n832), .C1(G294), .C2(new_n769), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1127), .B(new_n1128), .C1(new_n334), .C2(new_n774), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n762), .A2(G87), .B1(G107), .B2(new_n753), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n822), .B2(new_n750), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n941), .A2(G150), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1132), .A2(KEYINPUT53), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n819), .A2(G132), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1132), .A2(KEYINPUT53), .B1(G159), .B2(new_n773), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n295), .B1(new_n765), .B2(new_n201), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G125), .B2(new_n769), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .A4(new_n1137), .ZN(new_n1138));
  XOR2_X1   g0938(.A(KEYINPUT54), .B(G143), .Z(new_n1139));
  AOI22_X1  g0939(.A1(G137), .A2(new_n753), .B1(new_n780), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(G128), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1140), .B1(new_n1141), .B2(new_n750), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n1129), .A2(new_n1131), .B1(new_n1138), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1126), .B1(new_n1143), .B2(new_n748), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n1103), .B2(new_n797), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1107), .A2(new_n1123), .A3(new_n1145), .ZN(G378));
  NAND2_X1  g0946(.A1(new_n330), .A2(new_n669), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n628), .A2(new_n354), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1147), .B1(new_n628), .B2(new_n354), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  OR3_X1    g0951(.A1(new_n1148), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1151), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1154), .A2(new_n797), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n750), .A2(new_n250), .B1(new_n774), .B2(new_n203), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT116), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(G58), .A2(new_n766), .B1(new_n769), .B2(G283), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n295), .A2(G41), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n1033), .A3(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n752), .A2(new_n257), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n509), .A2(new_n776), .B1(new_n758), .B2(new_n436), .ZN(new_n1162));
  NOR4_X1   g0962(.A1(new_n1157), .A2(new_n1160), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1163), .A2(KEYINPUT58), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(KEYINPUT58), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1159), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1166), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1164), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n941), .A2(new_n1139), .B1(new_n773), .B2(G150), .ZN(new_n1169));
  INV_X1    g0969(.A(G132), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1169), .B1(new_n1170), .B2(new_n752), .ZN(new_n1171));
  INV_X1    g0971(.A(G125), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n1172), .A2(new_n750), .B1(new_n776), .B2(new_n1141), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1171), .B(new_n1173), .C1(G137), .C2(new_n780), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1177));
  XOR2_X1   g0977(.A(KEYINPUT117), .B(G124), .Z(new_n1178));
  OAI211_X1 g0978(.A(new_n287), .B(new_n277), .C1(new_n1178), .C2(new_n768), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G159), .B2(new_n766), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1176), .A2(new_n1177), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n841), .B1(new_n1168), .B2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n745), .B1(G50), .B2(new_n1124), .ZN(new_n1183));
  NOR3_X1   g0983(.A1(new_n1155), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT118), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n886), .A2(new_n877), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1186), .B(G330), .C1(new_n874), .C2(new_n875), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1154), .A2(KEYINPUT119), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(new_n913), .C2(new_n917), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n915), .A2(new_n914), .A3(new_n916), .ZN(new_n1192));
  OAI21_X1  g0992(.A(KEYINPUT102), .B1(new_n903), .B2(new_n912), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1192), .B(new_n1193), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1191), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1185), .B1(new_n1197), .B2(new_n744), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT57), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n1122), .B2(new_n1113), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n733), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1122), .A2(new_n1113), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT57), .B1(new_n1197), .B2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1198), .B1(new_n1202), .B2(new_n1204), .ZN(G375));
  XOR2_X1   g1005(.A(new_n743), .B(KEYINPUT120), .Z(new_n1206));
  NAND2_X1  g1006(.A1(new_n1119), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n746), .B1(new_n203), .B2(new_n817), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n377), .B1(new_n765), .B2(new_n334), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1209), .B(new_n1035), .C1(G303), .C2(new_n769), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n509), .B2(new_n758), .C1(new_n775), .C2(new_n750), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n762), .A2(G97), .B1(G283), .B2(new_n819), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n250), .B2(new_n752), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n753), .A2(new_n1139), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1214), .B1(new_n950), .B2(new_n776), .C1(new_n763), .C2(new_n783), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n295), .B1(new_n768), .B2(new_n1141), .C1(new_n202), .C2(new_n765), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G50), .B2(new_n773), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n1170), .B2(new_n750), .C1(new_n325), .C2(new_n758), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n1211), .A2(new_n1213), .B1(new_n1215), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT121), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n748), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1208), .B1(new_n1222), .B2(new_n1223), .C1(new_n878), .C2(new_n797), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1207), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT122), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1207), .A2(KEYINPUT122), .A3(new_n1224), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1113), .A2(new_n1119), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1120), .A2(new_n995), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1229), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT123), .ZN(G381));
  NAND3_X1  g1033(.A1(new_n1016), .A2(new_n807), .A3(new_n1059), .ZN(new_n1234));
  OR4_X1    g1034(.A1(G384), .A2(G390), .A3(G387), .A4(new_n1234), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1235), .A2(G381), .A3(G378), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(G375), .A2(KEYINPUT124), .ZN(new_n1237));
  OR2_X1    g1037(.A1(G375), .A2(KEYINPUT124), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(G407));
  AND3_X1   g1039(.A1(new_n1107), .A2(new_n1123), .A3(new_n1145), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n671), .A2(G213), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1238), .A2(new_n1240), .A3(new_n1237), .A4(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(G407), .A2(G213), .A3(new_n1243), .ZN(G409));
  AOI21_X1  g1044(.A(new_n1230), .B1(KEYINPUT60), .B2(new_n1120), .ZN(new_n1245));
  OR2_X1    g1045(.A1(new_n1118), .A2(new_n892), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1246), .A2(KEYINPUT60), .A3(new_n1112), .A4(new_n1116), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n733), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1207), .A2(KEYINPUT122), .A3(new_n1224), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT122), .B1(new_n1207), .B2(new_n1224), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n1245), .A2(new_n1248), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(G384), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1229), .B(G384), .C1(new_n1245), .C2(new_n1248), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1242), .A2(G2897), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1253), .A2(new_n1254), .A3(new_n1256), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(G378), .B(new_n1198), .C1(new_n1202), .C2(new_n1204), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1184), .B1(new_n1197), .B2(new_n1206), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1197), .A2(new_n995), .A3(new_n1203), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1240), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1262), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1241), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT61), .B1(new_n1261), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT63), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(new_n1268), .B2(new_n1255), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n993), .A2(new_n995), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n743), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1010), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(G390), .A2(new_n1274), .A3(new_n968), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT125), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1087), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1276), .B1(G387), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G387), .A2(new_n1277), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G393), .A2(G396), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1234), .ZN(new_n1281));
  AND4_X1   g1081(.A1(new_n1275), .A2(new_n1278), .A3(new_n1279), .A4(new_n1281), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n1275), .A2(new_n1279), .B1(new_n1278), .B2(new_n1281), .ZN(new_n1283));
  OR2_X1    g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1242), .B1(new_n1262), .B2(new_n1266), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1255), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1285), .A2(KEYINPUT63), .A3(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1269), .A2(new_n1271), .A3(new_n1284), .A4(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT62), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1285), .A2(new_n1289), .A3(new_n1286), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT61), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(new_n1285), .B2(new_n1260), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1289), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(new_n1290), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1288), .B1(new_n1294), .B2(new_n1284), .ZN(G405));
  INV_X1    g1095(.A(new_n1262), .ZN(new_n1296));
  AOI22_X1  g1096(.A1(new_n1191), .A2(new_n1196), .B1(new_n1113), .B2(new_n1122), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1201), .B(new_n733), .C1(new_n1297), .C2(KEYINPUT57), .ZN(new_n1298));
  AOI21_X1  g1098(.A(G378), .B1(new_n1298), .B2(new_n1198), .ZN(new_n1299));
  NOR3_X1   g1099(.A1(new_n1296), .A2(new_n1299), .A3(new_n1286), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(G375), .A2(new_n1240), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1255), .B1(new_n1301), .B2(new_n1262), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1284), .B1(new_n1300), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT127), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n1284), .B(KEYINPUT127), .C1(new_n1300), .C2(new_n1302), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1286), .B1(new_n1296), .B2(new_n1299), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1301), .A2(new_n1255), .A3(new_n1262), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1307), .A2(new_n1308), .A3(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT126), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1307), .A2(new_n1308), .A3(new_n1309), .A4(KEYINPUT126), .ZN(new_n1313));
  AOI22_X1  g1113(.A1(new_n1305), .A2(new_n1306), .B1(new_n1312), .B2(new_n1313), .ZN(G402));
endmodule


