

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738;

  BUF_X1 U368 ( .A(n537), .Z(n539) );
  XNOR2_X1 U369 ( .A(n427), .B(KEYINPUT89), .ZN(n548) );
  XNOR2_X1 U370 ( .A(n464), .B(n465), .ZN(n726) );
  INV_X1 U371 ( .A(G953), .ZN(n728) );
  INV_X2 U372 ( .A(G143), .ZN(n410) );
  NOR2_X2 U373 ( .A1(n622), .A2(n710), .ZN(n625) );
  XNOR2_X2 U374 ( .A(n531), .B(n530), .ZN(n533) );
  XNOR2_X1 U375 ( .A(n355), .B(n354), .ZN(n544) );
  XNOR2_X1 U376 ( .A(n505), .B(n504), .ZN(n521) );
  XNOR2_X1 U377 ( .A(n516), .B(KEYINPUT38), .ZN(n658) );
  NAND2_X1 U378 ( .A1(n348), .A2(n392), .ZN(n427) );
  XNOR2_X1 U379 ( .A(n402), .B(n401), .ZN(n523) );
  XNOR2_X1 U380 ( .A(n726), .B(n466), .ZN(n484) );
  XNOR2_X1 U381 ( .A(n484), .B(n485), .ZN(n699) );
  XOR2_X1 U382 ( .A(G137), .B(KEYINPUT72), .Z(n492) );
  XNOR2_X1 U383 ( .A(G101), .B(KEYINPUT67), .ZN(n414) );
  XNOR2_X1 U384 ( .A(n673), .B(n477), .ZN(n524) );
  OR2_X2 U385 ( .A1(n699), .A2(G902), .ZN(n385) );
  NOR2_X1 U386 ( .A1(n463), .A2(n351), .ZN(n368) );
  NAND2_X1 U387 ( .A1(n370), .A2(n369), .ZN(n366) );
  XNOR2_X1 U388 ( .A(G122), .B(G116), .ZN(n417) );
  INV_X1 U389 ( .A(G146), .ZN(n466) );
  NOR2_X1 U390 ( .A1(n521), .A2(n634), .ZN(n532) );
  XNOR2_X1 U391 ( .A(n468), .B(G137), .ZN(n377) );
  AND2_X1 U392 ( .A1(n544), .A2(n545), .ZN(n546) );
  XNOR2_X1 U393 ( .A(G140), .B(KEYINPUT10), .ZN(n400) );
  XOR2_X1 U394 ( .A(KEYINPUT71), .B(G131), .Z(n464) );
  XNOR2_X1 U395 ( .A(n439), .B(n403), .ZN(n440) );
  XNOR2_X1 U396 ( .A(G113), .B(G143), .ZN(n437) );
  INV_X1 U397 ( .A(n493), .ZN(n360) );
  XNOR2_X1 U398 ( .A(n399), .B(n525), .ZN(n667) );
  INV_X1 U399 ( .A(n346), .ZN(n381) );
  INV_X1 U400 ( .A(n657), .ZN(n380) );
  NAND2_X1 U401 ( .A1(n616), .A2(n390), .ZN(n382) );
  OR2_X1 U402 ( .A1(n616), .A2(n393), .ZN(n392) );
  INV_X1 U403 ( .A(KEYINPUT30), .ZN(n373) );
  XNOR2_X1 U404 ( .A(n499), .B(KEYINPUT25), .ZN(n401) );
  OR2_X2 U405 ( .A1(n707), .A2(G902), .ZN(n402) );
  XNOR2_X1 U406 ( .A(n376), .B(G113), .ZN(n467) );
  XNOR2_X1 U407 ( .A(KEYINPUT3), .B(G119), .ZN(n376) );
  XOR2_X1 U408 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n453) );
  INV_X1 U409 ( .A(G134), .ZN(n444) );
  XOR2_X1 U410 ( .A(KEYINPUT101), .B(KEYINPUT103), .Z(n447) );
  INV_X1 U411 ( .A(n658), .ZN(n582) );
  NAND2_X1 U412 ( .A1(n365), .A2(n364), .ZN(n502) );
  NAND2_X1 U413 ( .A1(n345), .A2(n367), .ZN(n364) );
  BUF_X1 U414 ( .A(n697), .Z(n706) );
  XNOR2_X1 U415 ( .A(n483), .B(n482), .ZN(n485) );
  XNOR2_X1 U416 ( .A(n388), .B(n386), .ZN(n483) );
  AND2_X1 U417 ( .A1(n606), .A2(G953), .ZN(n710) );
  INV_X1 U418 ( .A(KEYINPUT83), .ZN(n655) );
  XOR2_X1 U419 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n438) );
  INV_X1 U420 ( .A(n405), .ZN(n407) );
  XNOR2_X1 U421 ( .A(KEYINPUT81), .B(KEYINPUT18), .ZN(n405) );
  OR2_X1 U422 ( .A1(n660), .A2(n522), .ZN(n463) );
  NOR2_X1 U423 ( .A1(n589), .A2(n588), .ZN(n591) );
  XNOR2_X1 U424 ( .A(KEYINPUT7), .B(KEYINPUT102), .ZN(n446) );
  NAND2_X1 U425 ( .A1(n658), .A2(n657), .ZN(n663) );
  NOR2_X1 U426 ( .A1(n523), .A2(n522), .ZN(n353) );
  XNOR2_X1 U427 ( .A(n377), .B(n467), .ZN(n473) );
  INV_X1 U428 ( .A(G110), .ZN(n415) );
  XNOR2_X1 U429 ( .A(n487), .B(n404), .ZN(n491) );
  XNOR2_X1 U430 ( .A(KEYINPUT99), .B(KEYINPUT74), .ZN(n404) );
  XNOR2_X1 U431 ( .A(G128), .B(G110), .ZN(n486) );
  XNOR2_X1 U432 ( .A(G119), .B(KEYINPUT24), .ZN(n488) );
  XOR2_X1 U433 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n489) );
  XNOR2_X1 U434 ( .A(n359), .B(n441), .ZN(n603) );
  XNOR2_X1 U435 ( .A(n440), .B(n360), .ZN(n359) );
  XNOR2_X1 U436 ( .A(n492), .B(n480), .ZN(n388) );
  XNOR2_X1 U437 ( .A(n479), .B(n387), .ZN(n386) );
  XNOR2_X1 U438 ( .A(G140), .B(G107), .ZN(n479) );
  XNOR2_X1 U439 ( .A(KEYINPUT80), .B(KEYINPUT96), .ZN(n387) );
  NOR2_X1 U440 ( .A1(n598), .A2(KEYINPUT79), .ZN(n597) );
  NOR2_X1 U441 ( .A1(n381), .A2(n380), .ZN(n379) );
  NOR2_X1 U442 ( .A1(n559), .A2(n511), .ZN(n549) );
  AND2_X1 U443 ( .A1(n555), .A2(n375), .ZN(n374) );
  XNOR2_X1 U444 ( .A(n553), .B(n373), .ZN(n372) );
  INV_X1 U445 ( .A(n554), .ZN(n375) );
  OR2_X1 U446 ( .A1(n541), .A2(n542), .ZN(n579) );
  XNOR2_X1 U447 ( .A(KEYINPUT76), .B(KEYINPUT77), .ZN(n418) );
  XNOR2_X1 U448 ( .A(n451), .B(n356), .ZN(n456) );
  NOR2_X1 U449 ( .A1(n670), .A2(n513), .ZN(n514) );
  OR2_X1 U450 ( .A1(n688), .A2(n584), .ZN(n585) );
  NAND2_X1 U451 ( .A1(n363), .A2(n362), .ZN(n520) );
  INV_X1 U452 ( .A(KEYINPUT105), .ZN(n354) );
  NAND2_X1 U453 ( .A1(n502), .A2(n350), .ZN(n355) );
  XNOR2_X1 U454 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U455 ( .A1(n695), .A2(G953), .ZN(n696) );
  AND2_X1 U456 ( .A1(n368), .A2(n478), .ZN(n345) );
  NAND2_X1 U457 ( .A1(n425), .A2(n391), .ZN(n346) );
  XOR2_X1 U458 ( .A(KEYINPUT73), .B(G469), .Z(n347) );
  AND2_X1 U459 ( .A1(n382), .A2(n379), .ZN(n348) );
  AND2_X1 U460 ( .A1(n670), .A2(n524), .ZN(n349) );
  NAND2_X1 U461 ( .A1(n374), .A2(n372), .ZN(n577) );
  AND2_X1 U462 ( .A1(n500), .A2(n674), .ZN(n350) );
  XNOR2_X1 U463 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n351) );
  INV_X1 U464 ( .A(n599), .ZN(n391) );
  XNOR2_X1 U465 ( .A(KEYINPUT84), .B(KEYINPUT45), .ZN(n352) );
  XNOR2_X2 U466 ( .A(n353), .B(KEYINPUT68), .ZN(n669) );
  NAND2_X1 U467 ( .A1(n532), .A2(n378), .ZN(n394) );
  INV_X1 U468 ( .A(n465), .ZN(n356) );
  NOR2_X2 U469 ( .A1(n667), .A2(n537), .ZN(n526) );
  XNOR2_X2 U470 ( .A(n357), .B(n597), .ZN(n654) );
  NAND2_X1 U471 ( .A1(n727), .A2(n711), .ZN(n357) );
  XNOR2_X1 U472 ( .A(n358), .B(KEYINPUT87), .ZN(n384) );
  NAND2_X1 U473 ( .A1(n546), .A2(n547), .ZN(n358) );
  OR2_X2 U474 ( .A1(n566), .A2(n434), .ZN(n371) );
  XNOR2_X2 U475 ( .A(n361), .B(n476), .ZN(n673) );
  NAND2_X1 U476 ( .A1(n610), .A2(n475), .ZN(n361) );
  NOR2_X2 U477 ( .A1(n607), .A2(n710), .ZN(n609) );
  NOR2_X1 U478 ( .A1(n735), .A2(n738), .ZN(n587) );
  NAND2_X1 U479 ( .A1(n367), .A2(n368), .ZN(n362) );
  INV_X1 U480 ( .A(n366), .ZN(n363) );
  NAND2_X1 U481 ( .A1(n366), .A2(n478), .ZN(n365) );
  INV_X1 U482 ( .A(n539), .ZN(n367) );
  NAND2_X1 U483 ( .A1(n463), .A2(n351), .ZN(n369) );
  NAND2_X1 U484 ( .A1(n537), .A2(n351), .ZN(n370) );
  XNOR2_X2 U485 ( .A(n371), .B(KEYINPUT0), .ZN(n537) );
  NOR2_X2 U486 ( .A1(n577), .A2(n582), .ZN(n578) );
  INV_X1 U487 ( .A(n737), .ZN(n378) );
  AND2_X1 U488 ( .A1(n382), .A2(n346), .ZN(n389) );
  XNOR2_X2 U489 ( .A(n421), .B(n719), .ZN(n616) );
  XNOR2_X1 U490 ( .A(n383), .B(n352), .ZN(n711) );
  AND2_X2 U491 ( .A1(n596), .A2(n595), .ZN(n727) );
  NAND2_X1 U492 ( .A1(n398), .A2(n384), .ZN(n383) );
  XNOR2_X2 U493 ( .A(n564), .B(KEYINPUT1), .ZN(n670) );
  XNOR2_X2 U494 ( .A(n385), .B(n347), .ZN(n564) );
  NAND2_X1 U495 ( .A1(n389), .A2(n392), .ZN(n516) );
  NOR2_X1 U496 ( .A1(n425), .A2(n391), .ZN(n390) );
  INV_X1 U497 ( .A(n425), .ZN(n393) );
  NAND2_X1 U498 ( .A1(n532), .A2(KEYINPUT44), .ZN(n395) );
  NAND2_X1 U499 ( .A1(n394), .A2(n397), .ZN(n396) );
  NAND2_X1 U500 ( .A1(n396), .A2(n395), .ZN(n398) );
  INV_X1 U501 ( .A(KEYINPUT44), .ZN(n397) );
  NAND2_X1 U502 ( .A1(n669), .A2(n349), .ZN(n399) );
  AND2_X1 U503 ( .A1(n669), .A2(n670), .ZN(n535) );
  XNOR2_X1 U504 ( .A(n435), .B(n400), .ZN(n493) );
  XNOR2_X2 U505 ( .A(G146), .B(G125), .ZN(n435) );
  AND2_X1 U506 ( .A1(G214), .A2(n469), .ZN(n403) );
  INV_X1 U507 ( .A(KEYINPUT46), .ZN(n586) );
  XNOR2_X1 U508 ( .A(KEYINPUT28), .B(KEYINPUT111), .ZN(n562) );
  XNOR2_X1 U509 ( .A(KEYINPUT48), .B(KEYINPUT86), .ZN(n590) );
  INV_X1 U510 ( .A(n481), .ZN(n482) );
  XNOR2_X1 U511 ( .A(n563), .B(n562), .ZN(n565) );
  XNOR2_X1 U512 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U513 ( .A(KEYINPUT17), .B(KEYINPUT91), .ZN(n406) );
  XNOR2_X1 U514 ( .A(n407), .B(n406), .ZN(n409) );
  XNOR2_X1 U515 ( .A(n435), .B(KEYINPUT92), .ZN(n408) );
  XNOR2_X1 U516 ( .A(n408), .B(n409), .ZN(n413) );
  XNOR2_X2 U517 ( .A(n410), .B(G128), .ZN(n445) );
  NAND2_X1 U518 ( .A1(G224), .A2(n728), .ZN(n411) );
  XNOR2_X1 U519 ( .A(n445), .B(n411), .ZN(n412) );
  XNOR2_X1 U520 ( .A(n413), .B(n412), .ZN(n416) );
  XNOR2_X1 U521 ( .A(n414), .B(KEYINPUT4), .ZN(n471) );
  XNOR2_X1 U522 ( .A(n415), .B(G104), .ZN(n717) );
  XNOR2_X1 U523 ( .A(n471), .B(n717), .ZN(n481) );
  XNOR2_X1 U524 ( .A(n416), .B(n481), .ZN(n421) );
  XNOR2_X1 U525 ( .A(n417), .B(G107), .ZN(n449) );
  XNOR2_X1 U526 ( .A(n418), .B(KEYINPUT16), .ZN(n419) );
  XNOR2_X1 U527 ( .A(n449), .B(n419), .ZN(n420) );
  XNOR2_X1 U528 ( .A(n420), .B(n467), .ZN(n719) );
  XNOR2_X1 U529 ( .A(KEYINPUT15), .B(G902), .ZN(n599) );
  INV_X1 U530 ( .A(G902), .ZN(n475) );
  INV_X1 U531 ( .A(G237), .ZN(n422) );
  NAND2_X1 U532 ( .A1(n475), .A2(n422), .ZN(n426) );
  NAND2_X1 U533 ( .A1(n426), .A2(G210), .ZN(n424) );
  INV_X1 U534 ( .A(KEYINPUT93), .ZN(n423) );
  XNOR2_X1 U535 ( .A(n424), .B(n423), .ZN(n425) );
  NAND2_X1 U536 ( .A1(n426), .A2(G214), .ZN(n657) );
  XNOR2_X1 U537 ( .A(KEYINPUT66), .B(KEYINPUT19), .ZN(n428) );
  XNOR2_X1 U538 ( .A(n548), .B(n428), .ZN(n566) );
  NAND2_X1 U539 ( .A1(G234), .A2(G237), .ZN(n429) );
  XNOR2_X1 U540 ( .A(KEYINPUT14), .B(n429), .ZN(n431) );
  NAND2_X1 U541 ( .A1(G952), .A2(n431), .ZN(n687) );
  NOR2_X1 U542 ( .A1(G953), .A2(n687), .ZN(n508) );
  NOR2_X1 U543 ( .A1(G898), .A2(n728), .ZN(n430) );
  XOR2_X1 U544 ( .A(KEYINPUT94), .B(n430), .Z(n720) );
  NAND2_X1 U545 ( .A1(G902), .A2(n431), .ZN(n506) );
  NOR2_X1 U546 ( .A1(n720), .A2(n506), .ZN(n432) );
  OR2_X1 U547 ( .A1(n508), .A2(n432), .ZN(n433) );
  XNOR2_X1 U548 ( .A(n433), .B(KEYINPUT95), .ZN(n434) );
  XNOR2_X1 U549 ( .A(n464), .B(G104), .ZN(n436) );
  XNOR2_X1 U550 ( .A(n436), .B(G122), .ZN(n441) );
  XNOR2_X1 U551 ( .A(n438), .B(n437), .ZN(n439) );
  NOR2_X1 U552 ( .A1(G953), .A2(G237), .ZN(n469) );
  NOR2_X1 U553 ( .A1(G902), .A2(n603), .ZN(n443) );
  XNOR2_X1 U554 ( .A(KEYINPUT13), .B(G475), .ZN(n442) );
  XOR2_X1 U555 ( .A(n443), .B(n442), .Z(n541) );
  INV_X1 U556 ( .A(n541), .ZN(n527) );
  XNOR2_X2 U557 ( .A(n445), .B(n444), .ZN(n465) );
  XNOR2_X1 U558 ( .A(n446), .B(KEYINPUT9), .ZN(n448) );
  XNOR2_X1 U559 ( .A(n448), .B(n447), .ZN(n450) );
  XNOR2_X1 U560 ( .A(n450), .B(n449), .ZN(n451) );
  NAND2_X1 U561 ( .A1(G234), .A2(n728), .ZN(n452) );
  XNOR2_X1 U562 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U563 ( .A(KEYINPUT70), .B(n454), .Z(n495) );
  NAND2_X1 U564 ( .A1(G217), .A2(n495), .ZN(n455) );
  XNOR2_X1 U565 ( .A(n456), .B(n455), .ZN(n703) );
  NOR2_X1 U566 ( .A1(n703), .A2(G902), .ZN(n457) );
  XOR2_X1 U567 ( .A(n457), .B(G478), .Z(n542) );
  NOR2_X1 U568 ( .A1(n527), .A2(n542), .ZN(n459) );
  INV_X1 U569 ( .A(KEYINPUT104), .ZN(n458) );
  XNOR2_X1 U570 ( .A(n459), .B(n458), .ZN(n660) );
  NAND2_X1 U571 ( .A1(G234), .A2(n599), .ZN(n460) );
  XNOR2_X1 U572 ( .A(KEYINPUT20), .B(n460), .ZN(n498) );
  NAND2_X1 U573 ( .A1(n498), .A2(G221), .ZN(n462) );
  INV_X1 U574 ( .A(KEYINPUT21), .ZN(n461) );
  XNOR2_X1 U575 ( .A(n462), .B(n461), .ZN(n675) );
  INV_X1 U576 ( .A(n675), .ZN(n522) );
  XOR2_X1 U577 ( .A(KEYINPUT5), .B(G116), .Z(n468) );
  NAND2_X1 U578 ( .A1(n469), .A2(G210), .ZN(n470) );
  XNOR2_X1 U579 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U580 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U581 ( .A(n484), .B(n474), .ZN(n610) );
  XOR2_X1 U582 ( .A(G472), .B(KEYINPUT75), .Z(n476) );
  INV_X1 U583 ( .A(KEYINPUT6), .ZN(n477) );
  INV_X1 U584 ( .A(n524), .ZN(n478) );
  NAND2_X1 U585 ( .A1(G227), .A2(n728), .ZN(n480) );
  INV_X1 U586 ( .A(n670), .ZN(n500) );
  XNOR2_X1 U587 ( .A(n486), .B(KEYINPUT23), .ZN(n487) );
  XNOR2_X1 U588 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U589 ( .A(n491), .B(n490), .ZN(n494) );
  XNOR2_X1 U590 ( .A(n493), .B(n492), .ZN(n724) );
  XNOR2_X1 U591 ( .A(n724), .B(n494), .ZN(n497) );
  NAND2_X1 U592 ( .A1(G221), .A2(n495), .ZN(n496) );
  XNOR2_X1 U593 ( .A(n497), .B(n496), .ZN(n707) );
  NAND2_X1 U594 ( .A1(G217), .A2(n498), .ZN(n499) );
  INV_X1 U595 ( .A(n523), .ZN(n674) );
  XNOR2_X1 U596 ( .A(n544), .B(G101), .ZN(G3) );
  AND2_X1 U597 ( .A1(n670), .A2(n523), .ZN(n501) );
  NAND2_X1 U598 ( .A1(n502), .A2(n501), .ZN(n505) );
  INV_X1 U599 ( .A(KEYINPUT64), .ZN(n503) );
  XNOR2_X1 U600 ( .A(n503), .B(KEYINPUT32), .ZN(n504) );
  XOR2_X1 U601 ( .A(n521), .B(G119), .Z(G21) );
  OR2_X1 U602 ( .A1(n728), .A2(n506), .ZN(n507) );
  NOR2_X1 U603 ( .A1(G900), .A2(n507), .ZN(n509) );
  NOR2_X1 U604 ( .A1(n509), .A2(n508), .ZN(n554) );
  NOR2_X1 U605 ( .A1(n554), .A2(n522), .ZN(n510) );
  NAND2_X1 U606 ( .A1(n523), .A2(n510), .ZN(n559) );
  XNOR2_X1 U607 ( .A(KEYINPUT108), .B(n579), .ZN(n643) );
  INV_X1 U608 ( .A(n643), .ZN(n641) );
  NAND2_X1 U609 ( .A1(n524), .A2(n641), .ZN(n511) );
  NAND2_X1 U610 ( .A1(n549), .A2(n657), .ZN(n512) );
  XOR2_X1 U611 ( .A(KEYINPUT109), .B(n512), .Z(n513) );
  XNOR2_X1 U612 ( .A(n514), .B(KEYINPUT110), .ZN(n515) );
  XNOR2_X1 U613 ( .A(n515), .B(KEYINPUT43), .ZN(n517) );
  INV_X1 U614 ( .A(n516), .ZN(n556) );
  NOR2_X1 U615 ( .A1(n517), .A2(n556), .ZN(n594) );
  XOR2_X1 U616 ( .A(n594), .B(G140), .Z(G42) );
  XNOR2_X1 U617 ( .A(n673), .B(KEYINPUT106), .ZN(n561) );
  OR2_X1 U618 ( .A1(n670), .A2(n674), .ZN(n518) );
  NOR2_X1 U619 ( .A1(n561), .A2(n518), .ZN(n519) );
  AND2_X1 U620 ( .A1(n520), .A2(n519), .ZN(n634) );
  INV_X1 U621 ( .A(KEYINPUT33), .ZN(n525) );
  XNOR2_X1 U622 ( .A(n526), .B(KEYINPUT34), .ZN(n529) );
  NAND2_X1 U623 ( .A1(n527), .A2(n542), .ZN(n528) );
  XNOR2_X1 U624 ( .A(KEYINPUT107), .B(n528), .ZN(n557) );
  NAND2_X1 U625 ( .A1(n529), .A2(n557), .ZN(n531) );
  XNOR2_X1 U626 ( .A(KEYINPUT35), .B(KEYINPUT82), .ZN(n530) );
  BUF_X1 U627 ( .A(n533), .Z(n737) );
  NAND2_X1 U628 ( .A1(n533), .A2(KEYINPUT44), .ZN(n534) );
  XNOR2_X1 U629 ( .A(n534), .B(KEYINPUT88), .ZN(n547) );
  NAND2_X1 U630 ( .A1(n535), .A2(n673), .ZN(n536) );
  XNOR2_X1 U631 ( .A(n536), .B(KEYINPUT100), .ZN(n680) );
  NOR2_X1 U632 ( .A1(n680), .A2(n539), .ZN(n538) );
  XNOR2_X1 U633 ( .A(n538), .B(KEYINPUT31), .ZN(n645) );
  NAND2_X1 U634 ( .A1(n669), .A2(n564), .ZN(n552) );
  NOR2_X1 U635 ( .A1(n552), .A2(n673), .ZN(n540) );
  NAND2_X1 U636 ( .A1(n367), .A2(n540), .ZN(n629) );
  NAND2_X1 U637 ( .A1(n645), .A2(n629), .ZN(n543) );
  NAND2_X1 U638 ( .A1(n542), .A2(n541), .ZN(n646) );
  NAND2_X1 U639 ( .A1(n579), .A2(n646), .ZN(n662) );
  NAND2_X1 U640 ( .A1(n543), .A2(n662), .ZN(n545) );
  NAND2_X1 U641 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U642 ( .A(KEYINPUT36), .B(n550), .Z(n551) );
  NAND2_X1 U643 ( .A1(n551), .A2(n670), .ZN(n650) );
  INV_X1 U644 ( .A(n552), .ZN(n555) );
  NAND2_X1 U645 ( .A1(n657), .A2(n561), .ZN(n553) );
  NAND2_X1 U646 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U647 ( .A1(n577), .A2(n558), .ZN(n640) );
  INV_X1 U648 ( .A(n559), .ZN(n560) );
  NAND2_X1 U649 ( .A1(n561), .A2(n560), .ZN(n563) );
  NAND2_X1 U650 ( .A1(n565), .A2(n564), .ZN(n584) );
  BUF_X1 U651 ( .A(n566), .Z(n567) );
  NOR2_X1 U652 ( .A1(n584), .A2(n567), .ZN(n635) );
  AND2_X1 U653 ( .A1(n635), .A2(n662), .ZN(n569) );
  INV_X1 U654 ( .A(KEYINPUT47), .ZN(n568) );
  XNOR2_X1 U655 ( .A(n569), .B(n568), .ZN(n570) );
  NOR2_X1 U656 ( .A1(n640), .A2(n570), .ZN(n571) );
  NAND2_X1 U657 ( .A1(n571), .A2(KEYINPUT78), .ZN(n575) );
  INV_X1 U658 ( .A(n571), .ZN(n573) );
  INV_X1 U659 ( .A(KEYINPUT78), .ZN(n572) );
  NAND2_X1 U660 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U661 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U662 ( .A1(n650), .A2(n576), .ZN(n589) );
  XNOR2_X1 U663 ( .A(n578), .B(KEYINPUT39), .ZN(n592) );
  NOR2_X1 U664 ( .A1(n579), .A2(n592), .ZN(n581) );
  XNOR2_X1 U665 ( .A(KEYINPUT40), .B(KEYINPUT112), .ZN(n580) );
  XNOR2_X1 U666 ( .A(n581), .B(n580), .ZN(n735) );
  NOR2_X1 U667 ( .A1(n660), .A2(n663), .ZN(n583) );
  XNOR2_X1 U668 ( .A(KEYINPUT41), .B(n583), .ZN(n688) );
  XOR2_X1 U669 ( .A(KEYINPUT42), .B(n585), .Z(n738) );
  XNOR2_X1 U670 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U671 ( .A(n591), .B(n590), .ZN(n596) );
  OR2_X1 U672 ( .A1(n646), .A2(n592), .ZN(n651) );
  INV_X1 U673 ( .A(n651), .ZN(n593) );
  NOR2_X1 U674 ( .A1(n594), .A2(n593), .ZN(n595) );
  INV_X1 U675 ( .A(KEYINPUT2), .ZN(n598) );
  NAND2_X1 U676 ( .A1(n598), .A2(KEYINPUT79), .ZN(n653) );
  AND2_X1 U677 ( .A1(n653), .A2(n391), .ZN(n600) );
  AND2_X2 U678 ( .A1(n654), .A2(n600), .ZN(n697) );
  AND2_X2 U679 ( .A1(n697), .A2(G475), .ZN(n605) );
  XNOR2_X1 U680 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n601) );
  XNOR2_X1 U681 ( .A(n601), .B(KEYINPUT59), .ZN(n602) );
  XOR2_X1 U682 ( .A(n603), .B(n602), .Z(n604) );
  XNOR2_X1 U683 ( .A(n605), .B(n604), .ZN(n607) );
  INV_X1 U684 ( .A(G952), .ZN(n606) );
  XOR2_X1 U685 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n608) );
  XNOR2_X1 U686 ( .A(n609), .B(n608), .ZN(G60) );
  INV_X1 U687 ( .A(KEYINPUT63), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n697), .A2(G472), .ZN(n612) );
  XOR2_X1 U689 ( .A(KEYINPUT62), .B(n610), .Z(n611) );
  XNOR2_X1 U690 ( .A(n612), .B(n611), .ZN(n613) );
  NOR2_X2 U691 ( .A1(n613), .A2(n710), .ZN(n614) );
  XNOR2_X1 U692 ( .A(n615), .B(n614), .ZN(G57) );
  NAND2_X1 U693 ( .A1(n697), .A2(G210), .ZN(n621) );
  XOR2_X1 U694 ( .A(KEYINPUT90), .B(KEYINPUT55), .Z(n618) );
  XNOR2_X1 U695 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n617) );
  XNOR2_X1 U696 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U697 ( .A(n616), .B(n619), .ZN(n620) );
  XNOR2_X1 U698 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U699 ( .A(KEYINPUT122), .B(KEYINPUT56), .ZN(n623) );
  XOR2_X1 U700 ( .A(n623), .B(KEYINPUT85), .Z(n624) );
  XNOR2_X1 U701 ( .A(n625), .B(n624), .ZN(G51) );
  NOR2_X1 U702 ( .A1(n629), .A2(n643), .ZN(n626) );
  XOR2_X1 U703 ( .A(G104), .B(n626), .Z(G6) );
  XOR2_X1 U704 ( .A(KEYINPUT115), .B(KEYINPUT27), .Z(n628) );
  XNOR2_X1 U705 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n627) );
  XNOR2_X1 U706 ( .A(n628), .B(n627), .ZN(n633) );
  NOR2_X1 U707 ( .A1(n629), .A2(n646), .ZN(n631) );
  XNOR2_X1 U708 ( .A(G107), .B(KEYINPUT26), .ZN(n630) );
  XNOR2_X1 U709 ( .A(n631), .B(n630), .ZN(n632) );
  XOR2_X1 U710 ( .A(n633), .B(n632), .Z(G9) );
  XOR2_X1 U711 ( .A(G110), .B(n634), .Z(G12) );
  XOR2_X1 U712 ( .A(KEYINPUT29), .B(KEYINPUT116), .Z(n638) );
  INV_X1 U713 ( .A(n646), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n635), .A2(n636), .ZN(n637) );
  XNOR2_X1 U715 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U716 ( .A(G128), .B(n639), .ZN(G30) );
  XOR2_X1 U717 ( .A(G143), .B(n640), .Z(G45) );
  NAND2_X1 U718 ( .A1(n635), .A2(n641), .ZN(n642) );
  XNOR2_X1 U719 ( .A(n642), .B(G146), .ZN(G48) );
  NOR2_X1 U720 ( .A1(n643), .A2(n645), .ZN(n644) );
  XOR2_X1 U721 ( .A(G113), .B(n644), .Z(G15) );
  NOR2_X1 U722 ( .A1(n646), .A2(n645), .ZN(n648) );
  XNOR2_X1 U723 ( .A(G116), .B(KEYINPUT117), .ZN(n647) );
  XNOR2_X1 U724 ( .A(n648), .B(n647), .ZN(G18) );
  XOR2_X1 U725 ( .A(G125), .B(KEYINPUT37), .Z(n649) );
  XNOR2_X1 U726 ( .A(n650), .B(n649), .ZN(G27) );
  XNOR2_X1 U727 ( .A(G134), .B(KEYINPUT118), .ZN(n652) );
  XNOR2_X1 U728 ( .A(n652), .B(n651), .ZN(G36) );
  NAND2_X1 U729 ( .A1(n654), .A2(n653), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n656), .B(n655), .ZN(n694) );
  NOR2_X1 U731 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U732 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U733 ( .A(KEYINPUT119), .B(n661), .Z(n666) );
  INV_X1 U734 ( .A(n662), .ZN(n664) );
  NOR2_X1 U735 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U736 ( .A1(n666), .A2(n665), .ZN(n668) );
  BUF_X1 U737 ( .A(n667), .Z(n689) );
  NOR2_X1 U738 ( .A1(n668), .A2(n689), .ZN(n684) );
  NOR2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U740 ( .A(n671), .B(KEYINPUT50), .ZN(n672) );
  NOR2_X1 U741 ( .A1(n673), .A2(n672), .ZN(n678) );
  NOR2_X1 U742 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U743 ( .A(n676), .B(KEYINPUT49), .ZN(n677) );
  NAND2_X1 U744 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U745 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U746 ( .A(KEYINPUT51), .B(n681), .ZN(n682) );
  NOR2_X1 U747 ( .A1(n682), .A2(n688), .ZN(n683) );
  NOR2_X1 U748 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U749 ( .A(n685), .B(KEYINPUT52), .ZN(n686) );
  NOR2_X1 U750 ( .A1(n687), .A2(n686), .ZN(n691) );
  NOR2_X1 U751 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U752 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U753 ( .A(n692), .B(KEYINPUT120), .ZN(n693) );
  NAND2_X1 U754 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U755 ( .A(n696), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U756 ( .A1(n706), .A2(G469), .ZN(n701) );
  XOR2_X1 U757 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n698) );
  NOR2_X1 U758 ( .A1(n710), .A2(n702), .ZN(G54) );
  NAND2_X1 U759 ( .A1(n706), .A2(G478), .ZN(n704) );
  XNOR2_X1 U760 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U761 ( .A1(n710), .A2(n705), .ZN(G63) );
  NAND2_X1 U762 ( .A1(n706), .A2(G217), .ZN(n708) );
  XNOR2_X1 U763 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U764 ( .A1(n710), .A2(n709), .ZN(G66) );
  NAND2_X1 U765 ( .A1(n711), .A2(n728), .ZN(n712) );
  XNOR2_X1 U766 ( .A(n712), .B(KEYINPUT126), .ZN(n716) );
  NAND2_X1 U767 ( .A1(G953), .A2(G224), .ZN(n713) );
  XNOR2_X1 U768 ( .A(KEYINPUT61), .B(n713), .ZN(n714) );
  NAND2_X1 U769 ( .A1(n714), .A2(G898), .ZN(n715) );
  NAND2_X1 U770 ( .A1(n716), .A2(n715), .ZN(n723) );
  XOR2_X1 U771 ( .A(G101), .B(n717), .Z(n718) );
  XNOR2_X1 U772 ( .A(n719), .B(n718), .ZN(n721) );
  NAND2_X1 U773 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U774 ( .A(n723), .B(n722), .Z(G69) );
  XOR2_X1 U775 ( .A(KEYINPUT4), .B(n724), .Z(n725) );
  XOR2_X1 U776 ( .A(n726), .B(n725), .Z(n730) );
  XOR2_X1 U777 ( .A(n730), .B(n727), .Z(n729) );
  NAND2_X1 U778 ( .A1(n729), .A2(n728), .ZN(n734) );
  XNOR2_X1 U779 ( .A(G227), .B(n730), .ZN(n731) );
  NAND2_X1 U780 ( .A1(n731), .A2(G900), .ZN(n732) );
  NAND2_X1 U781 ( .A1(G953), .A2(n732), .ZN(n733) );
  NAND2_X1 U782 ( .A1(n734), .A2(n733), .ZN(G72) );
  XNOR2_X1 U783 ( .A(n735), .B(G131), .ZN(n736) );
  XNOR2_X1 U784 ( .A(n736), .B(KEYINPUT127), .ZN(G33) );
  XOR2_X1 U785 ( .A(n737), .B(G122), .Z(G24) );
  XOR2_X1 U786 ( .A(G137), .B(n738), .Z(G39) );
endmodule

