

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U557 ( .A(KEYINPUT23), .B(KEYINPUT65), .ZN(n523) );
  NOR2_X1 U558 ( .A1(n532), .A2(n531), .ZN(G160) );
  NOR2_X1 U559 ( .A1(n784), .A2(n869), .ZN(n744) );
  XNOR2_X1 U560 ( .A(n750), .B(n749), .ZN(n751) );
  NOR2_X1 U561 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U562 ( .A1(n528), .A2(G2104), .ZN(n903) );
  NOR2_X1 U563 ( .A1(G651), .A2(n651), .ZN(n667) );
  XNOR2_X1 U564 ( .A(n524), .B(n523), .ZN(n527) );
  INV_X1 U565 ( .A(G2105), .ZN(n528) );
  NAND2_X1 U566 ( .A1(G101), .A2(n903), .ZN(n524) );
  NOR2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n525) );
  XOR2_X2 U568 ( .A(KEYINPUT17), .B(n525), .Z(n906) );
  NAND2_X1 U569 ( .A1(G137), .A2(n906), .ZN(n526) );
  NAND2_X1 U570 ( .A1(n527), .A2(n526), .ZN(n532) );
  AND2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n899) );
  NAND2_X1 U572 ( .A1(G113), .A2(n899), .ZN(n530) );
  NOR2_X1 U573 ( .A1(G2104), .A2(n528), .ZN(n897) );
  NAND2_X1 U574 ( .A1(G125), .A2(n897), .ZN(n529) );
  NAND2_X1 U575 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U576 ( .A1(G102), .A2(n903), .ZN(n534) );
  NAND2_X1 U577 ( .A1(G114), .A2(n899), .ZN(n533) );
  NAND2_X1 U578 ( .A1(n534), .A2(n533), .ZN(n539) );
  NAND2_X1 U579 ( .A1(n906), .A2(G138), .ZN(n535) );
  XNOR2_X1 U580 ( .A(n535), .B(KEYINPUT96), .ZN(n537) );
  NAND2_X1 U581 ( .A1(G126), .A2(n897), .ZN(n536) );
  NAND2_X1 U582 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X2 U583 ( .A1(n539), .A2(n538), .ZN(G164) );
  XNOR2_X1 U584 ( .A(G2435), .B(G2446), .ZN(n549) );
  XOR2_X1 U585 ( .A(G2454), .B(G2430), .Z(n541) );
  XNOR2_X1 U586 ( .A(G2451), .B(G2443), .ZN(n540) );
  XNOR2_X1 U587 ( .A(n541), .B(n540), .ZN(n545) );
  XOR2_X1 U588 ( .A(G2427), .B(KEYINPUT113), .Z(n543) );
  XNOR2_X1 U589 ( .A(G1348), .B(G1341), .ZN(n542) );
  XNOR2_X1 U590 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U591 ( .A(n545), .B(n544), .Z(n547) );
  XNOR2_X1 U592 ( .A(KEYINPUT114), .B(G2438), .ZN(n546) );
  XNOR2_X1 U593 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U594 ( .A(n549), .B(n548), .ZN(n550) );
  AND2_X1 U595 ( .A1(n550), .A2(G14), .ZN(G401) );
  AND2_X1 U596 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U597 ( .A(G57), .ZN(G237) );
  INV_X1 U598 ( .A(G132), .ZN(G219) );
  INV_X1 U599 ( .A(G82), .ZN(G220) );
  NOR2_X1 U600 ( .A1(G651), .A2(G543), .ZN(n661) );
  NAND2_X1 U601 ( .A1(n661), .A2(G90), .ZN(n551) );
  XNOR2_X1 U602 ( .A(n551), .B(KEYINPUT68), .ZN(n553) );
  XOR2_X1 U603 ( .A(G543), .B(KEYINPUT0), .Z(n651) );
  INV_X1 U604 ( .A(G651), .ZN(n557) );
  NOR2_X1 U605 ( .A1(n651), .A2(n557), .ZN(n662) );
  NAND2_X1 U606 ( .A1(G77), .A2(n662), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U608 ( .A(n554), .B(KEYINPUT9), .ZN(n556) );
  NAND2_X1 U609 ( .A1(G52), .A2(n667), .ZN(n555) );
  NAND2_X1 U610 ( .A1(n556), .A2(n555), .ZN(n562) );
  NOR2_X1 U611 ( .A1(G543), .A2(n557), .ZN(n558) );
  XOR2_X1 U612 ( .A(KEYINPUT66), .B(n558), .Z(n559) );
  XNOR2_X1 U613 ( .A(KEYINPUT1), .B(n559), .ZN(n660) );
  NAND2_X1 U614 ( .A1(G64), .A2(n660), .ZN(n560) );
  XNOR2_X1 U615 ( .A(KEYINPUT67), .B(n560), .ZN(n561) );
  NOR2_X1 U616 ( .A1(n562), .A2(n561), .ZN(G171) );
  NAND2_X1 U617 ( .A1(n661), .A2(G89), .ZN(n563) );
  XNOR2_X1 U618 ( .A(n563), .B(KEYINPUT4), .ZN(n565) );
  NAND2_X1 U619 ( .A1(G76), .A2(n662), .ZN(n564) );
  NAND2_X1 U620 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U621 ( .A(n566), .B(KEYINPUT5), .ZN(n571) );
  NAND2_X1 U622 ( .A1(n667), .A2(G51), .ZN(n568) );
  NAND2_X1 U623 ( .A1(G63), .A2(n660), .ZN(n567) );
  NAND2_X1 U624 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U625 ( .A(KEYINPUT6), .B(n569), .Z(n570) );
  NAND2_X1 U626 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U627 ( .A(n572), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U628 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U629 ( .A1(G7), .A2(G661), .ZN(n573) );
  XOR2_X1 U630 ( .A(n573), .B(KEYINPUT10), .Z(n928) );
  NAND2_X1 U631 ( .A1(n928), .A2(G567), .ZN(n574) );
  XOR2_X1 U632 ( .A(KEYINPUT11), .B(n574), .Z(G234) );
  NAND2_X1 U633 ( .A1(n660), .A2(G56), .ZN(n575) );
  XOR2_X1 U634 ( .A(KEYINPUT14), .B(n575), .Z(n582) );
  NAND2_X1 U635 ( .A1(G81), .A2(n661), .ZN(n576) );
  XNOR2_X1 U636 ( .A(n576), .B(KEYINPUT72), .ZN(n577) );
  XNOR2_X1 U637 ( .A(n577), .B(KEYINPUT12), .ZN(n579) );
  NAND2_X1 U638 ( .A1(G68), .A2(n662), .ZN(n578) );
  NAND2_X1 U639 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U640 ( .A(KEYINPUT13), .B(n580), .Z(n581) );
  NOR2_X1 U641 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U642 ( .A1(n667), .A2(G43), .ZN(n583) );
  NAND2_X1 U643 ( .A1(n584), .A2(n583), .ZN(n748) );
  INV_X1 U644 ( .A(n748), .ZN(n1027) );
  NAND2_X1 U645 ( .A1(n1027), .A2(G860), .ZN(G153) );
  INV_X1 U646 ( .A(G171), .ZN(G301) );
  NAND2_X1 U647 ( .A1(G54), .A2(n667), .ZN(n591) );
  NAND2_X1 U648 ( .A1(n661), .A2(G92), .ZN(n586) );
  NAND2_X1 U649 ( .A1(G66), .A2(n660), .ZN(n585) );
  NAND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U651 ( .A1(G79), .A2(n662), .ZN(n587) );
  XNOR2_X1 U652 ( .A(KEYINPUT73), .B(n587), .ZN(n588) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U654 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U655 ( .A(n592), .B(KEYINPUT15), .ZN(n593) );
  XNOR2_X1 U656 ( .A(KEYINPUT74), .B(n593), .ZN(n1018) );
  INV_X1 U657 ( .A(G868), .ZN(n678) );
  AND2_X1 U658 ( .A1(n1018), .A2(n678), .ZN(n595) );
  NOR2_X1 U659 ( .A1(n678), .A2(G301), .ZN(n594) );
  NOR2_X1 U660 ( .A1(n595), .A2(n594), .ZN(G284) );
  NAND2_X1 U661 ( .A1(n660), .A2(G65), .ZN(n596) );
  XNOR2_X1 U662 ( .A(n596), .B(KEYINPUT70), .ZN(n603) );
  NAND2_X1 U663 ( .A1(G91), .A2(n661), .ZN(n598) );
  NAND2_X1 U664 ( .A1(G53), .A2(n667), .ZN(n597) );
  NAND2_X1 U665 ( .A1(n598), .A2(n597), .ZN(n601) );
  NAND2_X1 U666 ( .A1(G78), .A2(n662), .ZN(n599) );
  XNOR2_X1 U667 ( .A(KEYINPUT69), .B(n599), .ZN(n600) );
  NOR2_X1 U668 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U669 ( .A1(n603), .A2(n602), .ZN(n1008) );
  XOR2_X1 U670 ( .A(KEYINPUT71), .B(n1008), .Z(G299) );
  NAND2_X1 U671 ( .A1(G286), .A2(G868), .ZN(n605) );
  NAND2_X1 U672 ( .A1(G299), .A2(n678), .ZN(n604) );
  NAND2_X1 U673 ( .A1(n605), .A2(n604), .ZN(G297) );
  INV_X1 U674 ( .A(G559), .ZN(n606) );
  NOR2_X1 U675 ( .A1(G860), .A2(n606), .ZN(n607) );
  XNOR2_X1 U676 ( .A(KEYINPUT75), .B(n607), .ZN(n608) );
  NAND2_X1 U677 ( .A1(n608), .A2(n1018), .ZN(n609) );
  XNOR2_X1 U678 ( .A(n609), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U679 ( .A1(G868), .A2(n748), .ZN(n612) );
  NAND2_X1 U680 ( .A1(n1018), .A2(G868), .ZN(n610) );
  NOR2_X1 U681 ( .A1(G559), .A2(n610), .ZN(n611) );
  NOR2_X1 U682 ( .A1(n612), .A2(n611), .ZN(G282) );
  NAND2_X1 U683 ( .A1(G99), .A2(n903), .ZN(n614) );
  NAND2_X1 U684 ( .A1(G111), .A2(n899), .ZN(n613) );
  NAND2_X1 U685 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U686 ( .A(n615), .B(KEYINPUT77), .ZN(n617) );
  NAND2_X1 U687 ( .A1(G135), .A2(n906), .ZN(n616) );
  NAND2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n621) );
  XOR2_X1 U689 ( .A(KEYINPUT76), .B(KEYINPUT18), .Z(n619) );
  NAND2_X1 U690 ( .A1(G123), .A2(n897), .ZN(n618) );
  XNOR2_X1 U691 ( .A(n619), .B(n618), .ZN(n620) );
  NOR2_X1 U692 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U693 ( .A(n622), .B(KEYINPUT78), .ZN(n978) );
  XOR2_X1 U694 ( .A(G2096), .B(KEYINPUT79), .Z(n623) );
  XNOR2_X1 U695 ( .A(n978), .B(n623), .ZN(n624) );
  INV_X1 U696 ( .A(G2100), .ZN(n854) );
  NAND2_X1 U697 ( .A1(n624), .A2(n854), .ZN(G156) );
  NAND2_X1 U698 ( .A1(G93), .A2(n661), .ZN(n625) );
  XNOR2_X1 U699 ( .A(n625), .B(KEYINPUT80), .ZN(n633) );
  NAND2_X1 U700 ( .A1(G55), .A2(n667), .ZN(n626) );
  XNOR2_X1 U701 ( .A(n626), .B(KEYINPUT82), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n662), .A2(G80), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U704 ( .A1(G67), .A2(n660), .ZN(n629) );
  XNOR2_X1 U705 ( .A(KEYINPUT81), .B(n629), .ZN(n630) );
  NOR2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n679) );
  NAND2_X1 U708 ( .A1(n1018), .A2(G559), .ZN(n634) );
  XOR2_X1 U709 ( .A(n1027), .B(n634), .Z(n676) );
  NOR2_X1 U710 ( .A1(n676), .A2(G860), .ZN(n635) );
  XNOR2_X1 U711 ( .A(n635), .B(KEYINPUT83), .ZN(n636) );
  XNOR2_X1 U712 ( .A(n679), .B(n636), .ZN(G145) );
  NAND2_X1 U713 ( .A1(G86), .A2(n661), .ZN(n637) );
  XNOR2_X1 U714 ( .A(n637), .B(KEYINPUT86), .ZN(n646) );
  NAND2_X1 U715 ( .A1(G73), .A2(n662), .ZN(n638) );
  XOR2_X1 U716 ( .A(KEYINPUT87), .B(n638), .Z(n639) );
  XNOR2_X1 U717 ( .A(n639), .B(KEYINPUT2), .ZN(n641) );
  NAND2_X1 U718 ( .A1(G48), .A2(n667), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U720 ( .A1(G61), .A2(n660), .ZN(n642) );
  XNOR2_X1 U721 ( .A(KEYINPUT85), .B(n642), .ZN(n643) );
  NOR2_X1 U722 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U723 ( .A1(n646), .A2(n645), .ZN(G305) );
  NAND2_X1 U724 ( .A1(G49), .A2(n667), .ZN(n648) );
  NAND2_X1 U725 ( .A1(G74), .A2(G651), .ZN(n647) );
  NAND2_X1 U726 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U727 ( .A(KEYINPUT84), .B(n649), .ZN(n650) );
  NOR2_X1 U728 ( .A1(n660), .A2(n650), .ZN(n653) );
  NAND2_X1 U729 ( .A1(n651), .A2(G87), .ZN(n652) );
  NAND2_X1 U730 ( .A1(n653), .A2(n652), .ZN(G288) );
  NAND2_X1 U731 ( .A1(G88), .A2(n661), .ZN(n655) );
  NAND2_X1 U732 ( .A1(G75), .A2(n662), .ZN(n654) );
  NAND2_X1 U733 ( .A1(n655), .A2(n654), .ZN(n659) );
  NAND2_X1 U734 ( .A1(n667), .A2(G50), .ZN(n657) );
  NAND2_X1 U735 ( .A1(G62), .A2(n660), .ZN(n656) );
  NAND2_X1 U736 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U737 ( .A1(n659), .A2(n658), .ZN(G166) );
  INV_X1 U738 ( .A(G166), .ZN(G303) );
  AND2_X1 U739 ( .A1(G60), .A2(n660), .ZN(n666) );
  NAND2_X1 U740 ( .A1(G85), .A2(n661), .ZN(n664) );
  NAND2_X1 U741 ( .A1(G72), .A2(n662), .ZN(n663) );
  NAND2_X1 U742 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U743 ( .A1(n666), .A2(n665), .ZN(n669) );
  NAND2_X1 U744 ( .A1(n667), .A2(G47), .ZN(n668) );
  NAND2_X1 U745 ( .A1(n669), .A2(n668), .ZN(G290) );
  XOR2_X1 U746 ( .A(G288), .B(G299), .Z(n670) );
  XNOR2_X1 U747 ( .A(n679), .B(n670), .ZN(n671) );
  XOR2_X1 U748 ( .A(n671), .B(KEYINPUT88), .Z(n673) );
  XOR2_X1 U749 ( .A(G303), .B(KEYINPUT19), .Z(n672) );
  XNOR2_X1 U750 ( .A(n673), .B(n672), .ZN(n674) );
  XOR2_X1 U751 ( .A(n674), .B(G290), .Z(n675) );
  XNOR2_X1 U752 ( .A(G305), .B(n675), .ZN(n916) );
  XOR2_X1 U753 ( .A(n676), .B(n916), .Z(n677) );
  NOR2_X1 U754 ( .A1(n678), .A2(n677), .ZN(n681) );
  NOR2_X1 U755 ( .A1(G868), .A2(n679), .ZN(n680) );
  NOR2_X1 U756 ( .A1(n681), .A2(n680), .ZN(G295) );
  NAND2_X1 U757 ( .A1(G2078), .A2(G2084), .ZN(n682) );
  XNOR2_X1 U758 ( .A(n682), .B(KEYINPUT20), .ZN(n683) );
  XNOR2_X1 U759 ( .A(n683), .B(KEYINPUT89), .ZN(n684) );
  NAND2_X1 U760 ( .A1(n684), .A2(G2090), .ZN(n685) );
  XNOR2_X1 U761 ( .A(n685), .B(KEYINPUT21), .ZN(n686) );
  XNOR2_X1 U762 ( .A(n686), .B(KEYINPUT90), .ZN(n687) );
  NAND2_X1 U763 ( .A1(n687), .A2(G2072), .ZN(n688) );
  XOR2_X1 U764 ( .A(KEYINPUT91), .B(n688), .Z(G158) );
  XNOR2_X1 U765 ( .A(KEYINPUT92), .B(G44), .ZN(n689) );
  XNOR2_X1 U766 ( .A(n689), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U767 ( .A1(G220), .A2(G219), .ZN(n690) );
  XNOR2_X1 U768 ( .A(KEYINPUT22), .B(n690), .ZN(n691) );
  NAND2_X1 U769 ( .A1(n691), .A2(G96), .ZN(n692) );
  NOR2_X1 U770 ( .A1(n692), .A2(G218), .ZN(n693) );
  XNOR2_X1 U771 ( .A(n693), .B(KEYINPUT93), .ZN(n853) );
  NAND2_X1 U772 ( .A1(G2106), .A2(n853), .ZN(n697) );
  NAND2_X1 U773 ( .A1(G69), .A2(G120), .ZN(n694) );
  NOR2_X1 U774 ( .A1(G237), .A2(n694), .ZN(n695) );
  NAND2_X1 U775 ( .A1(G108), .A2(n695), .ZN(n852) );
  NAND2_X1 U776 ( .A1(G567), .A2(n852), .ZN(n696) );
  NAND2_X1 U777 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U778 ( .A(KEYINPUT94), .B(n698), .ZN(n927) );
  NAND2_X1 U779 ( .A1(G661), .A2(G483), .ZN(n699) );
  XOR2_X1 U780 ( .A(KEYINPUT95), .B(n699), .Z(n700) );
  NOR2_X1 U781 ( .A1(n927), .A2(n700), .ZN(n851) );
  NAND2_X1 U782 ( .A1(n851), .A2(G36), .ZN(G176) );
  NAND2_X1 U783 ( .A1(G40), .A2(G160), .ZN(n701) );
  XNOR2_X1 U784 ( .A(KEYINPUT97), .B(n701), .ZN(n737) );
  NOR2_X1 U785 ( .A1(G1384), .A2(G164), .ZN(n702) );
  XNOR2_X1 U786 ( .A(n702), .B(KEYINPUT64), .ZN(n736) );
  INV_X1 U787 ( .A(n736), .ZN(n703) );
  NAND2_X1 U788 ( .A1(n737), .A2(n703), .ZN(n734) );
  INV_X1 U789 ( .A(n734), .ZN(n844) );
  INV_X1 U790 ( .A(G2067), .ZN(n857) );
  XOR2_X1 U791 ( .A(n857), .B(KEYINPUT37), .Z(n841) );
  NAND2_X1 U792 ( .A1(n906), .A2(G140), .ZN(n704) );
  XNOR2_X1 U793 ( .A(n704), .B(KEYINPUT98), .ZN(n706) );
  NAND2_X1 U794 ( .A1(G104), .A2(n903), .ZN(n705) );
  NAND2_X1 U795 ( .A1(n706), .A2(n705), .ZN(n708) );
  XOR2_X1 U796 ( .A(KEYINPUT34), .B(KEYINPUT99), .Z(n707) );
  XNOR2_X1 U797 ( .A(n708), .B(n707), .ZN(n713) );
  NAND2_X1 U798 ( .A1(G116), .A2(n899), .ZN(n710) );
  NAND2_X1 U799 ( .A1(G128), .A2(n897), .ZN(n709) );
  NAND2_X1 U800 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U801 ( .A(KEYINPUT35), .B(n711), .Z(n712) );
  NOR2_X1 U802 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U803 ( .A(KEYINPUT36), .B(n714), .ZN(n910) );
  NOR2_X1 U804 ( .A1(n841), .A2(n910), .ZN(n998) );
  NAND2_X1 U805 ( .A1(n844), .A2(n998), .ZN(n839) );
  NAND2_X1 U806 ( .A1(n899), .A2(G107), .ZN(n715) );
  XNOR2_X1 U807 ( .A(n715), .B(KEYINPUT100), .ZN(n717) );
  NAND2_X1 U808 ( .A1(G119), .A2(n897), .ZN(n716) );
  NAND2_X1 U809 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U810 ( .A(n718), .B(KEYINPUT101), .ZN(n720) );
  NAND2_X1 U811 ( .A1(G95), .A2(n903), .ZN(n719) );
  NAND2_X1 U812 ( .A1(n720), .A2(n719), .ZN(n723) );
  NAND2_X1 U813 ( .A1(n906), .A2(G131), .ZN(n721) );
  XOR2_X1 U814 ( .A(KEYINPUT102), .B(n721), .Z(n722) );
  OR2_X1 U815 ( .A1(n723), .A2(n722), .ZN(n889) );
  AND2_X1 U816 ( .A1(n889), .A2(G1991), .ZN(n733) );
  NAND2_X1 U817 ( .A1(G117), .A2(n899), .ZN(n725) );
  NAND2_X1 U818 ( .A1(G141), .A2(n906), .ZN(n724) );
  NAND2_X1 U819 ( .A1(n725), .A2(n724), .ZN(n729) );
  NAND2_X1 U820 ( .A1(G105), .A2(n903), .ZN(n726) );
  XNOR2_X1 U821 ( .A(n726), .B(KEYINPUT103), .ZN(n727) );
  XNOR2_X1 U822 ( .A(n727), .B(KEYINPUT38), .ZN(n728) );
  NOR2_X1 U823 ( .A1(n729), .A2(n728), .ZN(n731) );
  NAND2_X1 U824 ( .A1(n897), .A2(G129), .ZN(n730) );
  NAND2_X1 U825 ( .A1(n731), .A2(n730), .ZN(n891) );
  AND2_X1 U826 ( .A1(n891), .A2(G1996), .ZN(n732) );
  NOR2_X1 U827 ( .A1(n733), .A2(n732), .ZN(n988) );
  NOR2_X1 U828 ( .A1(n988), .A2(n734), .ZN(n836) );
  INV_X1 U829 ( .A(n836), .ZN(n735) );
  NAND2_X1 U830 ( .A1(n839), .A2(n735), .ZN(n831) );
  NAND2_X1 U831 ( .A1(n737), .A2(n736), .ZN(n784) );
  NAND2_X1 U832 ( .A1(G8), .A2(n784), .ZN(n824) );
  NOR2_X1 U833 ( .A1(G1981), .A2(G305), .ZN(n738) );
  XOR2_X1 U834 ( .A(n738), .B(KEYINPUT24), .Z(n739) );
  NOR2_X1 U835 ( .A1(n824), .A2(n739), .ZN(n829) );
  NOR2_X1 U836 ( .A1(n784), .A2(n857), .ZN(n740) );
  XOR2_X1 U837 ( .A(n740), .B(KEYINPUT108), .Z(n742) );
  NAND2_X1 U838 ( .A1(n784), .A2(G1348), .ZN(n741) );
  NAND2_X1 U839 ( .A1(n742), .A2(n741), .ZN(n752) );
  INV_X1 U840 ( .A(G1996), .ZN(n869) );
  INV_X1 U841 ( .A(KEYINPUT26), .ZN(n743) );
  XNOR2_X1 U842 ( .A(n744), .B(n743), .ZN(n746) );
  NAND2_X1 U843 ( .A1(n784), .A2(G1341), .ZN(n745) );
  NAND2_X1 U844 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X2 U845 ( .A1(n748), .A2(n747), .ZN(n753) );
  NAND2_X1 U846 ( .A1(n753), .A2(n1018), .ZN(n750) );
  INV_X1 U847 ( .A(KEYINPUT107), .ZN(n749) );
  NAND2_X1 U848 ( .A1(n752), .A2(n751), .ZN(n756) );
  NOR2_X1 U849 ( .A1(n753), .A2(n1018), .ZN(n754) );
  XNOR2_X1 U850 ( .A(n754), .B(KEYINPUT109), .ZN(n755) );
  NAND2_X1 U851 ( .A1(n756), .A2(n755), .ZN(n763) );
  INV_X1 U852 ( .A(n784), .ZN(n770) );
  AND2_X1 U853 ( .A1(n770), .A2(G2072), .ZN(n758) );
  XNOR2_X1 U854 ( .A(KEYINPUT106), .B(KEYINPUT27), .ZN(n757) );
  XNOR2_X1 U855 ( .A(n758), .B(n757), .ZN(n760) );
  NAND2_X1 U856 ( .A1(n784), .A2(G1956), .ZN(n759) );
  NAND2_X1 U857 ( .A1(n760), .A2(n759), .ZN(n764) );
  NOR2_X1 U858 ( .A1(n1008), .A2(n764), .ZN(n761) );
  XOR2_X1 U859 ( .A(KEYINPUT110), .B(n761), .Z(n762) );
  NAND2_X1 U860 ( .A1(n763), .A2(n762), .ZN(n767) );
  NAND2_X1 U861 ( .A1(n1008), .A2(n764), .ZN(n765) );
  XNOR2_X1 U862 ( .A(n765), .B(KEYINPUT28), .ZN(n766) );
  NAND2_X1 U863 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U864 ( .A(n768), .B(KEYINPUT29), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n784), .A2(G1961), .ZN(n772) );
  XOR2_X1 U866 ( .A(G2078), .B(KEYINPUT25), .Z(n769) );
  XNOR2_X1 U867 ( .A(KEYINPUT104), .B(n769), .ZN(n954) );
  NAND2_X1 U868 ( .A1(n770), .A2(n954), .ZN(n771) );
  NAND2_X1 U869 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U870 ( .A(n773), .B(KEYINPUT105), .Z(n780) );
  NOR2_X1 U871 ( .A1(G301), .A2(n780), .ZN(n774) );
  XNOR2_X1 U872 ( .A(n776), .B(KEYINPUT111), .ZN(n797) );
  NOR2_X1 U873 ( .A1(G1966), .A2(n824), .ZN(n798) );
  NOR2_X1 U874 ( .A1(G2084), .A2(n784), .ZN(n799) );
  NOR2_X1 U875 ( .A1(n798), .A2(n799), .ZN(n777) );
  NAND2_X1 U876 ( .A1(G8), .A2(n777), .ZN(n778) );
  XNOR2_X1 U877 ( .A(KEYINPUT30), .B(n778), .ZN(n779) );
  NOR2_X1 U878 ( .A1(G168), .A2(n779), .ZN(n782) );
  AND2_X1 U879 ( .A1(G301), .A2(n780), .ZN(n781) );
  NOR2_X1 U880 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U881 ( .A(KEYINPUT31), .B(n783), .Z(n796) );
  INV_X1 U882 ( .A(G8), .ZN(n789) );
  NOR2_X1 U883 ( .A1(G2090), .A2(n784), .ZN(n786) );
  NOR2_X1 U884 ( .A1(G1971), .A2(n824), .ZN(n785) );
  NOR2_X1 U885 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U886 ( .A1(n787), .A2(G303), .ZN(n788) );
  OR2_X1 U887 ( .A1(n789), .A2(n788), .ZN(n791) );
  AND2_X1 U888 ( .A1(n796), .A2(n791), .ZN(n790) );
  NAND2_X1 U889 ( .A1(n797), .A2(n790), .ZN(n794) );
  INV_X1 U890 ( .A(n791), .ZN(n792) );
  OR2_X1 U891 ( .A1(n792), .A2(G286), .ZN(n793) );
  NAND2_X1 U892 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U893 ( .A(n795), .B(KEYINPUT32), .ZN(n820) );
  NAND2_X1 U894 ( .A1(n797), .A2(n796), .ZN(n803) );
  INV_X1 U895 ( .A(n798), .ZN(n801) );
  NAND2_X1 U896 ( .A1(G8), .A2(n799), .ZN(n800) );
  AND2_X1 U897 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U898 ( .A1(n803), .A2(n802), .ZN(n819) );
  NAND2_X1 U899 ( .A1(G1976), .A2(G288), .ZN(n1011) );
  AND2_X1 U900 ( .A1(n819), .A2(n1011), .ZN(n804) );
  NAND2_X1 U901 ( .A1(n820), .A2(n804), .ZN(n809) );
  INV_X1 U902 ( .A(n1011), .ZN(n806) );
  NOR2_X1 U903 ( .A1(G1976), .A2(G288), .ZN(n811) );
  NOR2_X1 U904 ( .A1(G1971), .A2(G303), .ZN(n805) );
  NOR2_X1 U905 ( .A1(n811), .A2(n805), .ZN(n1012) );
  OR2_X1 U906 ( .A1(n806), .A2(n1012), .ZN(n807) );
  INV_X1 U907 ( .A(KEYINPUT33), .ZN(n810) );
  AND2_X1 U908 ( .A1(n807), .A2(n810), .ZN(n808) );
  NAND2_X1 U909 ( .A1(n809), .A2(n808), .ZN(n818) );
  AND2_X1 U910 ( .A1(n810), .A2(n824), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n811), .A2(KEYINPUT33), .ZN(n812) );
  NOR2_X1 U912 ( .A1(n812), .A2(n824), .ZN(n814) );
  XOR2_X1 U913 ( .A(G1981), .B(G305), .Z(n1022) );
  INV_X1 U914 ( .A(n1022), .ZN(n813) );
  OR2_X1 U915 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U916 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U917 ( .A1(n818), .A2(n817), .ZN(n827) );
  NAND2_X1 U918 ( .A1(n820), .A2(n819), .ZN(n823) );
  NOR2_X1 U919 ( .A1(G2090), .A2(G303), .ZN(n821) );
  NAND2_X1 U920 ( .A1(G8), .A2(n821), .ZN(n822) );
  NAND2_X1 U921 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U922 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n828) );
  NOR2_X1 U924 ( .A1(n829), .A2(n828), .ZN(n830) );
  NOR2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n833) );
  XNOR2_X1 U926 ( .A(G1986), .B(G290), .ZN(n1007) );
  NAND2_X1 U927 ( .A1(n1007), .A2(n844), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n833), .A2(n832), .ZN(n847) );
  NOR2_X1 U929 ( .A1(G1996), .A2(n891), .ZN(n981) );
  NOR2_X1 U930 ( .A1(G1986), .A2(G290), .ZN(n834) );
  NOR2_X1 U931 ( .A1(G1991), .A2(n889), .ZN(n986) );
  NOR2_X1 U932 ( .A1(n834), .A2(n986), .ZN(n835) );
  NOR2_X1 U933 ( .A1(n836), .A2(n835), .ZN(n837) );
  NOR2_X1 U934 ( .A1(n981), .A2(n837), .ZN(n838) );
  XNOR2_X1 U935 ( .A(n838), .B(KEYINPUT39), .ZN(n840) );
  NAND2_X1 U936 ( .A1(n840), .A2(n839), .ZN(n842) );
  NAND2_X1 U937 ( .A1(n841), .A2(n910), .ZN(n995) );
  NAND2_X1 U938 ( .A1(n842), .A2(n995), .ZN(n843) );
  XNOR2_X1 U939 ( .A(KEYINPUT112), .B(n843), .ZN(n845) );
  NAND2_X1 U940 ( .A1(n845), .A2(n844), .ZN(n846) );
  NAND2_X1 U941 ( .A1(n847), .A2(n846), .ZN(n848) );
  XNOR2_X1 U942 ( .A(KEYINPUT40), .B(n848), .ZN(G329) );
  NAND2_X1 U943 ( .A1(G2106), .A2(n928), .ZN(G217) );
  AND2_X1 U944 ( .A1(G15), .A2(G2), .ZN(n849) );
  NAND2_X1 U945 ( .A1(G661), .A2(n849), .ZN(G259) );
  NAND2_X1 U946 ( .A1(G3), .A2(G1), .ZN(n850) );
  NAND2_X1 U947 ( .A1(n851), .A2(n850), .ZN(G188) );
  INV_X1 U949 ( .A(G120), .ZN(G236) );
  INV_X1 U950 ( .A(G96), .ZN(G221) );
  INV_X1 U951 ( .A(G69), .ZN(G235) );
  NOR2_X1 U952 ( .A1(n853), .A2(n852), .ZN(G325) );
  INV_X1 U953 ( .A(G325), .ZN(G261) );
  XOR2_X1 U954 ( .A(KEYINPUT42), .B(G2096), .Z(n856) );
  XOR2_X1 U955 ( .A(n854), .B(G2678), .Z(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n861) );
  XOR2_X1 U957 ( .A(KEYINPUT43), .B(G2090), .Z(n859) );
  XOR2_X1 U958 ( .A(n857), .B(G2072), .Z(n858) );
  XNOR2_X1 U959 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U960 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U961 ( .A(G2078), .B(G2084), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(G227) );
  INV_X1 U963 ( .A(G1971), .ZN(n1005) );
  XNOR2_X1 U964 ( .A(n1005), .B(G1961), .ZN(n865) );
  XNOR2_X1 U965 ( .A(G1986), .B(G1966), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U967 ( .A(n866), .B(G2474), .Z(n868) );
  XNOR2_X1 U968 ( .A(G1956), .B(G1976), .ZN(n867) );
  XNOR2_X1 U969 ( .A(n868), .B(n867), .ZN(n873) );
  XOR2_X1 U970 ( .A(KEYINPUT41), .B(G1981), .Z(n871) );
  XOR2_X1 U971 ( .A(n869), .B(G1991), .Z(n870) );
  XNOR2_X1 U972 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U973 ( .A(n873), .B(n872), .ZN(G229) );
  NAND2_X1 U974 ( .A1(G124), .A2(n897), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n874), .B(KEYINPUT44), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G112), .A2(n899), .ZN(n875) );
  XOR2_X1 U977 ( .A(KEYINPUT115), .B(n875), .Z(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n881) );
  NAND2_X1 U979 ( .A1(G100), .A2(n903), .ZN(n879) );
  NAND2_X1 U980 ( .A1(G136), .A2(n906), .ZN(n878) );
  NAND2_X1 U981 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U982 ( .A1(n881), .A2(n880), .ZN(G162) );
  NAND2_X1 U983 ( .A1(G118), .A2(n899), .ZN(n883) );
  NAND2_X1 U984 ( .A1(G130), .A2(n897), .ZN(n882) );
  NAND2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n888) );
  NAND2_X1 U986 ( .A1(G106), .A2(n903), .ZN(n885) );
  NAND2_X1 U987 ( .A1(G142), .A2(n906), .ZN(n884) );
  NAND2_X1 U988 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U989 ( .A(n886), .B(KEYINPUT45), .Z(n887) );
  NOR2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n890) );
  XNOR2_X1 U991 ( .A(n890), .B(n889), .ZN(n914) );
  XNOR2_X1 U992 ( .A(G162), .B(n891), .ZN(n892) );
  XNOR2_X1 U993 ( .A(n892), .B(n978), .ZN(n896) );
  XOR2_X1 U994 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n894) );
  XNOR2_X1 U995 ( .A(G160), .B(G164), .ZN(n893) );
  XNOR2_X1 U996 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U997 ( .A(n896), .B(n895), .ZN(n912) );
  NAND2_X1 U998 ( .A1(n897), .A2(G127), .ZN(n898) );
  XOR2_X1 U999 ( .A(KEYINPUT117), .B(n898), .Z(n901) );
  NAND2_X1 U1000 ( .A1(n899), .A2(G115), .ZN(n900) );
  NAND2_X1 U1001 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n902), .B(KEYINPUT47), .ZN(n905) );
  NAND2_X1 U1003 ( .A1(G103), .A2(n903), .ZN(n904) );
  NAND2_X1 U1004 ( .A1(n905), .A2(n904), .ZN(n909) );
  NAND2_X1 U1005 ( .A1(n906), .A2(G139), .ZN(n907) );
  XOR2_X1 U1006 ( .A(KEYINPUT116), .B(n907), .Z(n908) );
  NOR2_X1 U1007 ( .A1(n909), .A2(n908), .ZN(n989) );
  XNOR2_X1 U1008 ( .A(n910), .B(n989), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1010 ( .A(n914), .B(n913), .Z(n915) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n915), .ZN(G395) );
  XNOR2_X1 U1012 ( .A(G286), .B(n1018), .ZN(n917) );
  XNOR2_X1 U1013 ( .A(n917), .B(n916), .ZN(n919) );
  XOR2_X1 U1014 ( .A(n1027), .B(G171), .Z(n918) );
  XNOR2_X1 U1015 ( .A(n919), .B(n918), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n920), .ZN(G397) );
  NOR2_X1 U1017 ( .A1(G227), .A2(G229), .ZN(n921) );
  XNOR2_X1 U1018 ( .A(KEYINPUT49), .B(n921), .ZN(n922) );
  NOR2_X1 U1019 ( .A1(G401), .A2(n922), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n927), .ZN(n926) );
  XOR2_X1 U1023 ( .A(n926), .B(KEYINPUT118), .Z(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  INV_X1 U1025 ( .A(n927), .ZN(G319) );
  INV_X1 U1026 ( .A(G108), .ZN(G238) );
  INV_X1 U1027 ( .A(n928), .ZN(G223) );
  XOR2_X1 U1028 ( .A(G1976), .B(KEYINPUT126), .Z(n929) );
  XNOR2_X1 U1029 ( .A(G23), .B(n929), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(G1986), .B(G24), .ZN(n931) );
  XOR2_X1 U1031 ( .A(n1005), .B(G22), .Z(n930) );
  NOR2_X1 U1032 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1034 ( .A(n934), .B(KEYINPUT127), .ZN(n935) );
  XNOR2_X1 U1035 ( .A(KEYINPUT58), .B(n935), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(G1966), .B(G21), .ZN(n937) );
  XNOR2_X1 U1037 ( .A(G5), .B(G1961), .ZN(n936) );
  NOR2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n949) );
  XOR2_X1 U1040 ( .A(G1348), .B(KEYINPUT59), .Z(n940) );
  XNOR2_X1 U1041 ( .A(G4), .B(n940), .ZN(n942) );
  XNOR2_X1 U1042 ( .A(G20), .B(G1956), .ZN(n941) );
  NOR2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n946) );
  XNOR2_X1 U1044 ( .A(G1341), .B(G19), .ZN(n944) );
  XNOR2_X1 U1045 ( .A(G1981), .B(G6), .ZN(n943) );
  NOR2_X1 U1046 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1047 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1048 ( .A(KEYINPUT60), .B(n947), .ZN(n948) );
  NOR2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1050 ( .A(KEYINPUT61), .B(n950), .Z(n951) );
  NOR2_X1 U1051 ( .A1(G16), .A2(n951), .ZN(n976) );
  XOR2_X1 U1052 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n964) );
  XOR2_X1 U1053 ( .A(G1996), .B(G32), .Z(n953) );
  XOR2_X1 U1054 ( .A(G2067), .B(G26), .Z(n952) );
  NAND2_X1 U1055 ( .A1(n953), .A2(n952), .ZN(n956) );
  XNOR2_X1 U1056 ( .A(G27), .B(n954), .ZN(n955) );
  NOR2_X1 U1057 ( .A1(n956), .A2(n955), .ZN(n962) );
  XOR2_X1 U1058 ( .A(G33), .B(G2072), .Z(n957) );
  NAND2_X1 U1059 ( .A1(n957), .A2(G28), .ZN(n960) );
  XNOR2_X1 U1060 ( .A(G25), .B(G1991), .ZN(n958) );
  XNOR2_X1 U1061 ( .A(KEYINPUT120), .B(n958), .ZN(n959) );
  NOR2_X1 U1062 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1063 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1064 ( .A(n964), .B(n963), .ZN(n965) );
  XOR2_X1 U1065 ( .A(KEYINPUT53), .B(n965), .Z(n967) );
  XNOR2_X1 U1066 ( .A(G2090), .B(G35), .ZN(n966) );
  NOR2_X1 U1067 ( .A1(n967), .A2(n966), .ZN(n970) );
  XOR2_X1 U1068 ( .A(G2084), .B(G34), .Z(n968) );
  XNOR2_X1 U1069 ( .A(KEYINPUT54), .B(n968), .ZN(n969) );
  NAND2_X1 U1070 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1071 ( .A(KEYINPUT55), .B(n971), .Z(n973) );
  INV_X1 U1072 ( .A(G29), .ZN(n972) );
  NAND2_X1 U1073 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1074 ( .A1(G11), .A2(n974), .ZN(n975) );
  NOR2_X1 U1075 ( .A1(n976), .A2(n975), .ZN(n1004) );
  XOR2_X1 U1076 ( .A(G160), .B(G2084), .Z(n977) );
  NOR2_X1 U1077 ( .A1(n978), .A2(n977), .ZN(n984) );
  XNOR2_X1 U1078 ( .A(G2090), .B(G162), .ZN(n979) );
  XNOR2_X1 U1079 ( .A(n979), .B(KEYINPUT119), .ZN(n980) );
  NOR2_X1 U1080 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1081 ( .A(KEYINPUT51), .B(n982), .Z(n983) );
  NAND2_X1 U1082 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1083 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1084 ( .A1(n988), .A2(n987), .ZN(n994) );
  XOR2_X1 U1085 ( .A(G164), .B(G2078), .Z(n991) );
  XOR2_X1 U1086 ( .A(G2072), .B(n989), .Z(n990) );
  NOR2_X1 U1087 ( .A1(n991), .A2(n990), .ZN(n992) );
  XOR2_X1 U1088 ( .A(KEYINPUT50), .B(n992), .Z(n993) );
  NOR2_X1 U1089 ( .A1(n994), .A2(n993), .ZN(n996) );
  NAND2_X1 U1090 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1092 ( .A(KEYINPUT52), .B(n999), .ZN(n1001) );
  INV_X1 U1093 ( .A(KEYINPUT55), .ZN(n1000) );
  NAND2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1095 ( .A1(n1002), .A2(G29), .ZN(n1003) );
  NAND2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1034) );
  XOR2_X1 U1097 ( .A(KEYINPUT56), .B(G16), .Z(n1032) );
  NOR2_X1 U1098 ( .A1(G166), .A2(n1005), .ZN(n1006) );
  NOR2_X1 U1099 ( .A1(n1007), .A2(n1006), .ZN(n1010) );
  XOR2_X1 U1100 ( .A(G1956), .B(n1008), .Z(n1009) );
  NAND2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1104 ( .A(KEYINPUT123), .B(n1015), .Z(n1017) );
  XOR2_X1 U1105 ( .A(G301), .B(G1961), .Z(n1016) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1020) );
  XOR2_X1 U1107 ( .A(G1348), .B(n1018), .Z(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1109 ( .A(KEYINPUT124), .B(n1021), .ZN(n1026) );
  XNOR2_X1 U1110 ( .A(G1966), .B(G168), .ZN(n1023) );
  NAND2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1112 ( .A(n1024), .B(KEYINPUT57), .ZN(n1025) );
  NAND2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1029) );
  XOR2_X1 U1114 ( .A(G1341), .B(n1027), .Z(n1028) );
  NOR2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1116 ( .A(KEYINPUT125), .B(n1030), .Z(n1031) );
  NOR2_X1 U1117 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1118 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XOR2_X1 U1119 ( .A(n1035), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1120 ( .A(G150), .ZN(G311) );
endmodule

