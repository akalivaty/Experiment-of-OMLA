

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735;

  XNOR2_X1 U370 ( .A(n347), .B(n389), .ZN(n437) );
  XNOR2_X1 U371 ( .A(n348), .B(G119), .ZN(n347) );
  NOR2_X2 U372 ( .A1(n620), .A2(n636), .ZN(n621) );
  NOR2_X2 U373 ( .A1(n607), .A2(n636), .ZN(n608) );
  NOR2_X2 U374 ( .A1(n614), .A2(n636), .ZN(n615) );
  AND2_X2 U375 ( .A1(n591), .A2(KEYINPUT64), .ZN(n596) );
  NOR2_X2 U376 ( .A1(n625), .A2(n636), .ZN(n627) );
  XNOR2_X2 U377 ( .A(n724), .B(n350), .ZN(n463) );
  OR2_X2 U378 ( .A1(n655), .A2(n654), .ZN(n649) );
  NOR2_X2 U379 ( .A1(n598), .A2(n597), .ZN(n600) );
  XNOR2_X2 U380 ( .A(n427), .B(n426), .ZN(n491) );
  NOR2_X1 U381 ( .A1(n550), .A2(n549), .ZN(n562) );
  INV_X2 U382 ( .A(G953), .ZN(n725) );
  NOR2_X1 U383 ( .A1(n524), .A2(n523), .ZN(n700) );
  NOR2_X1 U384 ( .A1(n648), .A2(n563), .ZN(n555) );
  XNOR2_X1 U385 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U386 ( .A(n600), .B(n599), .ZN(n638) );
  NOR2_X1 U387 ( .A1(n733), .A2(n734), .ZN(n520) );
  NAND2_X1 U388 ( .A1(n425), .A2(n567), .ZN(n427) );
  XNOR2_X1 U389 ( .A(n377), .B(n376), .ZN(n447) );
  NAND2_X1 U390 ( .A1(n645), .A2(n638), .ZN(n642) );
  XNOR2_X2 U391 ( .A(n396), .B(n461), .ZN(n711) );
  XNOR2_X1 U392 ( .A(n535), .B(n534), .ZN(n539) );
  INV_X1 U393 ( .A(G475), .ZN(n363) );
  XNOR2_X1 U394 ( .A(n543), .B(n542), .ZN(n548) );
  INV_X1 U395 ( .A(KEYINPUT45), .ZN(n599) );
  NOR2_X1 U396 ( .A1(n541), .A2(n540), .ZN(n543) );
  NOR2_X1 U397 ( .A1(n565), .A2(n502), .ZN(n503) );
  XNOR2_X1 U398 ( .A(n479), .B(KEYINPUT68), .ZN(n513) );
  BUF_X1 U399 ( .A(n638), .Z(n717) );
  XNOR2_X1 U400 ( .A(n442), .B(n441), .ZN(n446) );
  INV_X1 U401 ( .A(KEYINPUT84), .ZN(n374) );
  INV_X1 U402 ( .A(G104), .ZN(n352) );
  AND2_X2 U403 ( .A1(n349), .A2(n409), .ZN(n629) );
  XNOR2_X1 U404 ( .A(n642), .B(KEYINPUT2), .ZN(n349) );
  NOR2_X1 U405 ( .A1(n531), .A2(n655), .ZN(n508) );
  NAND2_X1 U406 ( .A1(n522), .A2(n423), .ZN(n424) );
  XNOR2_X1 U407 ( .A(n364), .B(n363), .ZN(n365) );
  NOR2_X1 U408 ( .A1(n725), .A2(G952), .ZN(n636) );
  XNOR2_X1 U409 ( .A(n437), .B(n391), .ZN(n396) );
  XNOR2_X2 U410 ( .A(G116), .B(KEYINPUT3), .ZN(n348) );
  NOR2_X2 U411 ( .A1(n548), .A2(n547), .ZN(n645) );
  BUF_X1 U412 ( .A(n629), .Z(n633) );
  BUF_X1 U413 ( .A(n507), .Z(n529) );
  INV_X1 U414 ( .A(KEYINPUT82), .ZN(n534) );
  NOR2_X1 U415 ( .A1(G953), .A2(G237), .ZN(n433) );
  NAND2_X1 U416 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U417 ( .A(n353), .B(n352), .ZN(n355) );
  INV_X1 U418 ( .A(KEYINPUT48), .ZN(n542) );
  XNOR2_X1 U419 ( .A(G119), .B(G110), .ZN(n444) );
  XNOR2_X1 U420 ( .A(n355), .B(n354), .ZN(n361) );
  INV_X1 U421 ( .A(KEYINPUT109), .ZN(n514) );
  XNOR2_X1 U422 ( .A(n514), .B(KEYINPUT28), .ZN(n515) );
  XNOR2_X1 U423 ( .A(n446), .B(n445), .ZN(n449) );
  XNOR2_X1 U424 ( .A(n516), .B(n515), .ZN(n518) );
  INV_X1 U425 ( .A(n556), .ZN(n557) );
  XNOR2_X1 U426 ( .A(n366), .B(n365), .ZN(n528) );
  INV_X1 U427 ( .A(KEYINPUT104), .ZN(n383) );
  INV_X1 U428 ( .A(G146), .ZN(n350) );
  XNOR2_X1 U429 ( .A(n350), .B(G125), .ZN(n398) );
  XNOR2_X1 U430 ( .A(n398), .B(G140), .ZN(n351) );
  XNOR2_X1 U431 ( .A(n351), .B(KEYINPUT10), .ZN(n723) );
  NAND2_X1 U432 ( .A1(G214), .A2(n433), .ZN(n353) );
  XOR2_X1 U433 ( .A(G122), .B(G113), .Z(n354) );
  XOR2_X1 U434 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n357) );
  XNOR2_X1 U435 ( .A(KEYINPUT11), .B(KEYINPUT99), .ZN(n356) );
  XNOR2_X1 U436 ( .A(n357), .B(n356), .ZN(n359) );
  XNOR2_X1 U437 ( .A(G131), .B(G143), .ZN(n358) );
  XNOR2_X1 U438 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U439 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U440 ( .A(n723), .B(n362), .ZN(n617) );
  NOR2_X1 U441 ( .A1(G902), .A2(n617), .ZN(n366) );
  INV_X1 U442 ( .A(KEYINPUT13), .ZN(n364) );
  XOR2_X1 U443 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n368) );
  XNOR2_X1 U444 ( .A(G122), .B(KEYINPUT9), .ZN(n367) );
  XNOR2_X1 U445 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U446 ( .A(KEYINPUT102), .B(KEYINPUT7), .Z(n370) );
  XNOR2_X1 U447 ( .A(G116), .B(G107), .ZN(n369) );
  XNOR2_X1 U448 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U449 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U450 ( .A(G143), .B(G128), .ZN(n400) );
  XNOR2_X1 U451 ( .A(n400), .B(G134), .ZN(n432) );
  XNOR2_X1 U452 ( .A(n373), .B(n432), .ZN(n379) );
  XOR2_X1 U453 ( .A(KEYINPUT8), .B(KEYINPUT67), .Z(n377) );
  NAND2_X1 U454 ( .A1(G234), .A2(n725), .ZN(n375) );
  NAND2_X1 U455 ( .A1(n447), .A2(G217), .ZN(n378) );
  XNOR2_X1 U456 ( .A(n379), .B(n378), .ZN(n635) );
  INV_X1 U457 ( .A(G902), .ZN(n451) );
  NAND2_X1 U458 ( .A1(n635), .A2(n451), .ZN(n381) );
  XOR2_X1 U459 ( .A(KEYINPUT103), .B(G478), .Z(n380) );
  XNOR2_X1 U460 ( .A(n381), .B(n380), .ZN(n527) );
  NOR2_X1 U461 ( .A1(n528), .A2(n527), .ZN(n382) );
  XNOR2_X1 U462 ( .A(n383), .B(n382), .ZN(n652) );
  XNOR2_X1 U463 ( .A(KEYINPUT15), .B(G902), .ZN(n601) );
  NAND2_X1 U464 ( .A1(G234), .A2(n601), .ZN(n384) );
  XNOR2_X1 U465 ( .A(KEYINPUT20), .B(n384), .ZN(n452) );
  NAND2_X1 U466 ( .A1(n452), .A2(G221), .ZN(n385) );
  XOR2_X1 U467 ( .A(n385), .B(KEYINPUT21), .Z(n665) );
  INV_X1 U468 ( .A(n665), .ZN(n386) );
  NOR2_X1 U469 ( .A1(n652), .A2(n386), .ZN(n388) );
  INV_X1 U470 ( .A(KEYINPUT105), .ZN(n387) );
  XNOR2_X1 U471 ( .A(n388), .B(n387), .ZN(n425) );
  XNOR2_X1 U472 ( .A(G113), .B(KEYINPUT91), .ZN(n389) );
  XNOR2_X1 U473 ( .A(KEYINPUT71), .B(KEYINPUT16), .ZN(n390) );
  XNOR2_X1 U474 ( .A(n390), .B(G122), .ZN(n391) );
  XNOR2_X1 U475 ( .A(G107), .B(G104), .ZN(n393) );
  INV_X1 U476 ( .A(G110), .ZN(n392) );
  XNOR2_X1 U477 ( .A(n393), .B(n392), .ZN(n395) );
  XNOR2_X1 U478 ( .A(G101), .B(KEYINPUT73), .ZN(n394) );
  XNOR2_X1 U479 ( .A(n395), .B(n394), .ZN(n461) );
  INV_X1 U480 ( .A(KEYINPUT66), .ZN(n397) );
  XNOR2_X1 U481 ( .A(n397), .B(KEYINPUT4), .ZN(n429) );
  XNOR2_X1 U482 ( .A(n398), .B(n429), .ZN(n402) );
  XNOR2_X1 U483 ( .A(KEYINPUT78), .B(KEYINPUT90), .ZN(n399) );
  XNOR2_X1 U484 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U485 ( .A(n402), .B(n401), .ZN(n407) );
  XOR2_X1 U486 ( .A(KEYINPUT17), .B(KEYINPUT77), .Z(n405) );
  NAND2_X1 U487 ( .A1(G224), .A2(n725), .ZN(n403) );
  XNOR2_X1 U488 ( .A(n403), .B(KEYINPUT18), .ZN(n404) );
  XNOR2_X1 U489 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U490 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U491 ( .A(n711), .B(n408), .ZN(n604) );
  INV_X1 U492 ( .A(n601), .ZN(n409) );
  OR2_X2 U493 ( .A1(n604), .A2(n409), .ZN(n413) );
  INV_X1 U494 ( .A(G237), .ZN(n410) );
  NAND2_X1 U495 ( .A1(n451), .A2(n410), .ZN(n414) );
  NAND2_X1 U496 ( .A1(n414), .A2(G210), .ZN(n411) );
  XNOR2_X1 U497 ( .A(n411), .B(KEYINPUT92), .ZN(n412) );
  XNOR2_X2 U498 ( .A(n413), .B(n412), .ZN(n507) );
  NAND2_X1 U499 ( .A1(n414), .A2(G214), .ZN(n415) );
  XNOR2_X1 U500 ( .A(n415), .B(KEYINPUT93), .ZN(n654) );
  OR2_X2 U501 ( .A1(n507), .A2(n654), .ZN(n418) );
  INV_X1 U502 ( .A(KEYINPUT75), .ZN(n416) );
  XNOR2_X1 U503 ( .A(n416), .B(KEYINPUT19), .ZN(n417) );
  XNOR2_X2 U504 ( .A(n418), .B(n417), .ZN(n522) );
  NAND2_X1 U505 ( .A1(G234), .A2(G237), .ZN(n419) );
  XNOR2_X1 U506 ( .A(n419), .B(KEYINPUT14), .ZN(n420) );
  AND2_X1 U507 ( .A1(n420), .A2(G952), .ZN(n680) );
  AND2_X1 U508 ( .A1(n680), .A2(n725), .ZN(n476) );
  NAND2_X1 U509 ( .A1(G902), .A2(n420), .ZN(n472) );
  XOR2_X1 U510 ( .A(G898), .B(KEYINPUT94), .Z(n716) );
  NAND2_X1 U511 ( .A1(G953), .A2(n716), .ZN(n712) );
  NOR2_X1 U512 ( .A1(n472), .A2(n712), .ZN(n421) );
  NOR2_X1 U513 ( .A1(n476), .A2(n421), .ZN(n422) );
  XNOR2_X1 U514 ( .A(n422), .B(KEYINPUT95), .ZN(n423) );
  XNOR2_X2 U515 ( .A(n424), .B(KEYINPUT0), .ZN(n563) );
  INV_X1 U516 ( .A(n563), .ZN(n567) );
  INV_X1 U517 ( .A(KEYINPUT22), .ZN(n426) );
  XNOR2_X1 U518 ( .A(G137), .B(G131), .ZN(n428) );
  XNOR2_X1 U519 ( .A(n429), .B(n428), .ZN(n430) );
  INV_X1 U520 ( .A(n430), .ZN(n431) );
  XNOR2_X2 U521 ( .A(n432), .B(n431), .ZN(n724) );
  XOR2_X1 U522 ( .A(G101), .B(KEYINPUT5), .Z(n435) );
  NAND2_X1 U523 ( .A1(n433), .A2(G210), .ZN(n434) );
  XNOR2_X1 U524 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U525 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U526 ( .A(n463), .B(n438), .ZN(n622) );
  NAND2_X1 U527 ( .A1(n622), .A2(n451), .ZN(n440) );
  INV_X1 U528 ( .A(G472), .ZN(n439) );
  XNOR2_X2 U529 ( .A(n440), .B(n439), .ZN(n561) );
  XNOR2_X1 U530 ( .A(n561), .B(KEYINPUT6), .ZN(n551) );
  XOR2_X1 U531 ( .A(KEYINPUT23), .B(KEYINPUT96), .Z(n442) );
  XNOR2_X1 U532 ( .A(G137), .B(G128), .ZN(n441) );
  INV_X1 U533 ( .A(KEYINPUT24), .ZN(n443) );
  XNOR2_X1 U534 ( .A(n444), .B(n443), .ZN(n445) );
  NAND2_X1 U535 ( .A1(n447), .A2(G221), .ZN(n448) );
  XNOR2_X1 U536 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U537 ( .A(n450), .B(n723), .ZN(n631) );
  NAND2_X1 U538 ( .A1(n631), .A2(n451), .ZN(n458) );
  XOR2_X1 U539 ( .A(KEYINPUT76), .B(KEYINPUT97), .Z(n454) );
  NAND2_X1 U540 ( .A1(n452), .A2(G217), .ZN(n453) );
  XNOR2_X1 U541 ( .A(n454), .B(n453), .ZN(n456) );
  INV_X1 U542 ( .A(KEYINPUT25), .ZN(n455) );
  XNOR2_X1 U543 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U544 ( .A(n458), .B(n457), .ZN(n501) );
  BUF_X1 U545 ( .A(n501), .Z(n666) );
  XNOR2_X1 U546 ( .A(KEYINPUT69), .B(G469), .ZN(n466) );
  NAND2_X1 U547 ( .A1(G227), .A2(n725), .ZN(n459) );
  XNOR2_X1 U548 ( .A(n459), .B(G140), .ZN(n460) );
  XNOR2_X1 U549 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U550 ( .A(n463), .B(n462), .ZN(n611) );
  NOR2_X1 U551 ( .A1(G902), .A2(n611), .ZN(n464) );
  INV_X1 U552 ( .A(n464), .ZN(n465) );
  XNOR2_X1 U553 ( .A(n466), .B(n465), .ZN(n500) );
  XNOR2_X1 U554 ( .A(n500), .B(KEYINPUT1), .ZN(n550) );
  INV_X1 U555 ( .A(n550), .ZN(n662) );
  INV_X1 U556 ( .A(n662), .ZN(n483) );
  NAND2_X1 U557 ( .A1(n666), .A2(n483), .ZN(n467) );
  NOR2_X1 U558 ( .A1(n551), .A2(n467), .ZN(n468) );
  NAND2_X1 U559 ( .A1(n491), .A2(n468), .ZN(n571) );
  XOR2_X1 U560 ( .A(G101), .B(KEYINPUT113), .Z(n469) );
  XNOR2_X1 U561 ( .A(n571), .B(n469), .ZN(G3) );
  NOR2_X1 U562 ( .A1(n666), .A2(n662), .ZN(n470) );
  AND2_X1 U563 ( .A1(n561), .A2(n470), .ZN(n471) );
  AND2_X1 U564 ( .A1(n491), .A2(n471), .ZN(n576) );
  INV_X1 U565 ( .A(n576), .ZN(n592) );
  XNOR2_X1 U566 ( .A(n592), .B(G110), .ZN(G12) );
  NOR2_X1 U567 ( .A1(G900), .A2(n472), .ZN(n473) );
  NAND2_X1 U568 ( .A1(G953), .A2(n473), .ZN(n474) );
  XOR2_X1 U569 ( .A(KEYINPUT106), .B(n474), .Z(n475) );
  NOR2_X1 U570 ( .A1(n476), .A2(n475), .ZN(n477) );
  XOR2_X1 U571 ( .A(KEYINPUT81), .B(n477), .Z(n502) );
  NOR2_X1 U572 ( .A1(n666), .A2(n502), .ZN(n478) );
  NAND2_X1 U573 ( .A1(n478), .A2(n665), .ZN(n479) );
  INV_X1 U574 ( .A(n527), .ZN(n480) );
  NAND2_X1 U575 ( .A1(n528), .A2(n480), .ZN(n702) );
  NOR2_X1 U576 ( .A1(n513), .A2(n702), .ZN(n481) );
  NAND2_X1 U577 ( .A1(n551), .A2(n481), .ZN(n482) );
  NOR2_X1 U578 ( .A1(n482), .A2(n654), .ZN(n496) );
  XOR2_X1 U579 ( .A(n496), .B(KEYINPUT107), .Z(n484) );
  NAND2_X1 U580 ( .A1(n484), .A2(n483), .ZN(n485) );
  XNOR2_X1 U581 ( .A(n485), .B(KEYINPUT43), .ZN(n486) );
  XNOR2_X1 U582 ( .A(KEYINPUT108), .B(n486), .ZN(n487) );
  NAND2_X1 U583 ( .A1(n487), .A2(n529), .ZN(n545) );
  XNOR2_X1 U584 ( .A(G140), .B(KEYINPUT116), .ZN(n488) );
  XNOR2_X1 U585 ( .A(n545), .B(n488), .ZN(G42) );
  OR2_X1 U586 ( .A1(n666), .A2(n550), .ZN(n489) );
  NOR2_X1 U587 ( .A1(n489), .A2(n551), .ZN(n490) );
  NAND2_X1 U588 ( .A1(n491), .A2(n490), .ZN(n493) );
  XNOR2_X1 U589 ( .A(KEYINPUT80), .B(KEYINPUT32), .ZN(n492) );
  XNOR2_X2 U590 ( .A(n493), .B(n492), .ZN(n593) );
  XNOR2_X1 U591 ( .A(G119), .B(KEYINPUT126), .ZN(n494) );
  XNOR2_X1 U592 ( .A(n593), .B(n494), .ZN(G21) );
  INV_X1 U593 ( .A(KEYINPUT2), .ZN(n640) );
  INV_X1 U594 ( .A(n529), .ZN(n495) );
  NAND2_X1 U595 ( .A1(n496), .A2(n495), .ZN(n498) );
  XOR2_X1 U596 ( .A(KEYINPUT112), .B(KEYINPUT36), .Z(n497) );
  XNOR2_X1 U597 ( .A(n498), .B(n497), .ZN(n499) );
  NAND2_X1 U598 ( .A1(n499), .A2(n662), .ZN(n707) );
  INV_X1 U599 ( .A(n500), .ZN(n517) );
  NAND2_X1 U600 ( .A1(n665), .A2(n501), .ZN(n549) );
  INV_X1 U601 ( .A(n549), .ZN(n661) );
  NAND2_X1 U602 ( .A1(n517), .A2(n661), .ZN(n565) );
  XNOR2_X1 U603 ( .A(n503), .B(KEYINPUT74), .ZN(n506) );
  NOR2_X1 U604 ( .A1(n654), .A2(n561), .ZN(n504) );
  XNOR2_X1 U605 ( .A(KEYINPUT30), .B(n504), .ZN(n505) );
  NAND2_X1 U606 ( .A1(n506), .A2(n505), .ZN(n531) );
  XOR2_X1 U607 ( .A(KEYINPUT38), .B(n507), .Z(n655) );
  XNOR2_X1 U608 ( .A(n508), .B(KEYINPUT39), .ZN(n544) );
  NOR2_X1 U609 ( .A1(n702), .A2(n544), .ZN(n510) );
  XNOR2_X1 U610 ( .A(KEYINPUT40), .B(KEYINPUT110), .ZN(n509) );
  XNOR2_X1 U611 ( .A(n510), .B(n509), .ZN(n733) );
  NOR2_X1 U612 ( .A1(n652), .A2(n649), .ZN(n512) );
  XOR2_X1 U613 ( .A(KEYINPUT111), .B(KEYINPUT41), .Z(n511) );
  XNOR2_X1 U614 ( .A(n512), .B(n511), .ZN(n682) );
  NOR2_X1 U615 ( .A1(n513), .A2(n561), .ZN(n516) );
  NAND2_X1 U616 ( .A1(n518), .A2(n517), .ZN(n524) );
  NOR2_X1 U617 ( .A1(n682), .A2(n524), .ZN(n519) );
  XNOR2_X1 U618 ( .A(KEYINPUT42), .B(n519), .ZN(n734) );
  XNOR2_X1 U619 ( .A(n520), .B(KEYINPUT46), .ZN(n521) );
  NAND2_X1 U620 ( .A1(n707), .A2(n521), .ZN(n541) );
  INV_X1 U621 ( .A(n522), .ZN(n523) );
  INV_X1 U622 ( .A(n528), .ZN(n525) );
  NAND2_X1 U623 ( .A1(n525), .A2(n527), .ZN(n705) );
  AND2_X1 U624 ( .A1(n705), .A2(n702), .ZN(n650) );
  INV_X1 U625 ( .A(n650), .ZN(n568) );
  NAND2_X1 U626 ( .A1(n700), .A2(n568), .ZN(n526) );
  NAND2_X1 U627 ( .A1(n526), .A2(KEYINPUT47), .ZN(n533) );
  NAND2_X1 U628 ( .A1(n528), .A2(n527), .ZN(n556) );
  OR2_X1 U629 ( .A1(n556), .A2(n529), .ZN(n530) );
  NOR2_X1 U630 ( .A1(n531), .A2(n530), .ZN(n698) );
  XNOR2_X1 U631 ( .A(KEYINPUT83), .B(n698), .ZN(n532) );
  NAND2_X1 U632 ( .A1(n533), .A2(n532), .ZN(n535) );
  NOR2_X1 U633 ( .A1(KEYINPUT47), .A2(n650), .ZN(n536) );
  XNOR2_X1 U634 ( .A(n536), .B(KEYINPUT72), .ZN(n537) );
  NAND2_X1 U635 ( .A1(n700), .A2(n537), .ZN(n538) );
  NOR2_X1 U636 ( .A1(n544), .A2(n705), .ZN(n710) );
  INV_X1 U637 ( .A(n710), .ZN(n546) );
  NAND2_X1 U638 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U639 ( .A1(n562), .A2(n551), .ZN(n554) );
  INV_X1 U640 ( .A(KEYINPUT70), .ZN(n552) );
  XNOR2_X1 U641 ( .A(n552), .B(KEYINPUT33), .ZN(n553) );
  XNOR2_X1 U642 ( .A(n554), .B(n553), .ZN(n648) );
  XNOR2_X1 U643 ( .A(n555), .B(KEYINPUT34), .ZN(n558) );
  NAND2_X1 U644 ( .A1(n558), .A2(n557), .ZN(n560) );
  XNOR2_X1 U645 ( .A(KEYINPUT79), .B(KEYINPUT35), .ZN(n559) );
  XNOR2_X2 U646 ( .A(n560), .B(n559), .ZN(n628) );
  INV_X1 U647 ( .A(n628), .ZN(n574) );
  NOR2_X1 U648 ( .A1(n574), .A2(KEYINPUT86), .ZN(n573) );
  INV_X1 U649 ( .A(n561), .ZN(n669) );
  NAND2_X1 U650 ( .A1(n669), .A2(n562), .ZN(n672) );
  NOR2_X1 U651 ( .A1(n563), .A2(n672), .ZN(n564) );
  XNOR2_X1 U652 ( .A(n564), .B(KEYINPUT31), .ZN(n704) );
  NOR2_X1 U653 ( .A1(n669), .A2(n565), .ZN(n566) );
  NAND2_X1 U654 ( .A1(n567), .A2(n566), .ZN(n692) );
  NAND2_X1 U655 ( .A1(n704), .A2(n692), .ZN(n569) );
  NAND2_X1 U656 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U657 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U658 ( .A1(n573), .A2(n572), .ZN(n586) );
  NAND2_X1 U659 ( .A1(n574), .A2(KEYINPUT86), .ZN(n575) );
  NAND2_X1 U660 ( .A1(n575), .A2(KEYINPUT44), .ZN(n584) );
  NOR2_X1 U661 ( .A1(n576), .A2(KEYINPUT87), .ZN(n577) );
  AND2_X1 U662 ( .A1(n628), .A2(n577), .ZN(n578) );
  NAND2_X1 U663 ( .A1(n578), .A2(n593), .ZN(n582) );
  INV_X1 U664 ( .A(KEYINPUT44), .ZN(n587) );
  NAND2_X1 U665 ( .A1(n587), .A2(KEYINPUT64), .ZN(n580) );
  INV_X1 U666 ( .A(KEYINPUT86), .ZN(n579) );
  NOR2_X1 U667 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U668 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U669 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U670 ( .A1(n586), .A2(n585), .ZN(n598) );
  NAND2_X1 U671 ( .A1(n628), .A2(KEYINPUT87), .ZN(n588) );
  NAND2_X1 U672 ( .A1(n588), .A2(n587), .ZN(n590) );
  NAND2_X1 U673 ( .A1(n593), .A2(n592), .ZN(n589) );
  NAND2_X1 U674 ( .A1(n590), .A2(n589), .ZN(n591) );
  AND2_X1 U675 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U676 ( .A1(n594), .A2(KEYINPUT64), .ZN(n595) );
  NOR2_X1 U677 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U678 ( .A1(n629), .A2(G210), .ZN(n606) );
  XNOR2_X1 U679 ( .A(KEYINPUT89), .B(KEYINPUT54), .ZN(n602) );
  XNOR2_X1 U680 ( .A(n602), .B(KEYINPUT55), .ZN(n603) );
  XNOR2_X1 U681 ( .A(n604), .B(n603), .ZN(n605) );
  XNOR2_X1 U682 ( .A(n606), .B(n605), .ZN(n607) );
  XNOR2_X1 U683 ( .A(n608), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U684 ( .A1(n629), .A2(G469), .ZN(n613) );
  XNOR2_X1 U685 ( .A(KEYINPUT121), .B(KEYINPUT57), .ZN(n609) );
  XNOR2_X1 U686 ( .A(n609), .B(KEYINPUT58), .ZN(n610) );
  XNOR2_X1 U687 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U688 ( .A(n613), .B(n612), .ZN(n614) );
  XNOR2_X1 U689 ( .A(n615), .B(KEYINPUT122), .ZN(G54) );
  NAND2_X1 U690 ( .A1(n629), .A2(G475), .ZN(n619) );
  XNOR2_X1 U691 ( .A(KEYINPUT65), .B(KEYINPUT59), .ZN(n616) );
  XNOR2_X1 U692 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U693 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U694 ( .A(n621), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U695 ( .A1(n629), .A2(G472), .ZN(n624) );
  XOR2_X1 U696 ( .A(n622), .B(KEYINPUT62), .Z(n623) );
  XNOR2_X1 U697 ( .A(n624), .B(n623), .ZN(n625) );
  XOR2_X1 U698 ( .A(KEYINPUT88), .B(KEYINPUT63), .Z(n626) );
  XNOR2_X1 U699 ( .A(n627), .B(n626), .ZN(G57) );
  XNOR2_X1 U700 ( .A(n628), .B(G122), .ZN(G24) );
  NAND2_X1 U701 ( .A1(n633), .A2(G217), .ZN(n630) );
  XOR2_X1 U702 ( .A(n631), .B(n630), .Z(n632) );
  NOR2_X1 U703 ( .A1(n632), .A2(n636), .ZN(G66) );
  NAND2_X1 U704 ( .A1(n633), .A2(G478), .ZN(n634) );
  XOR2_X1 U705 ( .A(n635), .B(n634), .Z(n637) );
  NOR2_X1 U706 ( .A1(n637), .A2(n636), .ZN(G63) );
  XNOR2_X1 U707 ( .A(n717), .B(KEYINPUT85), .ZN(n639) );
  NOR2_X1 U708 ( .A1(n639), .A2(KEYINPUT2), .ZN(n644) );
  NOR2_X1 U709 ( .A1(n640), .A2(KEYINPUT85), .ZN(n641) );
  AND2_X1 U710 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U711 ( .A1(n644), .A2(n643), .ZN(n647) );
  NOR2_X1 U712 ( .A1(n645), .A2(KEYINPUT2), .ZN(n646) );
  NOR2_X1 U713 ( .A1(n647), .A2(n646), .ZN(n687) );
  OR2_X1 U714 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U715 ( .A(KEYINPUT118), .B(n651), .ZN(n653) );
  NAND2_X1 U716 ( .A1(n653), .A2(n652), .ZN(n658) );
  AND2_X1 U717 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U718 ( .A1(KEYINPUT118), .A2(n656), .ZN(n657) );
  NAND2_X1 U719 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U720 ( .A1(n648), .A2(n659), .ZN(n660) );
  XOR2_X1 U721 ( .A(KEYINPUT119), .B(n660), .Z(n677) );
  NOR2_X1 U722 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U723 ( .A(n663), .B(KEYINPUT50), .ZN(n664) );
  XNOR2_X1 U724 ( .A(n664), .B(KEYINPUT117), .ZN(n671) );
  NOR2_X1 U725 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U726 ( .A(KEYINPUT49), .B(n667), .Z(n668) );
  NOR2_X1 U727 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U728 ( .A1(n671), .A2(n670), .ZN(n673) );
  NAND2_X1 U729 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U730 ( .A(KEYINPUT51), .B(n674), .ZN(n675) );
  NOR2_X1 U731 ( .A1(n682), .A2(n675), .ZN(n676) );
  NOR2_X1 U732 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U733 ( .A(n678), .B(KEYINPUT52), .ZN(n679) );
  XOR2_X1 U734 ( .A(n679), .B(KEYINPUT120), .Z(n681) );
  NAND2_X1 U735 ( .A1(n681), .A2(n680), .ZN(n685) );
  NOR2_X1 U736 ( .A1(n682), .A2(n648), .ZN(n683) );
  NOR2_X1 U737 ( .A1(n683), .A2(G953), .ZN(n684) );
  NAND2_X1 U738 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U739 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U740 ( .A(n688), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U741 ( .A1(n702), .A2(n692), .ZN(n689) );
  XOR2_X1 U742 ( .A(G104), .B(n689), .Z(G6) );
  XOR2_X1 U743 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n691) );
  XNOR2_X1 U744 ( .A(G107), .B(KEYINPUT26), .ZN(n690) );
  XNOR2_X1 U745 ( .A(n691), .B(n690), .ZN(n694) );
  NOR2_X1 U746 ( .A1(n705), .A2(n692), .ZN(n693) );
  XOR2_X1 U747 ( .A(n694), .B(n693), .Z(G9) );
  XOR2_X1 U748 ( .A(G128), .B(KEYINPUT29), .Z(n697) );
  INV_X1 U749 ( .A(n705), .ZN(n695) );
  NAND2_X1 U750 ( .A1(n700), .A2(n695), .ZN(n696) );
  XNOR2_X1 U751 ( .A(n697), .B(n696), .ZN(G30) );
  XOR2_X1 U752 ( .A(G143), .B(n698), .Z(G45) );
  INV_X1 U753 ( .A(n702), .ZN(n699) );
  NAND2_X1 U754 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U755 ( .A(n701), .B(G146), .ZN(G48) );
  NOR2_X1 U756 ( .A1(n702), .A2(n704), .ZN(n703) );
  XOR2_X1 U757 ( .A(G113), .B(n703), .Z(G15) );
  NOR2_X1 U758 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U759 ( .A(G116), .B(n706), .Z(G18) );
  XNOR2_X1 U760 ( .A(KEYINPUT37), .B(KEYINPUT115), .ZN(n708) );
  XNOR2_X1 U761 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X1 U762 ( .A(G125), .B(n709), .ZN(G27) );
  XOR2_X1 U763 ( .A(G134), .B(n710), .Z(G36) );
  XOR2_X1 U764 ( .A(n711), .B(KEYINPUT124), .Z(n713) );
  NAND2_X1 U765 ( .A1(n713), .A2(n712), .ZN(n722) );
  NAND2_X1 U766 ( .A1(G953), .A2(G224), .ZN(n714) );
  XOR2_X1 U767 ( .A(KEYINPUT61), .B(n714), .Z(n715) );
  NOR2_X1 U768 ( .A1(n716), .A2(n715), .ZN(n720) );
  NAND2_X1 U769 ( .A1(n717), .A2(n725), .ZN(n718) );
  XNOR2_X1 U770 ( .A(n718), .B(KEYINPUT123), .ZN(n719) );
  NOR2_X1 U771 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U772 ( .A(n722), .B(n721), .ZN(G69) );
  XNOR2_X1 U773 ( .A(n724), .B(n723), .ZN(n727) );
  XOR2_X1 U774 ( .A(n645), .B(n727), .Z(n726) );
  NAND2_X1 U775 ( .A1(n726), .A2(n725), .ZN(n732) );
  XNOR2_X1 U776 ( .A(G227), .B(n727), .ZN(n728) );
  NAND2_X1 U777 ( .A1(n728), .A2(G900), .ZN(n729) );
  NAND2_X1 U778 ( .A1(G953), .A2(n729), .ZN(n730) );
  XOR2_X1 U779 ( .A(KEYINPUT125), .B(n730), .Z(n731) );
  NAND2_X1 U780 ( .A1(n732), .A2(n731), .ZN(G72) );
  XOR2_X1 U781 ( .A(G131), .B(n733), .Z(G33) );
  XNOR2_X1 U782 ( .A(G137), .B(KEYINPUT127), .ZN(n735) );
  XNOR2_X1 U783 ( .A(n735), .B(n734), .ZN(G39) );
endmodule

