//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  INV_X1    g000(.A(G107), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(KEYINPUT83), .A3(G104), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n190));
  NAND4_X1  g004(.A1(new_n190), .A2(new_n187), .A3(KEYINPUT83), .A4(G104), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n187), .A2(G104), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n189), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT4), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G101), .ZN(new_n196));
  INV_X1    g010(.A(G116), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT70), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT70), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G116), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n198), .A2(new_n200), .A3(G119), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT69), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n202), .B1(new_n197), .B2(G119), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n197), .A2(G119), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT69), .ZN(new_n205));
  AND3_X1   g019(.A1(new_n201), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  XOR2_X1   g020(.A(KEYINPUT2), .B(G113), .Z(new_n207));
  AND2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n206), .A2(new_n207), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n196), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT85), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n194), .A2(KEYINPUT84), .A3(G101), .ZN(new_n212));
  INV_X1    g026(.A(G101), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n189), .A2(new_n193), .A3(new_n213), .A4(new_n191), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(KEYINPUT4), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT84), .B1(new_n194), .B2(G101), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n211), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n216), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n214), .A2(KEYINPUT4), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT85), .A4(new_n212), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n210), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(G110), .B(G122), .ZN(new_n223));
  INV_X1    g037(.A(G104), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(G107), .ZN(new_n225));
  OAI21_X1  g039(.A(G101), .B1(new_n225), .B2(new_n192), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n214), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT5), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n204), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n201), .A2(new_n205), .A3(new_n203), .ZN(new_n231));
  OAI211_X1 g045(.A(G113), .B(new_n230), .C1(new_n231), .C2(new_n229), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n206), .A2(new_n207), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n228), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT89), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT89), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n228), .A2(new_n232), .A3(new_n236), .A4(new_n233), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n222), .A2(new_n223), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n223), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n241), .B1(new_n221), .B2(new_n238), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(new_n242), .A3(KEYINPUT6), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT6), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n244), .B(new_n241), .C1(new_n221), .C2(new_n238), .ZN(new_n245));
  INV_X1    g059(.A(G146), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G143), .ZN(new_n247));
  INV_X1    g061(.A(G143), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G146), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  NOR2_X1   g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT64), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n250), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n247), .A2(new_n249), .A3(new_n251), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n254), .B1(new_n250), .B2(new_n253), .ZN(new_n258));
  OAI21_X1  g072(.A(G125), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n247), .A2(KEYINPUT1), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n250), .A2(new_n260), .A3(G128), .ZN(new_n261));
  INV_X1    g075(.A(G128), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n247), .B(new_n249), .C1(KEYINPUT1), .C2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G125), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT90), .B(G224), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n268), .A2(G953), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n267), .B(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n243), .A2(new_n245), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n267), .B1(KEYINPUT91), .B2(KEYINPUT7), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT7), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n272), .B1(new_n273), .B2(new_n269), .ZN(new_n274));
  OAI221_X1 g088(.A(KEYINPUT7), .B1(G953), .B2(new_n268), .C1(new_n267), .C2(KEYINPUT91), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n232), .A2(new_n233), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n227), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n234), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n223), .B(KEYINPUT8), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n274), .A2(new_n275), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(G902), .B1(new_n280), .B2(new_n240), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n271), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(G210), .B1(G237), .B2(G902), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT92), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n271), .A2(new_n281), .A3(new_n283), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n287), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT92), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G469), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  XNOR2_X1  g107(.A(G110), .B(G140), .ZN(new_n294));
  INV_X1    g108(.A(G227), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(G953), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n294), .B(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n214), .A2(new_n261), .A3(new_n263), .A4(new_n226), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT10), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n299), .B(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n217), .A2(new_n220), .ZN(new_n302));
  INV_X1    g116(.A(new_n257), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n250), .A2(new_n253), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT64), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n303), .A2(new_n305), .A3(new_n196), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n301), .B1(new_n302), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT11), .ZN(new_n309));
  INV_X1    g123(.A(G134), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n309), .B1(new_n310), .B2(G137), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(G137), .ZN(new_n312));
  INV_X1    g126(.A(G137), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(KEYINPUT11), .A3(G134), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n311), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G131), .ZN(new_n316));
  INV_X1    g130(.A(G131), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n311), .A2(new_n314), .A3(new_n317), .A4(new_n312), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n316), .A2(KEYINPUT66), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT66), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n315), .A2(new_n320), .A3(G131), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT87), .B1(new_n308), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT87), .ZN(new_n324));
  INV_X1    g138(.A(new_n322), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n306), .B1(new_n217), .B2(new_n220), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n324), .B(new_n325), .C1(new_n326), .C2(new_n301), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n302), .A2(new_n307), .ZN(new_n329));
  INV_X1    g143(.A(new_n301), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n322), .B(KEYINPUT86), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n298), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n297), .B1(new_n308), .B2(new_n331), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n227), .A2(new_n264), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n299), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n325), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT12), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n337), .B(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n292), .B(new_n293), .C1(new_n333), .C2(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n298), .B1(new_n332), .B2(new_n339), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n342), .B1(new_n328), .B2(new_n334), .ZN(new_n343));
  OAI21_X1  g157(.A(G469), .B1(new_n343), .B2(G902), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT9), .B(G234), .ZN(new_n346));
  OAI21_X1  g160(.A(G221), .B1(new_n346), .B2(G902), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n347), .B(KEYINPUT82), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(G214), .B1(G237), .B2(G902), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(KEYINPUT88), .ZN(new_n352));
  NOR3_X1   g166(.A1(new_n291), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G478), .ZN(new_n354));
  OR2_X1    g168(.A1(new_n354), .A2(KEYINPUT15), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n262), .A2(G143), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n248), .A2(G128), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(G134), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n198), .A2(new_n200), .A3(G122), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n197), .A2(G122), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n360), .A2(new_n187), .A3(new_n362), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n363), .A2(KEYINPUT97), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n363), .A2(KEYINPUT97), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n359), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n360), .B1(KEYINPUT14), .B2(new_n361), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n367), .B(KEYINPUT98), .C1(KEYINPUT14), .C2(new_n360), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n360), .A2(KEYINPUT98), .A3(KEYINPUT14), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(new_n187), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n368), .A2(new_n370), .A3(KEYINPUT99), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT99), .B1(new_n368), .B2(new_n370), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n366), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n248), .A2(G128), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT13), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n374), .B1(new_n357), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT94), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n377), .B1(new_n356), .B2(KEYINPUT13), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n377), .B(new_n374), .C1(new_n357), .C2(new_n375), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G134), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT95), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n376), .A2(new_n378), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT95), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n383), .A2(new_n384), .A3(G134), .A4(new_n380), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n360), .A2(new_n362), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G107), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n388), .A2(new_n363), .B1(new_n310), .B2(new_n358), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n386), .A2(KEYINPUT96), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT96), .B1(new_n386), .B2(new_n389), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n373), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G217), .ZN(new_n393));
  NOR3_X1   g207(.A1(new_n346), .A2(new_n393), .A3(G953), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n373), .B(new_n394), .C1(new_n390), .C2(new_n391), .ZN(new_n397));
  AOI21_X1  g211(.A(G902), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT100), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI211_X1 g214(.A(KEYINPUT100), .B(G902), .C1(new_n396), .C2(new_n397), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n355), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OR2_X1    g216(.A1(new_n401), .A2(new_n355), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(G113), .B(G122), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(new_n224), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(G237), .A2(G953), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G214), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n248), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(G143), .A3(G214), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AND2_X1   g226(.A1(KEYINPUT18), .A2(G131), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n412), .B(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n265), .A2(G140), .ZN(new_n415));
  INV_X1    g229(.A(G140), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G125), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT77), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT77), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n415), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n421), .A3(new_n246), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT78), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n423), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n415), .A2(new_n417), .A3(KEYINPUT75), .ZN(new_n428));
  OR3_X1    g242(.A1(new_n416), .A2(KEYINPUT75), .A3(G125), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT93), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT93), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n428), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n431), .A2(G146), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n414), .B1(new_n427), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n412), .A2(G131), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT17), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n410), .A2(new_n317), .A3(new_n411), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT16), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n440), .B1(new_n428), .B2(new_n429), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n416), .A3(G125), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(KEYINPUT76), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n442), .A2(G146), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT76), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n443), .B(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n246), .B1(new_n447), .B2(new_n441), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n412), .A2(KEYINPUT17), .A3(G131), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n439), .A2(new_n445), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n407), .B1(new_n435), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n426), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n434), .B1(new_n453), .B2(new_n424), .ZN(new_n454));
  INV_X1    g268(.A(new_n414), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(new_n406), .A3(new_n450), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n293), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G475), .ZN(new_n460));
  INV_X1    g274(.A(G953), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n461), .A2(G952), .ZN(new_n462));
  INV_X1    g276(.A(G234), .ZN(new_n463));
  INV_X1    g277(.A(G237), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI211_X1 g280(.A(new_n293), .B(new_n461), .C1(G234), .C2(G237), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(G898), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n431), .A2(KEYINPUT19), .A3(new_n433), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT19), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n419), .A2(new_n421), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n471), .A2(new_n246), .A3(new_n473), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n447), .A2(new_n441), .A3(new_n246), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(new_n436), .B2(new_n438), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n474), .A2(new_n476), .B1(new_n454), .B2(new_n455), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n457), .B1(new_n477), .B2(new_n406), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT20), .ZN(new_n479));
  NOR2_X1   g293(.A1(G475), .A2(G902), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n479), .B1(new_n478), .B2(new_n480), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n460), .B(new_n470), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n404), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n264), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT67), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n486), .B1(new_n310), .B2(G137), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n313), .A2(KEYINPUT67), .A3(G134), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n488), .A3(new_n312), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT68), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n489), .A2(new_n490), .A3(G131), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n490), .B1(new_n489), .B2(G131), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n485), .B(new_n318), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT65), .B1(new_n257), .B2(new_n258), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT65), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n305), .A2(new_n255), .A3(new_n495), .A4(new_n256), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n493), .B1(new_n497), .B2(new_n322), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT30), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n231), .B(new_n207), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n303), .A2(new_n319), .A3(new_n321), .A4(new_n305), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n493), .A2(new_n503), .A3(KEYINPUT30), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n493), .A2(new_n503), .A3(new_n501), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n408), .A2(G210), .ZN(new_n507));
  XOR2_X1   g321(.A(new_n507), .B(KEYINPUT27), .Z(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT26), .B(G101), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n505), .A2(new_n506), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT31), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n498), .A2(new_n502), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT28), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n506), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n493), .A2(new_n503), .A3(KEYINPUT28), .A4(new_n501), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n510), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT31), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n505), .A2(new_n520), .A3(new_n506), .A4(new_n511), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n513), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(G472), .A2(G902), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT71), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT32), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT71), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n522), .A2(new_n527), .A3(new_n523), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT72), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n506), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n493), .A2(new_n503), .A3(KEYINPUT72), .A4(new_n501), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n493), .A2(new_n503), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n502), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT28), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT29), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n510), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n536), .A2(new_n516), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n537), .B1(new_n518), .B2(new_n510), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n511), .B1(new_n505), .B2(new_n506), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n539), .B(new_n293), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G472), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT73), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT73), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n542), .A2(new_n545), .A3(G472), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n522), .A2(KEYINPUT32), .A3(new_n523), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n529), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n445), .A2(new_n448), .ZN(new_n550));
  XNOR2_X1  g364(.A(G119), .B(G128), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT74), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XOR2_X1   g367(.A(KEYINPUT24), .B(G110), .Z(new_n554));
  INV_X1    g368(.A(KEYINPUT23), .ZN(new_n555));
  INV_X1    g369(.A(G119), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n555), .B1(new_n556), .B2(G128), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n262), .A2(KEYINPUT23), .A3(G119), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n557), .B(new_n558), .C1(G119), .C2(new_n262), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n553), .A2(new_n554), .B1(G110), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n550), .A2(new_n560), .ZN(new_n561));
  OAI22_X1  g375(.A1(new_n553), .A2(new_n554), .B1(G110), .B2(new_n559), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n562), .B(new_n445), .C1(new_n453), .C2(new_n424), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT22), .B(G137), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n461), .A2(G221), .A3(G234), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n565), .B(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n561), .A2(new_n563), .A3(new_n567), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n293), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT25), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT25), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n569), .A2(new_n573), .A3(new_n293), .A4(new_n570), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n393), .B1(G234), .B2(new_n293), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT79), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n569), .A2(new_n570), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT80), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n575), .A2(G902), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n572), .A2(KEYINPUT79), .A3(new_n574), .A4(new_n575), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n579), .A2(new_n581), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT80), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n578), .A2(new_n582), .A3(new_n583), .A4(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n549), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(KEYINPUT81), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT81), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n549), .B2(new_n587), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n353), .B(new_n484), .C1(new_n589), .C2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(G101), .ZN(G3));
  AND2_X1   g407(.A1(new_n525), .A2(new_n528), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n522), .A2(new_n293), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT101), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n522), .A2(KEYINPUT101), .A3(new_n293), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n597), .A2(G472), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n594), .A2(new_n587), .A3(new_n599), .ZN(new_n600));
  OR2_X1    g414(.A1(new_n600), .A2(new_n350), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n396), .A2(new_n397), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT33), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n396), .A2(new_n604), .A3(new_n397), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n603), .A2(G478), .A3(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n354), .A2(new_n293), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n607), .B1(new_n398), .B2(new_n354), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(G475), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n458), .B2(new_n293), .ZN(new_n611));
  INV_X1    g425(.A(new_n482), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n470), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n283), .B1(new_n271), .B2(new_n281), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n351), .B1(new_n289), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n601), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT34), .B(G104), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  OAI21_X1  g437(.A(new_n612), .B1(new_n481), .B2(KEYINPUT102), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT102), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n482), .A2(new_n625), .A3(new_n613), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n611), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n404), .A2(new_n627), .A3(new_n470), .ZN(new_n628));
  OR3_X1    g442(.A1(new_n628), .A2(KEYINPUT103), .A3(new_n618), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT103), .B1(new_n628), .B2(new_n618), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n601), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(KEYINPUT35), .B(G107), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  NOR2_X1   g447(.A1(new_n568), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT104), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(new_n564), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n581), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n578), .A2(new_n583), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n483), .ZN(new_n639));
  AND4_X1   g453(.A1(new_n402), .A2(new_n638), .A3(new_n639), .A4(new_n403), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n640), .A2(new_n594), .A3(new_n599), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n353), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT37), .B(G110), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G12));
  OAI211_X1 g458(.A(new_n638), .B(new_n351), .C1(new_n289), .C2(new_n617), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n350), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(G900), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n466), .B1(new_n467), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n404), .A2(new_n627), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n646), .A2(new_n549), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G128), .ZN(G30));
  XNOR2_X1  g467(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n291), .B(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n460), .B1(new_n481), .B2(new_n482), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n404), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n351), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n658), .A2(new_n659), .A3(new_n638), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n510), .B1(new_n505), .B2(new_n506), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n293), .B1(new_n535), .B2(new_n511), .ZN(new_n662));
  OAI21_X1  g476(.A(G472), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n529), .A2(new_n548), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(KEYINPUT106), .B1(new_n656), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n655), .A2(new_n667), .A3(new_n664), .A4(new_n660), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n648), .B(KEYINPUT39), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n350), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT40), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n666), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n666), .A2(KEYINPUT107), .A3(new_n668), .A4(new_n671), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n248), .ZN(G45));
  AND4_X1   g491(.A1(new_n657), .A2(new_n606), .A3(new_n608), .A4(new_n649), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n646), .A2(new_n549), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT108), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n646), .A2(new_n549), .A3(new_n681), .A4(new_n678), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G146), .ZN(G48));
  OAI21_X1  g498(.A(new_n293), .B1(new_n333), .B2(new_n340), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G469), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n341), .ZN(new_n687));
  INV_X1    g501(.A(new_n347), .ZN(new_n688));
  OAI21_X1  g502(.A(KEYINPUT109), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT109), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n686), .A2(new_n690), .A3(new_n347), .A4(new_n341), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n689), .A2(new_n549), .A3(new_n587), .A4(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n620), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT41), .B(G113), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G15));
  INV_X1    g509(.A(new_n692), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n629), .A2(new_n630), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G116), .ZN(G18));
  AOI21_X1  g513(.A(new_n659), .B1(new_n285), .B2(new_n287), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n689), .A2(new_n700), .A3(new_n691), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n549), .A2(new_n640), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  NAND2_X1  g519(.A1(new_n689), .A2(new_n691), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT111), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n708), .B1(new_n658), .B2(new_n618), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n614), .B1(new_n402), .B2(new_n403), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n700), .A2(new_n710), .A3(KEYINPUT111), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n586), .A2(KEYINPUT110), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n585), .A2(new_n582), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT110), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n714), .A2(new_n715), .A3(new_n578), .A4(new_n583), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n595), .A2(G472), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n536), .A2(new_n516), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n513), .B(new_n521), .C1(new_n719), .C2(new_n511), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n523), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n469), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n707), .A2(new_n712), .A3(new_n724), .ZN(new_n725));
  XOR2_X1   g539(.A(KEYINPUT112), .B(G122), .Z(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G24));
  AND4_X1   g541(.A1(new_n638), .A2(new_n678), .A3(new_n721), .A4(new_n718), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n689), .A2(new_n728), .A3(new_n700), .A4(new_n691), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G125), .ZN(G27));
  INV_X1    g544(.A(new_n588), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT42), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n659), .B1(new_n288), .B2(new_n290), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n688), .B1(new_n341), .B2(new_n344), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n731), .A2(new_n732), .A3(new_n735), .A4(new_n678), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n733), .A2(new_n678), .A3(new_n734), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n524), .A2(new_n526), .ZN(new_n739));
  INV_X1    g553(.A(new_n546), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n545), .B1(new_n542), .B2(G472), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n739), .B(new_n548), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n738), .B1(new_n742), .B2(new_n717), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n742), .A2(new_n717), .A3(new_n738), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n737), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n736), .B1(new_n746), .B2(new_n732), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n317), .ZN(G33));
  NAND3_X1  g562(.A1(new_n731), .A2(new_n651), .A3(new_n735), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G134), .ZN(G36));
  AND2_X1   g564(.A1(new_n343), .A2(KEYINPUT45), .ZN(new_n751));
  OAI21_X1  g565(.A(G469), .B1(new_n343), .B2(KEYINPUT45), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(G469), .A2(G902), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT46), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n753), .A2(KEYINPUT46), .A3(new_n754), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n341), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n347), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n669), .ZN(new_n761));
  INV_X1    g575(.A(new_n733), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n614), .A2(new_n606), .A3(new_n608), .ZN(new_n763));
  XOR2_X1   g577(.A(new_n763), .B(KEYINPUT43), .Z(new_n764));
  NAND2_X1  g578(.A1(new_n594), .A2(new_n599), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n765), .A3(new_n638), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n762), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n761), .B(new_n768), .C1(new_n767), .C2(new_n766), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G137), .ZN(G39));
  INV_X1    g584(.A(new_n760), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT47), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n771), .B1(KEYINPUT114), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n678), .A2(new_n586), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n762), .A2(new_n549), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(KEYINPUT114), .B(KEYINPUT47), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n773), .B(new_n775), .C1(new_n771), .C2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G140), .ZN(G42));
  NOR3_X1   g592(.A1(new_n664), .A2(new_n586), .A3(new_n465), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n707), .A2(new_n779), .A3(new_n733), .ZN(new_n780));
  AOI211_X1 g594(.A(new_n657), .B(new_n780), .C1(new_n606), .C2(new_n608), .ZN(new_n781));
  XOR2_X1   g595(.A(new_n781), .B(KEYINPUT122), .Z(new_n782));
  OAI21_X1  g596(.A(new_n773), .B1(new_n771), .B2(new_n776), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n783), .B1(new_n349), .B2(new_n687), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n764), .A2(new_n466), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n723), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n733), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT121), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n785), .A2(new_n706), .A3(new_n762), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n790), .A2(new_n638), .A3(new_n722), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n786), .A2(new_n659), .A3(new_n656), .A4(new_n707), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT50), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n792), .A2(new_n793), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n782), .A2(new_n789), .A3(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n782), .A2(KEYINPUT51), .A3(new_n789), .A4(new_n796), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n742), .A2(new_n717), .A3(new_n738), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(new_n743), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n790), .A2(new_n803), .ZN(new_n804));
  XOR2_X1   g618(.A(new_n804), .B(KEYINPUT48), .Z(new_n805));
  NAND2_X1  g619(.A1(new_n786), .A2(new_n701), .ZN(new_n806));
  INV_X1    g620(.A(new_n615), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n806), .B(new_n462), .C1(new_n780), .C2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n799), .A2(new_n800), .A3(new_n809), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n696), .A2(new_n697), .B1(new_n701), .B2(new_n703), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n600), .A2(new_n616), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n696), .A2(new_n619), .B1(new_n353), .B2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n811), .A2(new_n813), .A3(new_n592), .A4(new_n725), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT42), .B1(new_n802), .B2(new_n737), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n401), .A2(new_n355), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n398), .B(new_n399), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n816), .B1(new_n817), .B2(new_n355), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n818), .A2(new_n627), .A3(new_n638), .A4(new_n649), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n350), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n820), .A2(new_n549), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n728), .A2(new_n734), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n733), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n815), .A2(new_n823), .A3(new_n736), .A4(new_n749), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT115), .B1(new_n404), .B2(new_n614), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n827));
  AOI211_X1 g641(.A(new_n827), .B(new_n657), .C1(new_n402), .C2(new_n403), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n470), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(new_n600), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n825), .B(new_n353), .C1(new_n830), .C2(new_n641), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n827), .B1(new_n818), .B2(new_n657), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n404), .A2(KEYINPUT115), .A3(new_n614), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n469), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n594), .A2(new_n587), .A3(new_n599), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n353), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n642), .A3(KEYINPUT116), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n831), .A2(new_n837), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n814), .A2(new_n824), .A3(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n729), .A2(new_n652), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT117), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n638), .A2(new_n648), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n734), .A2(new_n843), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n700), .A2(new_n710), .A3(KEYINPUT111), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT111), .B1(new_n700), .B2(new_n710), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n664), .B(new_n844), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n712), .A2(KEYINPUT118), .A3(new_n664), .A4(new_n844), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n842), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n729), .A2(new_n652), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT117), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n841), .A2(new_n851), .A3(new_n683), .A4(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(KEYINPUT119), .B(KEYINPUT52), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n849), .A2(new_n850), .B1(new_n680), .B2(new_n682), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n856), .B1(new_n857), .B2(new_n840), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n855), .B1(new_n858), .B2(KEYINPUT120), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n860));
  AOI211_X1 g674(.A(new_n860), .B(new_n856), .C1(new_n857), .C2(new_n840), .ZN(new_n861));
  OAI211_X1 g675(.A(KEYINPUT53), .B(new_n839), .C1(new_n859), .C2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n857), .A2(KEYINPUT52), .A3(new_n840), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT52), .B1(new_n857), .B2(new_n840), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI22_X1  g680(.A1(new_n820), .A2(new_n549), .B1(new_n728), .B2(new_n734), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n749), .B1(new_n762), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n747), .A2(new_n868), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n813), .A2(new_n592), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n831), .A2(new_n837), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n698), .A2(new_n704), .A3(new_n725), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n869), .A2(new_n870), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n863), .B1(new_n866), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n862), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n866), .A2(new_n873), .A3(new_n863), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n839), .B1(new_n859), .B2(new_n861), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n877), .B1(new_n863), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n876), .B1(new_n879), .B2(new_n875), .ZN(new_n880));
  OAI22_X1  g694(.A1(new_n810), .A2(new_n880), .B1(G952), .B2(G953), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n687), .A2(KEYINPUT49), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n763), .A2(new_n348), .A3(new_n352), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n882), .A2(new_n717), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n687), .A2(KEYINPUT49), .ZN(new_n885));
  OR3_X1    g699(.A1(new_n884), .A2(new_n664), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n881), .B1(new_n655), .B2(new_n886), .ZN(G75));
  AOI21_X1  g701(.A(new_n293), .B1(new_n862), .B2(new_n874), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(G210), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT56), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n243), .A2(new_n245), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT123), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n270), .B(KEYINPUT55), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n893), .B(new_n894), .Z(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n461), .A2(G952), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n895), .B1(new_n889), .B2(new_n890), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(G51));
  NAND2_X1  g714(.A1(new_n862), .A2(new_n874), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(new_n875), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n754), .B(KEYINPUT57), .ZN(new_n903));
  OAI22_X1  g717(.A1(new_n902), .A2(new_n903), .B1(new_n333), .B2(new_n340), .ZN(new_n904));
  INV_X1    g718(.A(new_n753), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n888), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n898), .B1(new_n904), .B2(new_n906), .ZN(G54));
  AND2_X1   g721(.A1(KEYINPUT58), .A2(G475), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n888), .A2(new_n478), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n478), .B1(new_n888), .B2(new_n908), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n909), .A2(new_n910), .A3(new_n898), .ZN(G60));
  INV_X1    g725(.A(new_n898), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n603), .A2(new_n605), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n607), .B(KEYINPUT59), .Z(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n912), .B1(new_n902), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n913), .B1(new_n880), .B2(new_n914), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(G63));
  NAND2_X1  g732(.A1(G217), .A2(G902), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT60), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n920), .B1(new_n862), .B2(new_n874), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n912), .B1(new_n921), .B2(new_n579), .ZN(new_n922));
  INV_X1    g736(.A(new_n920), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n901), .A2(new_n636), .A3(new_n923), .ZN(new_n924));
  OAI211_X1 g738(.A(KEYINPUT124), .B(KEYINPUT61), .C1(new_n922), .C2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n901), .A2(new_n636), .A3(new_n923), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n927), .B(new_n912), .C1(new_n579), .C2(new_n921), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT61), .B1(new_n928), .B2(KEYINPUT124), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n926), .A2(new_n929), .ZN(G66));
  NOR2_X1   g744(.A1(new_n268), .A2(new_n468), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n931), .A2(new_n461), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n870), .A2(new_n872), .A3(new_n871), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n933), .B2(new_n461), .ZN(new_n934));
  INV_X1    g748(.A(G898), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n893), .B1(new_n935), .B2(G953), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n934), .B(new_n936), .ZN(G69));
  NAND2_X1  g751(.A1(new_n500), .A2(new_n504), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n471), .A2(new_n473), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT125), .Z(new_n940));
  XNOR2_X1  g754(.A(new_n938), .B(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n589), .A2(new_n591), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n832), .A2(new_n807), .A3(new_n833), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n943), .A2(new_n670), .A3(new_n733), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n777), .B(new_n769), .C1(new_n942), .C2(new_n944), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n841), .A2(new_n683), .A3(new_n854), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n946), .A2(new_n674), .A3(new_n675), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n946), .A2(new_n674), .A3(KEYINPUT62), .A4(new_n675), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n945), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n941), .B1(new_n951), .B2(G953), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(KEYINPUT126), .ZN(new_n953));
  INV_X1    g767(.A(new_n941), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n761), .A2(new_n712), .A3(new_n803), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n769), .A2(new_n955), .A3(new_n749), .ZN(new_n956));
  INV_X1    g770(.A(new_n747), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n956), .A2(new_n957), .A3(new_n777), .A4(new_n946), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n958), .A2(new_n461), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n461), .A2(G900), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n954), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n962), .B(new_n941), .C1(new_n951), .C2(G953), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n953), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(G953), .B1(new_n295), .B2(new_n647), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT127), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n953), .A2(new_n961), .A3(new_n966), .A4(new_n963), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(G72));
  INV_X1    g784(.A(new_n512), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n971), .A2(new_n541), .ZN(new_n972));
  NAND2_X1  g786(.A1(G472), .A2(G902), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT63), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n898), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n505), .A2(new_n506), .A3(new_n510), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n958), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n661), .B2(new_n951), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n975), .B1(new_n978), .B2(new_n933), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n879), .A2(new_n974), .A3(new_n972), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(G57));
endmodule


