//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1281, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1340, new_n1341,
    new_n1342;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(KEYINPUT64), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g0012(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n204), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n209), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT65), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT66), .B(G244), .ZN(new_n221));
  AND2_X1   g0021(.A1(new_n221), .A2(G77), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G116), .A2(G270), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n223), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n206), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n220), .A2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G68), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT67), .ZN(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  XNOR2_X1  g0047(.A(KEYINPUT8), .B(G58), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT69), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G20), .ZN(new_n252));
  INV_X1    g0052(.A(G58), .ZN(new_n253));
  OR3_X1    g0053(.A1(new_n249), .A2(new_n253), .A3(KEYINPUT8), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n250), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G50), .ZN(new_n256));
  INV_X1    g0056(.A(G68), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(new_n253), .A3(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n258), .A2(G20), .B1(G150), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n255), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n212), .A2(new_n213), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT70), .ZN(new_n265));
  OR2_X1    g0065(.A1(KEYINPUT68), .A2(G1), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT68), .A2(G1), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n266), .A2(G13), .A3(G20), .A4(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(G50), .ZN(new_n269));
  AND3_X1   g0069(.A1(new_n212), .A2(new_n213), .A3(new_n262), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT68), .B(G1), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n270), .B1(new_n204), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n269), .B1(new_n273), .B2(G50), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n265), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n264), .A2(KEYINPUT70), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n251), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  AOI21_X1  g0080(.A(G1698), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G222), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(new_n280), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G223), .A3(G1698), .ZN(new_n284));
  INV_X1    g0084(.A(G77), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n282), .B(new_n284), .C1(new_n285), .C2(new_n283), .ZN(new_n286));
  AND2_X1   g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n287), .B1(new_n212), .B2(new_n213), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(G274), .B1(new_n287), .B2(new_n210), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G41), .A2(G45), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n290), .A2(G1), .A3(new_n291), .ZN(new_n292));
  AND2_X1   g0092(.A1(G1), .A2(G13), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G41), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n295), .B1(new_n271), .B2(new_n291), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n292), .B1(new_n297), .B2(G226), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n289), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n299), .A2(G169), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n277), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G274), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(new_n293), .B2(new_n294), .ZN(new_n305));
  INV_X1    g0105(.A(new_n291), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n305), .A2(new_n203), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G238), .ZN(new_n308));
  NAND2_X1  g0108(.A1(G33), .A2(G97), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(G226), .A2(G1698), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n232), .B2(G1698), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n310), .B1(new_n312), .B2(new_n283), .ZN(new_n313));
  INV_X1    g0113(.A(new_n288), .ZN(new_n314));
  OAI221_X1 g0114(.A(new_n307), .B1(new_n296), .B2(new_n308), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT13), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n312), .A2(new_n283), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n309), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n292), .B1(new_n318), .B2(new_n288), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT13), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n297), .A2(G238), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G200), .ZN(new_n324));
  INV_X1    g0124(.A(G190), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n252), .A2(G77), .ZN(new_n327));
  INV_X1    g0127(.A(new_n259), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n327), .B1(new_n204), .B2(G68), .C1(new_n256), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n263), .ZN(new_n330));
  XOR2_X1   g0130(.A(new_n330), .B(KEYINPUT11), .Z(new_n331));
  NOR2_X1   g0131(.A1(new_n268), .A2(G68), .ZN(new_n332));
  XOR2_X1   g0132(.A(new_n332), .B(KEYINPUT12), .Z(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n257), .B2(new_n272), .ZN(new_n334));
  NOR3_X1   g0134(.A1(new_n326), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n303), .B1(new_n324), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT15), .B(G87), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n252), .ZN(new_n339));
  XOR2_X1   g0139(.A(new_n339), .B(KEYINPUT74), .Z(new_n340));
  INV_X1    g0140(.A(KEYINPUT73), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n248), .B1(new_n341), .B2(new_n328), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n341), .B2(new_n328), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n204), .B2(new_n285), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n263), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n268), .A2(G77), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(new_n273), .B2(G77), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n221), .B(new_n295), .C1(new_n271), .C2(new_n291), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n307), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT71), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT71), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n350), .A2(new_n307), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G1698), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n232), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n308), .A2(G1698), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n356), .A2(new_n357), .B1(new_n279), .B2(new_n280), .ZN(new_n358));
  AND2_X1   g0158(.A1(KEYINPUT3), .A2(G33), .ZN(new_n359));
  NOR2_X1   g0159(.A1(KEYINPUT3), .A2(G33), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n359), .A2(new_n360), .A3(G107), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n288), .ZN(new_n363));
  AND4_X1   g0163(.A1(KEYINPUT72), .A2(new_n352), .A3(new_n354), .A4(new_n363), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n351), .A2(KEYINPUT71), .B1(new_n362), .B2(new_n288), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT72), .B1(new_n365), .B2(new_n354), .ZN(new_n366));
  OAI21_X1  g0166(.A(G190), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n352), .A2(new_n354), .A3(new_n363), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT72), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n365), .A2(KEYINPUT72), .A3(new_n354), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(G200), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n349), .A2(new_n367), .A3(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n300), .B1(new_n364), .B2(new_n366), .ZN(new_n374));
  INV_X1    g0174(.A(G169), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n370), .A2(new_n375), .A3(new_n371), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n348), .A3(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n331), .A2(new_n334), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT14), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n323), .A2(new_n380), .A3(G169), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n316), .A2(new_n322), .A3(G179), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n380), .B1(new_n323), .B2(G169), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n379), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n336), .A2(new_n373), .A3(new_n377), .A4(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT9), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n275), .B2(new_n276), .ZN(new_n388));
  INV_X1    g0188(.A(G200), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n389), .B1(new_n289), .B2(new_n298), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(G190), .B2(new_n299), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n264), .A2(KEYINPUT70), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n392), .A2(KEYINPUT9), .A3(new_n265), .A4(new_n274), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT10), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT10), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n388), .A2(new_n391), .A3(new_n393), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n259), .A2(G159), .ZN(new_n400));
  XNOR2_X1  g0200(.A(G58), .B(G68), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT75), .B1(new_n401), .B2(G20), .ZN(new_n402));
  AND2_X1   g0202(.A1(G58), .A2(G68), .ZN(new_n403));
  NOR2_X1   g0203(.A1(G58), .A2(G68), .ZN(new_n404));
  OAI211_X1 g0204(.A(KEYINPUT75), .B(G20), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n400), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n279), .A2(new_n204), .A3(new_n280), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT7), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n279), .A2(KEYINPUT7), .A3(new_n204), .A4(new_n280), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n257), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n399), .B1(new_n407), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n359), .A2(new_n360), .ZN(new_n414));
  AOI21_X1  g0214(.A(KEYINPUT7), .B1(new_n414), .B2(new_n204), .ZN(new_n415));
  INV_X1    g0215(.A(new_n411), .ZN(new_n416));
  OAI21_X1  g0216(.A(G68), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(G20), .B1(new_n403), .B2(new_n404), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT75), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n420), .A2(new_n405), .B1(G159), .B2(new_n259), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n417), .A2(new_n421), .A3(KEYINPUT16), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n413), .A2(new_n263), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n250), .A2(new_n254), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n272), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n268), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n307), .B1(new_n296), .B2(new_n232), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n283), .A2(G226), .A3(G1698), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n283), .A2(G223), .A3(new_n355), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G33), .A2(G87), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT76), .ZN(new_n435));
  XNOR2_X1  g0235(.A(new_n434), .B(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n432), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n288), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n431), .A2(new_n438), .A3(G179), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n430), .B1(new_n288), .B2(new_n437), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n439), .B1(new_n375), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n429), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT18), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT18), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n429), .A2(new_n444), .A3(new_n441), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n431), .A2(new_n438), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G200), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n440), .A2(G190), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n423), .A2(new_n448), .A3(new_n449), .A4(new_n428), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT17), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n431), .A2(new_n438), .A3(G190), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n389), .B1(new_n431), .B2(new_n438), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n455), .A2(KEYINPUT17), .A3(new_n423), .A4(new_n428), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n398), .A2(new_n446), .A3(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n386), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT79), .ZN(new_n461));
  AND2_X1   g0261(.A1(KEYINPUT4), .A2(G244), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n355), .B(new_n462), .C1(new_n359), .C2(new_n360), .ZN(new_n463));
  INV_X1    g0263(.A(G283), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n251), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(G244), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n467), .B1(new_n279), .B2(new_n280), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n463), .B(new_n466), .C1(new_n468), .C2(KEYINPUT4), .ZN(new_n469));
  OAI21_X1  g0269(.A(G250), .B1(new_n359), .B2(new_n360), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n355), .B1(new_n470), .B2(KEYINPUT4), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n461), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G250), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n473), .B1(new_n279), .B2(new_n280), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT4), .ZN(new_n475));
  OAI21_X1  g0275(.A(G1698), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n465), .B1(new_n281), .B2(new_n462), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n475), .B1(new_n414), .B2(new_n467), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT79), .A4(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n472), .A2(new_n479), .A3(new_n288), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT5), .ZN(new_n481));
  AOI21_X1  g0281(.A(G41), .B1(new_n481), .B2(KEYINPUT80), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT80), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT5), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n481), .A2(G41), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n266), .A2(new_n486), .A3(G45), .A4(new_n267), .ZN(new_n487));
  NOR3_X1   g0287(.A1(new_n485), .A2(new_n487), .A3(new_n290), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n287), .A2(new_n210), .ZN(new_n489));
  INV_X1    g0289(.A(G41), .ZN(new_n490));
  OAI21_X1  g0290(.A(G45), .B1(new_n490), .B2(KEYINPUT5), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n271), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n482), .A2(new_n484), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n489), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n488), .B1(G257), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n480), .A2(G190), .A3(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n271), .A2(new_n204), .ZN(new_n497));
  INV_X1    g0297(.A(G97), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n497), .A2(G13), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n266), .A2(G33), .A3(new_n267), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n270), .A2(new_n268), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n499), .B1(new_n501), .B2(new_n498), .ZN(new_n502));
  XOR2_X1   g0302(.A(G97), .B(G107), .Z(new_n503));
  XNOR2_X1  g0303(.A(KEYINPUT77), .B(KEYINPUT6), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n503), .A2(KEYINPUT78), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT6), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT77), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT77), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n498), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n507), .A2(new_n509), .A3(KEYINPUT78), .ZN(new_n512));
  XNOR2_X1  g0312(.A(G97), .B(G107), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n505), .A2(G20), .A3(new_n511), .A4(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(G107), .B1(new_n415), .B2(new_n416), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n259), .A2(G77), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n502), .B1(new_n518), .B2(new_n263), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n496), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n389), .B1(new_n480), .B2(new_n495), .ZN(new_n521));
  OAI21_X1  g0321(.A(KEYINPUT81), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n480), .A2(new_n495), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G200), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT81), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n524), .A2(new_n525), .A3(new_n519), .A4(new_n496), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n266), .A2(new_n267), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n528), .A2(new_n305), .A3(KEYINPUT83), .A4(G45), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT83), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n266), .A2(G45), .A3(new_n267), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(new_n290), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n489), .A2(new_n473), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n531), .ZN(new_n535));
  NOR2_X1   g0335(.A1(G238), .A2(G1698), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n536), .B1(new_n467), .B2(G1698), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n537), .A2(new_n283), .B1(G33), .B2(G116), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n535), .B1(new_n538), .B2(new_n314), .ZN(new_n539));
  OAI21_X1  g0339(.A(G200), .B1(new_n533), .B2(new_n539), .ZN(new_n540));
  NOR3_X1   g0340(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n541));
  AND2_X1   g0341(.A1(KEYINPUT84), .A2(KEYINPUT19), .ZN(new_n542));
  NOR2_X1   g0342(.A1(KEYINPUT84), .A2(KEYINPUT19), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n310), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n541), .B1(new_n544), .B2(new_n204), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n204), .B(G68), .C1(new_n359), .C2(new_n360), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n204), .A2(G33), .A3(G97), .ZN(new_n547));
  OR2_X1    g0347(.A1(KEYINPUT84), .A2(KEYINPUT19), .ZN(new_n548));
  NAND2_X1  g0348(.A1(KEYINPUT84), .A2(KEYINPUT19), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n263), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n497), .A2(G13), .A3(new_n337), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n270), .A2(G87), .A3(new_n268), .A4(new_n500), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n540), .A2(new_n555), .A3(KEYINPUT85), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT85), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G116), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n467), .A2(G1698), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(G238), .B2(G1698), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n558), .B1(new_n560), .B2(new_n414), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n561), .A2(new_n288), .B1(new_n534), .B2(new_n531), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n529), .A2(new_n532), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n389), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n557), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n562), .A2(G190), .A3(new_n563), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n556), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n562), .A2(new_n563), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n375), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n552), .B(new_n553), .C1(new_n337), .C2(new_n501), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n562), .A2(new_n300), .A3(new_n563), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT86), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT86), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n568), .A2(new_n576), .A3(new_n573), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n519), .B1(new_n523), .B2(new_n375), .ZN(new_n578));
  OAI21_X1  g0378(.A(KEYINPUT82), .B1(new_n523), .B2(G179), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT82), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n480), .A2(new_n495), .A3(new_n580), .A4(new_n300), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n527), .A2(new_n575), .A3(new_n577), .A4(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT23), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n204), .B2(G107), .ZN(new_n585));
  INV_X1    g0385(.A(G107), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(KEYINPUT23), .A3(G20), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n252), .A2(G116), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n204), .B(G87), .C1(new_n359), .C2(new_n360), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT22), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT22), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n283), .A2(new_n593), .A3(new_n204), .A4(G87), .ZN(new_n594));
  AOI211_X1 g0394(.A(KEYINPUT24), .B(new_n590), .C1(new_n592), .C2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT24), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n592), .A2(new_n594), .ZN(new_n597));
  INV_X1    g0397(.A(new_n590), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n263), .B1(new_n595), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n501), .A2(new_n586), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT25), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n268), .B2(G107), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n268), .A2(new_n602), .A3(G107), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT90), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(KEYINPUT90), .B(new_n602), .C1(new_n268), .C2(G107), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n601), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(G257), .B(G1698), .C1(new_n359), .C2(new_n360), .ZN(new_n609));
  OAI211_X1 g0409(.A(G250), .B(new_n355), .C1(new_n359), .C2(new_n360), .ZN(new_n610));
  INV_X1    g0410(.A(G294), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n609), .B(new_n610), .C1(new_n251), .C2(new_n611), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n494), .A2(G264), .B1(new_n612), .B2(new_n288), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n492), .A2(new_n305), .A3(new_n493), .ZN(new_n614));
  AOI21_X1  g0414(.A(G200), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n612), .A2(new_n288), .ZN(new_n616));
  OAI211_X1 g0416(.A(G264), .B(new_n295), .C1(new_n485), .C2(new_n487), .ZN(new_n617));
  AND4_X1   g0417(.A1(new_n325), .A2(new_n616), .A3(new_n614), .A4(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n600), .B(new_n608), .C1(new_n615), .C2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT92), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n616), .A2(new_n614), .A3(new_n617), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n389), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(G190), .B2(new_n622), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n624), .A2(KEYINPUT92), .A3(new_n600), .A4(new_n608), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT91), .ZN(new_n627));
  AOI21_X1  g0427(.A(G20), .B1(new_n279), .B2(new_n280), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n593), .B1(new_n628), .B2(G87), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n591), .A2(KEYINPUT22), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n598), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT24), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n597), .A2(new_n596), .A3(new_n598), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n270), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n606), .A2(new_n607), .ZN(new_n635));
  INV_X1    g0435(.A(new_n601), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n627), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n600), .A2(new_n608), .A3(KEYINPUT91), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n622), .A2(G169), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n300), .B2(new_n622), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n638), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n626), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(KEYINPUT87), .A2(G303), .ZN(new_n644));
  NOR2_X1   g0444(.A1(KEYINPUT87), .A2(G303), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n279), .B(new_n280), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  OAI211_X1 g0446(.A(G264), .B(G1698), .C1(new_n359), .C2(new_n360), .ZN(new_n647));
  OAI211_X1 g0447(.A(G257), .B(new_n355), .C1(new_n359), .C2(new_n360), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n288), .ZN(new_n650));
  OAI211_X1 g0450(.A(G270), .B(new_n295), .C1(new_n485), .C2(new_n487), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(new_n614), .A3(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n270), .A2(G116), .A3(new_n268), .A4(new_n500), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n268), .A2(G116), .ZN(new_n654));
  AOI21_X1  g0454(.A(G20), .B1(G33), .B2(G283), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n251), .A2(G97), .ZN(new_n656));
  INV_X1    g0456(.A(G116), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n655), .A2(new_n656), .B1(G20), .B2(new_n657), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n658), .A2(new_n263), .A3(KEYINPUT20), .ZN(new_n659));
  AOI21_X1  g0459(.A(KEYINPUT20), .B1(new_n658), .B2(new_n263), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n653), .B(new_n654), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n652), .A2(new_n661), .A3(G169), .ZN(new_n662));
  NOR2_X1   g0462(.A1(KEYINPUT88), .A2(KEYINPUT21), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n652), .A2(G200), .ZN(new_n665));
  INV_X1    g0465(.A(new_n661), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n650), .A2(G190), .A3(new_n651), .A4(new_n614), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n663), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n652), .A2(new_n661), .A3(G169), .A4(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n651), .A2(new_n614), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n671), .A2(new_n661), .A3(G179), .A4(new_n650), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n664), .A2(new_n668), .A3(new_n670), .A4(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT89), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n652), .A2(new_n300), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n662), .A2(new_n663), .B1(new_n675), .B2(new_n661), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT89), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n676), .A2(new_n677), .A3(new_n670), .A4(new_n668), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n643), .A2(new_n679), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n460), .A2(new_n583), .A3(new_n680), .ZN(G372));
  AND2_X1   g0481(.A1(new_n335), .A2(new_n324), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n385), .B1(new_n682), .B2(new_n377), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n457), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n446), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n303), .B1(new_n685), .B2(new_n398), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n540), .A2(new_n555), .A3(new_n567), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n573), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT26), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n568), .A2(new_n576), .A3(new_n573), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n576), .B1(new_n568), .B2(new_n573), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n691), .A2(new_n692), .A3(new_n582), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n690), .B1(new_n693), .B2(KEYINPUT26), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n527), .A2(new_n582), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n600), .A2(new_n608), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n641), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(new_n670), .A3(new_n676), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n626), .A2(new_n689), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n573), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n459), .B1(new_n694), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n686), .A2(new_n701), .ZN(G369));
  AND2_X1   g0502(.A1(new_n204), .A2(G13), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n528), .A2(new_n703), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n704), .A2(KEYINPUT27), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(KEYINPUT27), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(G213), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G343), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n666), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n710), .B1(new_n674), .B2(new_n678), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n664), .A2(new_n670), .A3(new_n672), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n711), .B1(new_n713), .B2(new_n710), .ZN(new_n714));
  INV_X1    g0514(.A(G330), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n709), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n638), .A2(new_n639), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n643), .A2(new_n718), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n642), .A2(new_n709), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT93), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT93), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n716), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n697), .A2(new_n717), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n712), .A2(new_n717), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT94), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n727), .B1(new_n721), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n726), .A2(new_n730), .ZN(G399));
  NAND2_X1  g0531(.A1(new_n207), .A2(new_n490), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n541), .A2(new_n657), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n732), .A2(G1), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(new_n218), .B2(new_n732), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT28), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  AND4_X1   g0537(.A1(new_n563), .A2(new_n562), .A3(new_n616), .A4(new_n617), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n675), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n737), .B1(new_n739), .B2(new_n523), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n480), .A2(new_n495), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n741), .A2(KEYINPUT30), .A3(new_n675), .A4(new_n738), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n569), .A2(new_n652), .A3(new_n300), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(new_n523), .A3(new_n622), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n740), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n717), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT31), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n745), .A2(KEYINPUT31), .A3(new_n717), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n679), .A2(new_n642), .A3(new_n626), .A4(new_n709), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n748), .B(new_n749), .C1(new_n750), .C2(new_n583), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n715), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n573), .A2(new_n688), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(new_n621), .B2(new_n625), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n642), .A2(new_n712), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n756), .A2(new_n527), .A3(new_n757), .A4(new_n582), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT26), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n575), .A2(new_n687), .A3(new_n759), .A4(new_n577), .ZN(new_n760));
  INV_X1    g0560(.A(new_n573), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n689), .A2(new_n581), .A3(new_n579), .A4(new_n578), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n761), .B1(new_n762), .B2(KEYINPUT26), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n758), .A2(new_n760), .A3(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(KEYINPUT29), .A3(new_n709), .ZN(new_n765));
  INV_X1    g0565(.A(new_n699), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n687), .B1(new_n522), .B2(new_n526), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n761), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n690), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n575), .A2(new_n687), .A3(KEYINPUT26), .A4(new_n577), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n717), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n765), .B1(new_n772), .B2(KEYINPUT29), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n754), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n736), .B1(new_n775), .B2(G1), .ZN(G364));
  AOI21_X1  g0576(.A(new_n203), .B1(new_n703), .B2(G45), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n732), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n716), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n714), .A2(new_n715), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G13), .A2(G33), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n204), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT95), .Z(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT100), .Z(new_n785));
  NAND2_X1  g0585(.A1(new_n714), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n207), .A2(new_n283), .ZN(new_n787));
  INV_X1    g0587(.A(G355), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n787), .A2(new_n788), .B1(G116), .B2(new_n207), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n243), .A2(G45), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n207), .A2(new_n414), .ZN(new_n791));
  INV_X1    g0591(.A(G45), .ZN(new_n792));
  INV_X1    g0592(.A(new_n218), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n789), .B1(new_n790), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n215), .B1(G20), .B2(new_n375), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n796), .A2(KEYINPUT96), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(KEYINPUT96), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n784), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n779), .B1(new_n795), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n204), .A2(G190), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n300), .A2(G200), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(G190), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n283), .B1(new_n805), .B2(new_n285), .C1(new_n808), .C2(new_n257), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n204), .A2(new_n325), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n389), .A2(G179), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n811), .A2(new_n803), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(G87), .A2(new_n813), .B1(new_n815), .B2(G107), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n810), .A2(new_n804), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n253), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n806), .A2(new_n325), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n809), .B(new_n818), .C1(G50), .C2(new_n819), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n300), .A2(new_n389), .A3(KEYINPUT97), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(KEYINPUT97), .B1(new_n300), .B2(new_n389), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n803), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(G159), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT32), .Z(new_n828));
  INV_X1    g0628(.A(new_n824), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n204), .B1(new_n829), .B2(G190), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(G97), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n820), .A2(new_n828), .A3(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(KEYINPUT33), .B(G317), .Z(new_n834));
  INV_X1    g0634(.A(new_n819), .ZN(new_n835));
  INV_X1    g0635(.A(G326), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n808), .A2(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n817), .ZN(new_n838));
  INV_X1    g0638(.A(new_n805), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G322), .A2(new_n838), .B1(new_n839), .B2(G311), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n464), .B2(new_n814), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n837), .B(new_n841), .C1(G329), .C2(new_n826), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n611), .B2(new_n830), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n812), .B(KEYINPUT98), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n283), .B1(new_n844), .B2(G303), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT99), .Z(new_n846));
  OAI21_X1  g0646(.A(new_n833), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n802), .B1(new_n847), .B2(new_n799), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n780), .A2(new_n781), .B1(new_n786), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G396));
  INV_X1    g0650(.A(new_n373), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n348), .A2(new_n717), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(new_n377), .B2(KEYINPUT101), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n377), .A2(KEYINPUT101), .A3(new_n852), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n851), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n772), .A2(new_n856), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n709), .B(new_n856), .C1(new_n694), .C2(new_n700), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n779), .B1(new_n859), .B2(new_n754), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n754), .B2(new_n859), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n799), .A2(new_n782), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n778), .B1(new_n862), .B2(new_n285), .ZN(new_n863));
  AOI22_X1  g0663(.A1(G143), .A2(new_n838), .B1(new_n839), .B2(G159), .ZN(new_n864));
  INV_X1    g0664(.A(G137), .ZN(new_n865));
  INV_X1    g0665(.A(G150), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n864), .B1(new_n835), .B2(new_n865), .C1(new_n866), .C2(new_n808), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT34), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n826), .A2(G132), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n414), .B1(new_n815), .B2(G68), .ZN(new_n870));
  INV_X1    g0670(.A(new_n844), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n869), .B(new_n870), .C1(new_n871), .C2(new_n256), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(G58), .B2(new_n831), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n283), .B1(new_n838), .B2(G294), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n844), .A2(G107), .B1(new_n826), .B2(G311), .ZN(new_n875));
  AOI22_X1  g0675(.A1(G87), .A2(new_n815), .B1(new_n839), .B2(G116), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n807), .A2(G283), .B1(new_n819), .B2(G303), .ZN(new_n877));
  AND4_X1   g0677(.A1(new_n874), .A2(new_n875), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n868), .A2(new_n873), .B1(new_n832), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n782), .ZN(new_n880));
  OAI221_X1 g0680(.A(new_n863), .B1(new_n800), .B2(new_n879), .C1(new_n856), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n861), .A2(new_n881), .ZN(G384));
  INV_X1    g0682(.A(KEYINPUT40), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n385), .A2(KEYINPUT102), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT102), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n885), .B(new_n379), .C1(new_n383), .C2(new_n384), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n378), .A2(new_n709), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n335), .B2(new_n324), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n884), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n887), .B1(new_n383), .B2(new_n384), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n751), .A2(new_n856), .A3(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n428), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT103), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n407), .B2(new_n412), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n417), .A2(new_n421), .A3(KEYINPUT103), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(new_n399), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n407), .A2(new_n412), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n270), .B1(new_n898), .B2(KEYINPUT16), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n893), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n441), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n450), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n900), .A2(new_n707), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT37), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n429), .A2(new_n708), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT37), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n442), .A2(new_n905), .A3(new_n906), .A4(new_n450), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n443), .A2(new_n445), .A3(new_n452), .A4(new_n456), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n903), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n908), .A2(new_n910), .A3(KEYINPUT38), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n908), .B2(new_n910), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n883), .B1(new_n892), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT105), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI211_X1 g0716(.A(KEYINPUT105), .B(new_n883), .C1(new_n892), .C2(new_n913), .ZN(new_n917));
  INV_X1    g0717(.A(new_n892), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n442), .A2(new_n905), .A3(new_n450), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT37), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n920), .A2(KEYINPUT104), .A3(new_n907), .ZN(new_n921));
  INV_X1    g0721(.A(new_n905), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n909), .A2(new_n922), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n921), .B(new_n923), .C1(KEYINPUT104), .C2(new_n920), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT38), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n911), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n883), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n916), .A2(new_n917), .B1(new_n918), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n459), .A2(new_n751), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT106), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n929), .A2(new_n931), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n932), .A2(new_n933), .A3(new_n715), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT39), .B1(new_n926), .B2(new_n927), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT39), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n911), .A2(new_n912), .A3(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n717), .B1(new_n884), .B2(new_n886), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n891), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n377), .A2(new_n717), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n941), .B1(new_n858), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n911), .B2(new_n912), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n446), .A2(new_n708), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n940), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n459), .B(new_n765), .C1(new_n772), .C2(KEYINPUT29), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n947), .A2(new_n686), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n946), .B(new_n948), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n934), .A2(new_n949), .B1(new_n528), .B2(new_n703), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n949), .B2(new_n934), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n505), .A2(new_n511), .A3(new_n514), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT35), .ZN(new_n953));
  OAI211_X1 g0753(.A(G116), .B(new_n216), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n953), .B2(new_n952), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT36), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n793), .B(G77), .C1(new_n253), .C2(new_n257), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n256), .A2(G68), .ZN(new_n958));
  AOI211_X1 g0758(.A(G13), .B(new_n528), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  OR3_X1    g0759(.A1(new_n951), .A2(new_n956), .A3(new_n959), .ZN(G367));
  AND2_X1   g0760(.A1(new_n721), .A2(new_n729), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n767), .B1(new_n519), .B2(new_n709), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n687), .A2(new_n717), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT42), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT43), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n582), .B1(new_n962), .B2(new_n642), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT107), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n717), .B1(new_n969), .B2(new_n970), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n709), .A2(new_n555), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n755), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n761), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n967), .A2(new_n968), .A3(new_n973), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n968), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n981));
  INV_X1    g0781(.A(new_n973), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n980), .B(new_n981), .C1(new_n966), .C2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n964), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n984), .B1(new_n726), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n726), .A2(new_n985), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n979), .A2(new_n987), .A3(new_n983), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n732), .B(KEYINPUT41), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n721), .A2(new_n729), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n961), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n716), .A2(KEYINPUT109), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n994), .B(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n775), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n730), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(KEYINPUT45), .B1(new_n730), .B2(new_n964), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT44), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n730), .B2(new_n964), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n999), .A2(new_n1000), .B1(new_n1002), .B2(KEYINPUT108), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n726), .A2(KEYINPUT110), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n730), .A2(new_n964), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(KEYINPUT44), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1007), .A2(KEYINPUT108), .A3(new_n1002), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n726), .A2(KEYINPUT110), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1004), .A2(new_n1005), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  AND3_X1   g0810(.A1(new_n1007), .A2(KEYINPUT108), .A3(new_n1002), .ZN(new_n1011));
  OAI211_X1 g0811(.A(KEYINPUT110), .B(new_n726), .C1(new_n1011), .C2(new_n1003), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n997), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n992), .B1(new_n1013), .B2(new_n774), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n777), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n990), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n831), .A2(G68), .ZN(new_n1017));
  INV_X1    g0817(.A(G159), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n283), .B1(new_n817), .B2(new_n866), .C1(new_n1018), .C2(new_n808), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G143), .B2(new_n819), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(KEYINPUT112), .B(G137), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n826), .A2(new_n1022), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n812), .A2(new_n253), .B1(new_n805), .B2(new_n256), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n814), .A2(new_n285), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1017), .A2(new_n1020), .A3(new_n1023), .A4(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(KEYINPUT46), .B1(new_n813), .B2(G116), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G311), .B2(new_n819), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n611), .B2(new_n808), .C1(new_n830), .C2(new_n586), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n844), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n826), .A2(G317), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n283), .B1(new_n839), .B2(G283), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n644), .A2(new_n645), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n1034), .A2(new_n838), .B1(new_n815), .B2(G97), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .A4(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1027), .B1(new_n1030), .B2(new_n1036), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT113), .Z(new_n1038));
  AOI21_X1  g0838(.A(new_n800), .B1(new_n1038), .B2(KEYINPUT47), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(KEYINPUT47), .B2(new_n1038), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n978), .A2(new_n785), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n238), .A2(new_n791), .B1(new_n207), .B2(new_n337), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n779), .B1(new_n801), .B2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT111), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1040), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1016), .A2(new_n1045), .ZN(G387));
  INV_X1    g0846(.A(new_n777), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n719), .A2(new_n720), .A3(new_n785), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n787), .A2(new_n733), .B1(G107), .B2(new_n207), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n235), .A2(new_n792), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n733), .B(new_n792), .C1(new_n257), .C2(new_n285), .ZN(new_n1051));
  XOR2_X1   g0851(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n1052));
  NOR3_X1   g0852(.A1(new_n1052), .A2(G50), .A3(new_n248), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1052), .B1(G50), .B2(new_n248), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n791), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1049), .B1(new_n1050), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n779), .B1(new_n1057), .B2(new_n801), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n256), .A2(new_n817), .B1(new_n812), .B2(new_n285), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n283), .B1(new_n814), .B2(new_n498), .C1(new_n835), .C2(new_n1018), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(G68), .C2(new_n839), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n831), .A2(new_n338), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n425), .A2(new_n807), .B1(new_n826), .B2(G150), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n283), .B1(new_n815), .B2(G116), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n826), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G317), .A2(new_n838), .B1(new_n839), .B2(new_n1034), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n819), .A2(G322), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n807), .A2(G311), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT48), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n831), .A2(G283), .B1(G294), .B2(new_n813), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT49), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1065), .B1(new_n836), .B2(new_n1066), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1064), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1058), .B1(new_n1079), .B2(new_n799), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n996), .A2(new_n1047), .B1(new_n1048), .B2(new_n1080), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n732), .B(KEYINPUT115), .Z(new_n1082));
  NAND2_X1  g0882(.A1(new_n997), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n996), .A2(new_n775), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1081), .B1(new_n1083), .B2(new_n1084), .ZN(G393));
  INV_X1    g0885(.A(new_n1082), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1013), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1010), .A2(new_n1012), .A3(new_n997), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n1047), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n964), .A2(new_n784), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT116), .Z(new_n1093));
  INV_X1    g0893(.A(new_n246), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n1094), .A2(new_n791), .B1(new_n498), .B2(new_n207), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n779), .B1(new_n801), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n414), .B1(new_n814), .B2(new_n586), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n812), .A2(new_n464), .B1(new_n805), .B2(new_n611), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1097), .B(new_n1098), .C1(new_n1034), .C2(new_n807), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n826), .A2(G322), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1099), .B(new_n1100), .C1(new_n657), .C2(new_n830), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n838), .A2(G311), .B1(G317), .B2(new_n819), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT52), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n831), .A2(G77), .ZN(new_n1104));
  INV_X1    g0904(.A(G87), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n283), .B1(new_n814), .B2(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n812), .A2(new_n257), .B1(new_n805), .B2(new_n248), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(G50), .C2(new_n807), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n826), .A2(G143), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1104), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n835), .A2(new_n866), .B1(new_n817), .B2(new_n1018), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(KEYINPUT117), .B(KEYINPUT51), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1111), .B(new_n1112), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n1101), .A2(new_n1103), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1096), .B1(new_n1114), .B2(new_n799), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1093), .A2(new_n1115), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1091), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1089), .A2(new_n1117), .ZN(G390));
  NAND2_X1  g0918(.A1(new_n753), .A2(new_n459), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1119), .A2(new_n947), .A3(new_n686), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n750), .A2(new_n583), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n748), .A2(new_n749), .ZN(new_n1122));
  OAI211_X1 g0922(.A(G330), .B(new_n856), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n941), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n764), .A2(new_n709), .A3(new_n856), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1125), .A2(new_n942), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n751), .A2(new_n891), .A3(G330), .A4(new_n856), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1124), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT118), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n858), .A2(new_n942), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1128), .A2(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1124), .A2(new_n1126), .A3(KEYINPUT118), .A4(new_n1127), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1120), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n943), .A2(new_n939), .B1(new_n935), .B2(new_n937), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n939), .B1(new_n926), .B2(new_n927), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n1126), .B2(new_n941), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1127), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1136), .A2(new_n1127), .A3(new_n1138), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1086), .B1(new_n1135), .B2(new_n1143), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1136), .A2(new_n1138), .A3(new_n1127), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1127), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n1134), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1144), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1147), .A2(new_n1047), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n862), .ZN(new_n1151));
  XOR2_X1   g0951(.A(KEYINPUT119), .B(KEYINPUT53), .Z(new_n1152));
  OR3_X1    g0952(.A1(new_n1152), .A2(new_n812), .A3(new_n866), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1022), .A2(new_n807), .B1(G128), .B2(new_n819), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1152), .B1(new_n812), .B2(new_n866), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n826), .A2(G125), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n414), .B1(new_n815), .B2(G50), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT54), .B(G143), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G132), .A2(new_n838), .B1(new_n839), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1157), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1156), .B(new_n1162), .C1(G159), .C2(new_n831), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1104), .B1(new_n657), .B2(new_n817), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT120), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n871), .A2(new_n1105), .B1(new_n1066), .B2(new_n611), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n283), .B1(new_n815), .B2(G68), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n498), .B2(new_n805), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n808), .A2(new_n586), .B1(new_n835), .B2(new_n464), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1166), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1163), .B1(new_n1165), .B2(new_n1170), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n779), .B1(new_n425), .B2(new_n1151), .C1(new_n1171), .C2(new_n800), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1172), .B(KEYINPUT121), .Z(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n938), .B2(new_n880), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1150), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1149), .A2(new_n1175), .ZN(G378));
  INV_X1    g0976(.A(new_n303), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n398), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n277), .A2(new_n707), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1179), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n398), .A2(new_n1177), .A3(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1180), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1183), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1181), .B1(new_n398), .B2(new_n1177), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1179), .B(new_n303), .C1(new_n395), .C2(new_n397), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1185), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1184), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT122), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1184), .A2(new_n1188), .A3(KEYINPUT122), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1193), .A2(new_n880), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n283), .A2(G41), .ZN(new_n1195));
  AOI211_X1 g0995(.A(G50), .B(new_n1195), .C1(new_n251), .C2(new_n490), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n338), .A2(new_n839), .B1(new_n815), .B2(G58), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n586), .B2(new_n817), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G283), .B2(new_n826), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1195), .B1(new_n285), .B2(new_n812), .C1(new_n835), .C2(new_n657), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G97), .B2(new_n807), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1017), .A3(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT58), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1196), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n812), .A2(new_n1159), .B1(new_n805), .B2(new_n865), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G128), .B2(new_n838), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n807), .A2(G132), .B1(new_n819), .B2(G125), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n866), .C2(new_n830), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n251), .B(new_n490), .C1(new_n814), .C2(new_n1018), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n826), .B2(G124), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1204), .B1(new_n1203), .B2(new_n1202), .C1(new_n1209), .C2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n799), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1215), .B(new_n779), .C1(G50), .C2(new_n1151), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1194), .A2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n715), .B1(new_n928), .B2(new_n918), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n917), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n377), .A2(KEYINPUT101), .A3(new_n852), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n373), .B1(new_n1220), .B2(new_n853), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n889), .B2(new_n890), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1222), .B(new_n751), .C1(new_n911), .C2(new_n912), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT105), .B1(new_n1223), .B2(new_n883), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1218), .B(new_n1193), .C1(new_n1219), .C2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n920), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT104), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1226), .A2(new_n1227), .B1(new_n909), .B2(new_n922), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT38), .B1(new_n1228), .B2(new_n921), .ZN(new_n1229));
  OAI21_X1  g1029(.A(KEYINPUT40), .B1(new_n1229), .B2(new_n911), .ZN(new_n1230));
  OAI21_X1  g1030(.A(G330), .B1(new_n1230), .B2(new_n892), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n916), .B2(new_n917), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n946), .B(new_n1225), .C1(new_n1232), .C2(new_n1189), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1218), .B1(new_n1219), .B2(new_n1224), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1189), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n946), .B1(new_n1237), .B2(new_n1225), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1234), .A2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1217), .B1(new_n1239), .B2(new_n1047), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1120), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1148), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT57), .B1(new_n1239), .B2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1225), .B1(new_n1232), .B2(new_n1189), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n946), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1246), .A2(KEYINPUT57), .A3(new_n1233), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1120), .B1(new_n1147), .B2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1082), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1240), .B1(new_n1243), .B2(new_n1250), .ZN(G375));
  NAND2_X1  g1051(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1252), .A2(new_n1120), .A3(new_n1133), .A4(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1135), .A2(new_n992), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n941), .A2(new_n782), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1256), .B(KEYINPUT123), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n779), .B1(new_n1151), .B2(G68), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n817), .A2(new_n464), .B1(new_n805), .B2(new_n586), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1259), .A2(new_n283), .A3(new_n1025), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n807), .A2(G116), .B1(new_n819), .B2(G294), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n844), .A2(G97), .B1(new_n826), .B2(G303), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1062), .A2(new_n1260), .A3(new_n1261), .A4(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n830), .A2(new_n256), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n844), .A2(G159), .B1(new_n826), .B2(G128), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n414), .B1(new_n815), .B2(G58), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n838), .A2(new_n1022), .B1(new_n839), .B2(G150), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n1160), .A2(new_n807), .B1(G132), .B2(new_n819), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .A4(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1263), .B1(new_n1264), .B2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1258), .B1(new_n799), .B2(new_n1270), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n1248), .A2(new_n1047), .B1(new_n1257), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1255), .A2(new_n1272), .ZN(G381));
  NAND4_X1  g1073(.A1(new_n1016), .A2(new_n1045), .A3(new_n1089), .A4(new_n1117), .ZN(new_n1274));
  NOR4_X1   g1074(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1150), .A2(new_n1174), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(new_n1144), .B2(new_n1148), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  OR2_X1    g1078(.A1(new_n1274), .A2(new_n1278), .ZN(new_n1279));
  OR2_X1    g1079(.A1(new_n1279), .A2(G375), .ZN(G407));
  INV_X1    g1080(.A(G213), .ZN(new_n1281));
  OR3_X1    g1081(.A1(new_n1281), .A2(KEYINPUT124), .A3(G343), .ZN(new_n1282));
  OAI21_X1  g1082(.A(KEYINPUT124), .B1(new_n1281), .B2(G343), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1284), .B(KEYINPUT125), .ZN(new_n1285));
  OR3_X1    g1085(.A1(G375), .A2(G378), .A3(new_n1285), .ZN(new_n1286));
  OAI211_X1 g1086(.A(G213), .B(new_n1286), .C1(new_n1279), .C2(G375), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1287), .B(KEYINPUT126), .ZN(G409));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1285), .ZN(new_n1290));
  OAI211_X1 g1090(.A(G378), .B(new_n1240), .C1(new_n1243), .C2(new_n1250), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1246), .A2(new_n1233), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1292), .A2(new_n1249), .A3(new_n991), .ZN(new_n1293));
  OAI22_X1  g1093(.A1(new_n1292), .A2(new_n777), .B1(new_n1194), .B2(new_n1216), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1277), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1290), .B1(new_n1291), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1254), .A2(KEYINPUT60), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT60), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1132), .A2(new_n1298), .A3(new_n1120), .A4(new_n1133), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1086), .B1(new_n1248), .B2(new_n1241), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1302), .A2(G384), .A3(new_n1272), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(G384), .B1(new_n1302), .B2(new_n1272), .ZN(new_n1305));
  OAI211_X1 g1105(.A(G2897), .B(new_n1290), .C1(new_n1304), .C2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1302), .A2(new_n1272), .ZN(new_n1307));
  INV_X1    g1107(.A(G384), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(G2897), .ZN(new_n1310));
  OAI211_X1 g1110(.A(new_n1309), .B(new_n1303), .C1(new_n1310), .C2(new_n1284), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1306), .A2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1289), .B1(new_n1296), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(KEYINPUT127), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1291), .A2(new_n1295), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1309), .A2(new_n1303), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1315), .A2(KEYINPUT62), .A3(new_n1285), .A4(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1284), .ZN(new_n1319));
  AOI211_X1 g1119(.A(new_n1319), .B(new_n1316), .C1(new_n1291), .C2(new_n1295), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1318), .B1(new_n1320), .B2(KEYINPUT62), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT127), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1322), .B(new_n1289), .C1(new_n1296), .C2(new_n1312), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1314), .A2(new_n1321), .A3(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n989), .B1(new_n1014), .B2(new_n777), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1045), .ZN(new_n1326));
  OAI21_X1  g1126(.A(G390), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(G393), .B(G396), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1274), .A2(new_n1327), .A3(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1328), .B1(new_n1274), .B2(new_n1327), .ZN(new_n1330));
  OR2_X1    g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1324), .A2(new_n1331), .ZN(new_n1332));
  NOR3_X1   g1132(.A1(new_n1329), .A2(new_n1330), .A3(KEYINPUT61), .ZN(new_n1333));
  OR2_X1    g1133(.A1(new_n1320), .A2(KEYINPUT63), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1296), .A2(KEYINPUT63), .A3(new_n1317), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1315), .A2(new_n1284), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1336), .A2(new_n1311), .A3(new_n1306), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1333), .A2(new_n1334), .A3(new_n1335), .A4(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1332), .A2(new_n1338), .ZN(G405));
  NAND2_X1  g1139(.A1(G375), .A2(new_n1277), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(new_n1291), .ZN(new_n1341));
  XNOR2_X1  g1141(.A(new_n1341), .B(new_n1317), .ZN(new_n1342));
  XNOR2_X1  g1142(.A(new_n1331), .B(new_n1342), .ZN(G402));
endmodule


