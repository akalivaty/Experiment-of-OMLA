

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589;

  XNOR2_X1 U323 ( .A(n324), .B(n323), .ZN(n327) );
  XNOR2_X1 U324 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U325 ( .A(n392), .B(KEYINPUT120), .Z(n291) );
  XOR2_X1 U326 ( .A(G85GAT), .B(G92GAT), .Z(n317) );
  AND2_X1 U327 ( .A1(n569), .A2(n430), .ZN(n431) );
  XNOR2_X1 U328 ( .A(n393), .B(n291), .ZN(n569) );
  INV_X1 U329 ( .A(KEYINPUT122), .ZN(n447) );
  XNOR2_X1 U330 ( .A(n307), .B(n306), .ZN(n578) );
  XNOR2_X1 U331 ( .A(n448), .B(n447), .ZN(n565) );
  XNOR2_X1 U332 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U333 ( .A(n455), .B(n454), .ZN(G1351GAT) );
  INV_X1 U334 ( .A(KEYINPUT55), .ZN(n432) );
  XNOR2_X1 U335 ( .A(KEYINPUT48), .B(KEYINPUT113), .ZN(n372) );
  XNOR2_X1 U336 ( .A(G106GAT), .B(G78GAT), .ZN(n292) );
  XNOR2_X1 U337 ( .A(n292), .B(G148GAT), .ZN(n422) );
  XNOR2_X1 U338 ( .A(G57GAT), .B(KEYINPUT69), .ZN(n293) );
  XNOR2_X1 U339 ( .A(n293), .B(KEYINPUT13), .ZN(n338) );
  XOR2_X1 U340 ( .A(n422), .B(n338), .Z(n307) );
  XOR2_X1 U341 ( .A(G176GAT), .B(G64GAT), .Z(n387) );
  XNOR2_X1 U342 ( .A(G204GAT), .B(n387), .ZN(n297) );
  XOR2_X1 U343 ( .A(KEYINPUT70), .B(KEYINPUT72), .Z(n295) );
  XNOR2_X1 U344 ( .A(KEYINPUT73), .B(KEYINPUT31), .ZN(n294) );
  XNOR2_X1 U345 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U346 ( .A(n297), .B(n296), .ZN(n299) );
  XOR2_X1 U347 ( .A(KEYINPUT71), .B(n317), .Z(n298) );
  XNOR2_X1 U348 ( .A(n299), .B(n298), .ZN(n301) );
  AND2_X1 U349 ( .A1(G230GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U350 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U351 ( .A(KEYINPUT33), .B(n302), .Z(n305) );
  XNOR2_X1 U352 ( .A(G99GAT), .B(G71GAT), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n303), .B(G120GAT), .ZN(n436) );
  XNOR2_X1 U354 ( .A(n436), .B(KEYINPUT32), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U356 ( .A(KEYINPUT9), .B(KEYINPUT77), .Z(n309) );
  XNOR2_X1 U357 ( .A(G99GAT), .B(KEYINPUT11), .ZN(n308) );
  XNOR2_X1 U358 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U359 ( .A(KEYINPUT10), .B(KEYINPUT64), .Z(n311) );
  XNOR2_X1 U360 ( .A(G190GAT), .B(KEYINPUT78), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U362 ( .A(n313), .B(n312), .ZN(n329) );
  XOR2_X1 U363 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n315) );
  XNOR2_X1 U364 ( .A(G36GAT), .B(G29GAT), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U366 ( .A(KEYINPUT7), .B(n316), .Z(n352) );
  XOR2_X1 U367 ( .A(KEYINPUT76), .B(n317), .Z(n319) );
  XOR2_X1 U368 ( .A(G43GAT), .B(G134GAT), .Z(n442) );
  XNOR2_X1 U369 ( .A(n442), .B(G218GAT), .ZN(n318) );
  XOR2_X1 U370 ( .A(n319), .B(n318), .Z(n320) );
  XNOR2_X1 U371 ( .A(n352), .B(n320), .ZN(n324) );
  NAND2_X1 U372 ( .A1(G232GAT), .A2(G233GAT), .ZN(n322) );
  INV_X1 U373 ( .A(KEYINPUT65), .ZN(n321) );
  XNOR2_X1 U374 ( .A(G50GAT), .B(KEYINPUT75), .ZN(n325) );
  XNOR2_X1 U375 ( .A(n325), .B(G162GAT), .ZN(n424) );
  XNOR2_X1 U376 ( .A(n424), .B(G106GAT), .ZN(n326) );
  XNOR2_X1 U377 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U378 ( .A(n329), .B(n328), .ZN(n545) );
  INV_X1 U379 ( .A(n545), .ZN(n561) );
  XNOR2_X1 U380 ( .A(KEYINPUT36), .B(n561), .ZN(n586) );
  XOR2_X1 U381 ( .A(KEYINPUT80), .B(G64GAT), .Z(n331) );
  XNOR2_X1 U382 ( .A(G155GAT), .B(G78GAT), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U384 ( .A(KEYINPUT14), .B(KEYINPUT81), .Z(n333) );
  XNOR2_X1 U385 ( .A(KEYINPUT79), .B(KEYINPUT12), .ZN(n332) );
  XNOR2_X1 U386 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U387 ( .A(n335), .B(n334), .ZN(n346) );
  XOR2_X1 U388 ( .A(G15GAT), .B(G127GAT), .Z(n440) );
  XOR2_X1 U389 ( .A(G71GAT), .B(n440), .Z(n337) );
  XOR2_X1 U390 ( .A(G1GAT), .B(G8GAT), .Z(n355) );
  XNOR2_X1 U391 ( .A(n355), .B(G183GAT), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n337), .B(n336), .ZN(n342) );
  XOR2_X1 U393 ( .A(n338), .B(KEYINPUT15), .Z(n340) );
  NAND2_X1 U394 ( .A1(G231GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U396 ( .A(n342), .B(n341), .Z(n344) );
  XNOR2_X1 U397 ( .A(G22GAT), .B(G211GAT), .ZN(n343) );
  XNOR2_X1 U398 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U399 ( .A(n346), .B(n345), .ZN(n557) );
  NOR2_X1 U400 ( .A1(n586), .A2(n557), .ZN(n347) );
  XOR2_X1 U401 ( .A(KEYINPUT45), .B(n347), .Z(n348) );
  NOR2_X1 U402 ( .A1(n578), .A2(n348), .ZN(n364) );
  XOR2_X1 U403 ( .A(G197GAT), .B(G15GAT), .Z(n350) );
  XNOR2_X1 U404 ( .A(G169GAT), .B(G113GAT), .ZN(n349) );
  XNOR2_X1 U405 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n363) );
  XOR2_X1 U407 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n354) );
  XNOR2_X1 U408 ( .A(KEYINPUT67), .B(KEYINPUT30), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n359) );
  XOR2_X1 U410 ( .A(G50GAT), .B(G43GAT), .Z(n357) );
  XOR2_X1 U411 ( .A(G141GAT), .B(G22GAT), .Z(n419) );
  XNOR2_X1 U412 ( .A(n419), .B(n355), .ZN(n356) );
  XNOR2_X1 U413 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U414 ( .A(n359), .B(n358), .Z(n361) );
  NAND2_X1 U415 ( .A1(G229GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n363), .B(n362), .ZN(n573) );
  INV_X1 U418 ( .A(n573), .ZN(n551) );
  NAND2_X1 U419 ( .A1(n364), .A2(n551), .ZN(n370) );
  XNOR2_X1 U420 ( .A(n578), .B(KEYINPUT41), .ZN(n553) );
  OR2_X1 U421 ( .A1(n551), .A2(n553), .ZN(n365) );
  XNOR2_X1 U422 ( .A(KEYINPUT46), .B(n365), .ZN(n367) );
  INV_X1 U423 ( .A(n557), .ZN(n581) );
  NOR2_X1 U424 ( .A1(n545), .A2(n581), .ZN(n366) );
  AND2_X1 U425 ( .A1(n367), .A2(n366), .ZN(n368) );
  XNOR2_X1 U426 ( .A(n368), .B(KEYINPUT47), .ZN(n369) );
  NAND2_X1 U427 ( .A1(n370), .A2(n369), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n372), .B(n371), .ZN(n532) );
  XNOR2_X1 U429 ( .A(G169GAT), .B(G183GAT), .ZN(n379) );
  XOR2_X1 U430 ( .A(KEYINPUT19), .B(KEYINPUT86), .Z(n374) );
  XNOR2_X1 U431 ( .A(KEYINPUT17), .B(KEYINPUT87), .ZN(n373) );
  XNOR2_X1 U432 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U433 ( .A(n375), .B(KEYINPUT88), .Z(n377) );
  XNOR2_X1 U434 ( .A(G190GAT), .B(KEYINPUT18), .ZN(n376) );
  XNOR2_X1 U435 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n443) );
  XNOR2_X1 U437 ( .A(G211GAT), .B(G218GAT), .ZN(n380) );
  XNOR2_X1 U438 ( .A(n380), .B(KEYINPUT91), .ZN(n381) );
  XOR2_X1 U439 ( .A(n381), .B(KEYINPUT21), .Z(n383) );
  XNOR2_X1 U440 ( .A(G197GAT), .B(G204GAT), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n383), .B(n382), .ZN(n429) );
  XNOR2_X1 U442 ( .A(n443), .B(n429), .ZN(n391) );
  XOR2_X1 U443 ( .A(KEYINPUT95), .B(G92GAT), .Z(n385) );
  XNOR2_X1 U444 ( .A(G36GAT), .B(G8GAT), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U446 ( .A(n387), .B(n386), .Z(n389) );
  NAND2_X1 U447 ( .A1(G226GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U449 ( .A(n391), .B(n390), .ZN(n493) );
  NOR2_X1 U450 ( .A1(n532), .A2(n493), .ZN(n393) );
  XNOR2_X1 U451 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n392) );
  XOR2_X1 U452 ( .A(G148GAT), .B(G120GAT), .Z(n395) );
  XNOR2_X1 U453 ( .A(G141GAT), .B(G127GAT), .ZN(n394) );
  XNOR2_X1 U454 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U455 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n397) );
  XNOR2_X1 U456 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n396) );
  XNOR2_X1 U457 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U458 ( .A(n399), .B(n398), .Z(n406) );
  XOR2_X1 U459 ( .A(G85GAT), .B(G162GAT), .Z(n403) );
  XOR2_X1 U460 ( .A(KEYINPUT84), .B(KEYINPUT0), .Z(n401) );
  XNOR2_X1 U461 ( .A(G113GAT), .B(KEYINPUT83), .ZN(n400) );
  XNOR2_X1 U462 ( .A(n401), .B(n400), .ZN(n437) );
  XNOR2_X1 U463 ( .A(G29GAT), .B(n437), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U465 ( .A(G134GAT), .B(n404), .ZN(n405) );
  XNOR2_X1 U466 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U467 ( .A(G57GAT), .B(KEYINPUT94), .Z(n408) );
  NAND2_X1 U468 ( .A1(G225GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U469 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U470 ( .A(n410), .B(n409), .Z(n415) );
  XOR2_X1 U471 ( .A(KEYINPUT3), .B(KEYINPUT93), .Z(n412) );
  XNOR2_X1 U472 ( .A(KEYINPUT92), .B(G155GAT), .ZN(n411) );
  XNOR2_X1 U473 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U474 ( .A(KEYINPUT2), .B(n413), .Z(n425) );
  XNOR2_X1 U475 ( .A(G1GAT), .B(n425), .ZN(n414) );
  XNOR2_X1 U476 ( .A(n415), .B(n414), .ZN(n570) );
  INV_X1 U477 ( .A(n570), .ZN(n530) );
  XOR2_X1 U478 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n417) );
  XNOR2_X1 U479 ( .A(KEYINPUT90), .B(KEYINPUT23), .ZN(n416) );
  XNOR2_X1 U480 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U481 ( .A(n419), .B(n418), .Z(n421) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U483 ( .A(n421), .B(n420), .ZN(n423) );
  XOR2_X1 U484 ( .A(n423), .B(n422), .Z(n427) );
  XNOR2_X1 U485 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U486 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n464) );
  NOR2_X1 U488 ( .A1(n530), .A2(n464), .ZN(n430) );
  XNOR2_X1 U489 ( .A(n432), .B(n431), .ZN(n446) );
  XOR2_X1 U490 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n434) );
  NAND2_X1 U491 ( .A1(G227GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U493 ( .A(n435), .B(G176GAT), .Z(n439) );
  XNOR2_X1 U494 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n441) );
  XOR2_X1 U496 ( .A(n441), .B(n440), .Z(n445) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n533) );
  NAND2_X1 U499 ( .A1(n446), .A2(n533), .ZN(n448) );
  INV_X1 U500 ( .A(n553), .ZN(n538) );
  NAND2_X1 U501 ( .A1(n565), .A2(n538), .ZN(n451) );
  XOR2_X1 U502 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n449) );
  XNOR2_X1 U503 ( .A(n449), .B(G176GAT), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n451), .B(n450), .ZN(G1349GAT) );
  NAND2_X1 U505 ( .A1(n545), .A2(n565), .ZN(n455) );
  XOR2_X1 U506 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n453) );
  INV_X1 U507 ( .A(G190GAT), .ZN(n452) );
  XNOR2_X1 U508 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n477) );
  OR2_X1 U509 ( .A1(n578), .A2(n551), .ZN(n456) );
  XNOR2_X1 U510 ( .A(n456), .B(KEYINPUT74), .ZN(n487) );
  XOR2_X1 U511 ( .A(n493), .B(KEYINPUT96), .Z(n457) );
  XNOR2_X1 U512 ( .A(KEYINPUT27), .B(n457), .ZN(n529) );
  XNOR2_X1 U513 ( .A(KEYINPUT28), .B(n464), .ZN(n536) );
  INV_X1 U514 ( .A(n533), .ZN(n497) );
  XNOR2_X1 U515 ( .A(KEYINPUT89), .B(n497), .ZN(n458) );
  NOR2_X1 U516 ( .A1(n536), .A2(n458), .ZN(n459) );
  NAND2_X1 U517 ( .A1(n529), .A2(n459), .ZN(n460) );
  NAND2_X1 U518 ( .A1(n530), .A2(n460), .ZN(n470) );
  NOR2_X1 U519 ( .A1(n493), .A2(n497), .ZN(n461) );
  NOR2_X1 U520 ( .A1(n464), .A2(n461), .ZN(n462) );
  XNOR2_X1 U521 ( .A(n462), .B(KEYINPUT97), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n463), .B(KEYINPUT25), .ZN(n467) );
  NAND2_X1 U523 ( .A1(n497), .A2(n464), .ZN(n465) );
  XOR2_X1 U524 ( .A(KEYINPUT26), .B(n465), .Z(n568) );
  AND2_X1 U525 ( .A1(n529), .A2(n568), .ZN(n466) );
  NOR2_X1 U526 ( .A1(n467), .A2(n466), .ZN(n468) );
  NAND2_X1 U527 ( .A1(n570), .A2(n468), .ZN(n469) );
  NAND2_X1 U528 ( .A1(n470), .A2(n469), .ZN(n484) );
  INV_X1 U529 ( .A(n484), .ZN(n474) );
  XOR2_X1 U530 ( .A(KEYINPUT16), .B(KEYINPUT82), .Z(n472) );
  NAND2_X1 U531 ( .A1(n581), .A2(n561), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n472), .B(n471), .ZN(n473) );
  NAND2_X1 U533 ( .A1(n474), .A2(n473), .ZN(n504) );
  NOR2_X1 U534 ( .A1(n487), .A2(n504), .ZN(n475) );
  XNOR2_X1 U535 ( .A(KEYINPUT98), .B(n475), .ZN(n482) );
  NAND2_X1 U536 ( .A1(n530), .A2(n482), .ZN(n476) );
  XNOR2_X1 U537 ( .A(n477), .B(n476), .ZN(G1324GAT) );
  XOR2_X1 U538 ( .A(G8GAT), .B(KEYINPUT99), .Z(n479) );
  INV_X1 U539 ( .A(n493), .ZN(n521) );
  NAND2_X1 U540 ( .A1(n482), .A2(n521), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n479), .B(n478), .ZN(G1325GAT) );
  XOR2_X1 U542 ( .A(G15GAT), .B(KEYINPUT35), .Z(n481) );
  NAND2_X1 U543 ( .A1(n533), .A2(n482), .ZN(n480) );
  XNOR2_X1 U544 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  NAND2_X1 U545 ( .A1(n482), .A2(n536), .ZN(n483) );
  XNOR2_X1 U546 ( .A(n483), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U547 ( .A1(n586), .A2(n484), .ZN(n485) );
  NAND2_X1 U548 ( .A1(n557), .A2(n485), .ZN(n486) );
  XOR2_X1 U549 ( .A(KEYINPUT37), .B(n486), .Z(n518) );
  NOR2_X1 U550 ( .A1(n487), .A2(n518), .ZN(n489) );
  XNOR2_X1 U551 ( .A(KEYINPUT38), .B(KEYINPUT101), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n489), .B(n488), .ZN(n501) );
  NOR2_X1 U553 ( .A1(n501), .A2(n570), .ZN(n492) );
  XNOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT100), .ZN(n490) );
  XNOR2_X1 U555 ( .A(n490), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U556 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  NOR2_X1 U557 ( .A1(n493), .A2(n501), .ZN(n494) );
  XOR2_X1 U558 ( .A(G36GAT), .B(n494), .Z(G1329GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT40), .B(KEYINPUT102), .Z(n496) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(KEYINPUT103), .ZN(n495) );
  XNOR2_X1 U561 ( .A(n496), .B(n495), .ZN(n499) );
  NOR2_X1 U562 ( .A1(n501), .A2(n497), .ZN(n498) );
  XOR2_X1 U563 ( .A(n499), .B(n498), .Z(G1330GAT) );
  INV_X1 U564 ( .A(n536), .ZN(n500) );
  NOR2_X1 U565 ( .A1(n501), .A2(n500), .ZN(n502) );
  XOR2_X1 U566 ( .A(G50GAT), .B(n502), .Z(n503) );
  XNOR2_X1 U567 ( .A(KEYINPUT104), .B(n503), .ZN(G1331GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT42), .B(KEYINPUT105), .Z(n506) );
  NAND2_X1 U569 ( .A1(n551), .A2(n538), .ZN(n517) );
  NOR2_X1 U570 ( .A1(n504), .A2(n517), .ZN(n512) );
  NAND2_X1 U571 ( .A1(n512), .A2(n530), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(n507), .ZN(G1332GAT) );
  NAND2_X1 U574 ( .A1(n521), .A2(n512), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n508), .B(KEYINPUT106), .ZN(n509) );
  XNOR2_X1 U576 ( .A(G64GAT), .B(n509), .ZN(G1333GAT) );
  XOR2_X1 U577 ( .A(G71GAT), .B(KEYINPUT107), .Z(n511) );
  NAND2_X1 U578 ( .A1(n512), .A2(n533), .ZN(n510) );
  XNOR2_X1 U579 ( .A(n511), .B(n510), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U581 ( .A1(n512), .A2(n536), .ZN(n513) );
  XNOR2_X1 U582 ( .A(n514), .B(n513), .ZN(n516) );
  XOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT108), .Z(n515) );
  XNOR2_X1 U584 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(KEYINPUT110), .ZN(n520) );
  NOR2_X1 U586 ( .A1(n518), .A2(n517), .ZN(n526) );
  NAND2_X1 U587 ( .A1(n526), .A2(n530), .ZN(n519) );
  XNOR2_X1 U588 ( .A(n520), .B(n519), .ZN(G1336GAT) );
  XOR2_X1 U589 ( .A(G92GAT), .B(KEYINPUT111), .Z(n523) );
  NAND2_X1 U590 ( .A1(n526), .A2(n521), .ZN(n522) );
  XNOR2_X1 U591 ( .A(n523), .B(n522), .ZN(G1337GAT) );
  NAND2_X1 U592 ( .A1(n526), .A2(n533), .ZN(n524) );
  XNOR2_X1 U593 ( .A(n524), .B(KEYINPUT112), .ZN(n525) );
  XNOR2_X1 U594 ( .A(G99GAT), .B(n525), .ZN(G1338GAT) );
  NAND2_X1 U595 ( .A1(n526), .A2(n536), .ZN(n527) );
  XNOR2_X1 U596 ( .A(n527), .B(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  NAND2_X1 U598 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U599 ( .A1(n532), .A2(n531), .ZN(n550) );
  NAND2_X1 U600 ( .A1(n533), .A2(n550), .ZN(n534) );
  XNOR2_X1 U601 ( .A(KEYINPUT114), .B(n534), .ZN(n535) );
  NOR2_X1 U602 ( .A1(n536), .A2(n535), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n573), .A2(n546), .ZN(n537) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U606 ( .A1(n546), .A2(n538), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U608 ( .A(G120GAT), .B(n541), .Z(G1341GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n543) );
  NAND2_X1 U610 ( .A1(n546), .A2(n581), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U612 ( .A(G127GAT), .B(n544), .Z(G1342GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U614 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U616 ( .A(G134GAT), .B(n549), .Z(G1343GAT) );
  NAND2_X1 U617 ( .A1(n550), .A2(n568), .ZN(n560) );
  NOR2_X1 U618 ( .A1(n551), .A2(n560), .ZN(n552) );
  XOR2_X1 U619 ( .A(G141GAT), .B(n552), .Z(G1344GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n560), .ZN(n555) );
  XNOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n556), .ZN(G1345GAT) );
  NOR2_X1 U624 ( .A1(n557), .A2(n560), .ZN(n558) );
  XOR2_X1 U625 ( .A(KEYINPUT118), .B(n558), .Z(n559) );
  XNOR2_X1 U626 ( .A(G155GAT), .B(n559), .ZN(G1346GAT) );
  NOR2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n563) );
  XNOR2_X1 U628 ( .A(G162GAT), .B(KEYINPUT119), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1347GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n573), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U632 ( .A(G183GAT), .B(KEYINPUT123), .Z(n567) );
  NAND2_X1 U633 ( .A1(n565), .A2(n581), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(G1350GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n575) );
  INV_X1 U636 ( .A(n568), .ZN(n572) );
  NAND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n584) );
  NAND2_X1 U639 ( .A1(n584), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n577) );
  XOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT60), .Z(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U644 ( .A1(n584), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NAND2_X1 U646 ( .A1(n581), .A2(n584), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(KEYINPUT126), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G211GAT), .B(n583), .ZN(G1354GAT) );
  INV_X1 U649 ( .A(n584), .ZN(n585) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n588) );
  XNOR2_X1 U651 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

