//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n810, new_n812, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009;
  INV_X1    g000(.A(G169gat), .ZN(new_n202));
  INV_X1    g001(.A(G176gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AOI21_X1  g003(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT26), .ZN(new_n208));
  AND3_X1   g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT66), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT66), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G190gat), .ZN(new_n213));
  INV_X1    g012(.A(G183gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT27), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT27), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G183gat), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n211), .A2(new_n213), .A3(new_n215), .A4(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT66), .B(G190gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT27), .B(G183gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n209), .A2(new_n220), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT23), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(G169gat), .B2(G176gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n227), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n207), .A2(KEYINPUT24), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT24), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n233), .A2(G183gat), .A3(G190gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n214), .A2(new_n210), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n231), .B1(new_n237), .B2(KEYINPUT65), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n232), .A2(new_n234), .B1(new_n214), .B2(new_n210), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT25), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n221), .A2(new_n214), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n235), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n227), .A2(new_n229), .A3(new_n230), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(KEYINPUT25), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n226), .B1(new_n242), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT71), .ZN(new_n249));
  INV_X1    g048(.A(G134gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G127gat), .ZN(new_n251));
  INV_X1    g050(.A(G127gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(G134gat), .ZN(new_n253));
  AND2_X1   g052(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n254));
  NOR2_X1   g053(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n251), .B(new_n253), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n257));
  INV_X1    g056(.A(G113gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n257), .B1(new_n258), .B2(G120gat), .ZN(new_n259));
  INV_X1    g058(.A(G120gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n260), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(G120gat), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n256), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G127gat), .B(G134gat), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n260), .A2(G113gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n258), .A2(G120gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n268), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n249), .B1(new_n267), .B2(new_n273), .ZN(new_n274));
  OR2_X1    g073(.A1(new_n254), .A2(new_n255), .ZN(new_n275));
  AND2_X1   g074(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n276), .A2(new_n263), .A3(new_n260), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n259), .A2(new_n261), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n268), .B(new_n275), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n272), .A2(new_n269), .ZN(new_n280));
  INV_X1    g079(.A(new_n268), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n279), .A2(KEYINPUT71), .A3(new_n282), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n248), .A2(KEYINPUT72), .A3(new_n274), .A4(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n285));
  NOR3_X1   g084(.A1(new_n267), .A2(new_n249), .A3(new_n273), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT71), .B1(new_n279), .B2(new_n282), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT25), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n245), .B1(new_n239), .B2(new_n240), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n235), .A2(new_n240), .A3(new_n236), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n225), .B1(new_n292), .B2(new_n246), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n274), .A2(KEYINPUT72), .A3(new_n283), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n288), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G227gat), .A2(G233gat), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n296), .B(KEYINPUT64), .Z(new_n297));
  NAND3_X1  g096(.A1(new_n284), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT32), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT33), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(G15gat), .B(G43gat), .Z(new_n302));
  XNOR2_X1  g101(.A(G71gat), .B(G99gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n299), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n304), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n298), .B(KEYINPUT32), .C1(new_n300), .C2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n284), .A2(new_n295), .ZN(new_n309));
  INV_X1    g108(.A(new_n297), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n311), .B(KEYINPUT34), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  OR2_X1    g112(.A1(new_n311), .A2(KEYINPUT34), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n311), .A2(KEYINPUT34), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n314), .A2(new_n305), .A3(new_n315), .A4(new_n307), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT86), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT81), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n319), .B1(G155gat), .B2(G162gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(G141gat), .B(G148gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT2), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n322), .B1(G155gat), .B2(G162gat), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n320), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G155gat), .B(G162gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  OR2_X1    g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(G141gat), .A2(G148gat), .ZN(new_n329));
  AND2_X1   g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n328), .B(new_n329), .C1(new_n330), .C2(new_n322), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(new_n325), .A3(new_n320), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT3), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT29), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  AND2_X1   g135(.A1(KEYINPUT76), .A2(G211gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(KEYINPUT76), .A2(G211gat), .ZN(new_n338));
  OAI21_X1  g137(.A(G218gat), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT75), .B(KEYINPUT22), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G204gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G197gat), .ZN(new_n343));
  INV_X1    g142(.A(G197gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G204gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n349));
  XNOR2_X1  g148(.A(G211gat), .B(G218gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n350), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n346), .B1(new_n339), .B2(new_n340), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n352), .B1(new_n353), .B2(KEYINPUT77), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n351), .A2(new_n354), .A3(KEYINPUT78), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT78), .B1(new_n351), .B2(new_n354), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n336), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n331), .A2(new_n325), .A3(new_n320), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n325), .B1(new_n331), .B2(new_n320), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n350), .B1(new_n348), .B2(new_n349), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n353), .A2(KEYINPUT77), .A3(new_n352), .ZN(new_n363));
  NOR3_X1   g162(.A1(new_n362), .A2(new_n363), .A3(KEYINPUT29), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n361), .B1(new_n364), .B2(KEYINPUT3), .ZN(new_n365));
  INV_X1    g164(.A(G228gat), .ZN(new_n366));
  INV_X1    g165(.A(G233gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n358), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n348), .A2(new_n350), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT29), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n352), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n333), .B1(new_n373), .B2(new_n334), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n368), .B1(new_n358), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(G22gat), .B1(new_n369), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n358), .A2(new_n365), .A3(new_n368), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT78), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n379), .B1(new_n362), .B2(new_n363), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n335), .B1(new_n380), .B2(new_n355), .ZN(new_n381));
  OAI22_X1  g180(.A1(new_n381), .A2(new_n374), .B1(new_n366), .B2(new_n367), .ZN(new_n382));
  INV_X1    g181(.A(G22gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n378), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(G78gat), .B(G106gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT31), .B(G50gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  AND4_X1   g186(.A1(new_n318), .A2(new_n377), .A3(new_n384), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n384), .A2(KEYINPUT86), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n389), .A2(new_n387), .B1(new_n377), .B2(new_n384), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n317), .A2(new_n391), .ZN(new_n392));
  NOR3_X1   g191(.A1(new_n267), .A2(KEYINPUT83), .A3(new_n273), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n394), .B1(new_n279), .B2(new_n282), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n334), .B1(new_n359), .B2(new_n360), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n327), .A2(KEYINPUT82), .A3(KEYINPUT3), .A4(new_n332), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n327), .A2(KEYINPUT3), .A3(new_n332), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT82), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n396), .A2(new_n397), .A3(new_n398), .A4(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n333), .A2(new_n282), .A3(new_n279), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT4), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT4), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n274), .A2(new_n405), .A3(new_n283), .A4(new_n333), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT5), .ZN(new_n408));
  NAND2_X1  g207(.A1(G225gat), .A2(G233gat), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n402), .A2(new_n407), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n274), .A2(KEYINPUT4), .A3(new_n283), .A4(new_n333), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n403), .A2(new_n405), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n402), .A2(new_n409), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT84), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT83), .B1(new_n267), .B2(new_n273), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n279), .A2(new_n394), .A3(new_n282), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(new_n361), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n403), .ZN(new_n418));
  INV_X1    g217(.A(new_n409), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n408), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n413), .A2(new_n414), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n414), .B1(new_n413), .B2(new_n420), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n410), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G1gat), .B(G29gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(KEYINPUT0), .ZN(new_n425));
  XNOR2_X1  g224(.A(G57gat), .B(G85gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n410), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n401), .A2(new_n398), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n397), .A2(new_n415), .A3(new_n416), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n409), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n412), .A2(new_n411), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT5), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT84), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n413), .A2(new_n414), .A3(new_n420), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n429), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n427), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT6), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n428), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n423), .A2(KEYINPUT6), .A3(new_n427), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT90), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n423), .A2(KEYINPUT90), .A3(KEYINPUT6), .A4(new_n427), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n443), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT35), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n380), .A2(new_n355), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(G226gat), .A2(G233gat), .ZN(new_n452));
  XOR2_X1   g251(.A(new_n452), .B(KEYINPUT79), .Z(new_n453));
  AOI21_X1  g252(.A(new_n453), .B1(new_n248), .B2(new_n371), .ZN(new_n454));
  INV_X1    g253(.A(new_n453), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n293), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n451), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n455), .B1(new_n293), .B2(KEYINPUT29), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n248), .A2(new_n453), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(new_n450), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G8gat), .B(G36gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(G64gat), .B(G92gat), .ZN(new_n463));
  XOR2_X1   g262(.A(new_n462), .B(new_n463), .Z(new_n464));
  OR2_X1    g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n461), .A2(KEYINPUT30), .A3(new_n464), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n461), .A2(new_n464), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT30), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT80), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT80), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n468), .A2(new_n472), .A3(new_n469), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n467), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n392), .A2(new_n448), .A3(new_n449), .A4(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT73), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n308), .A2(new_n312), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n316), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n477), .B1(new_n308), .B2(new_n312), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n479), .A2(new_n391), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT85), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n442), .B1(new_n439), .B2(new_n440), .ZN(new_n483));
  AOI211_X1 g282(.A(new_n427), .B(new_n429), .C1(new_n437), .C2(new_n438), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n428), .A2(new_n441), .A3(KEYINPUT85), .A4(new_n442), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(new_n486), .A3(new_n444), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n481), .A2(new_n487), .A3(new_n474), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT35), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n476), .B1(new_n489), .B2(KEYINPUT92), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT92), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n488), .A2(new_n491), .A3(KEYINPUT35), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT91), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT37), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n458), .A2(new_n450), .A3(new_n459), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n450), .B1(new_n458), .B2(new_n459), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT88), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT88), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n461), .A2(new_n499), .A3(new_n494), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT38), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n495), .A2(new_n496), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n464), .B1(new_n503), .B2(KEYINPUT37), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n501), .A2(KEYINPUT89), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n443), .A2(new_n446), .A3(new_n505), .A4(new_n447), .ZN(new_n506));
  INV_X1    g305(.A(new_n468), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n499), .B1(new_n461), .B2(new_n494), .ZN(new_n508));
  AOI211_X1 g307(.A(KEYINPUT88), .B(KEYINPUT37), .C1(new_n457), .C2(new_n460), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n504), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n507), .B1(new_n510), .B2(KEYINPUT38), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n504), .B(new_n502), .C1(new_n508), .C2(new_n509), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT89), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n506), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n391), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n409), .B1(new_n402), .B2(new_n407), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT39), .B1(new_n418), .B2(new_n419), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT39), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n427), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n522), .A3(KEYINPUT40), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT87), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT87), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n520), .A2(new_n522), .A3(new_n525), .A4(KEYINPUT40), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT40), .B1(new_n520), .B2(new_n522), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n528), .B1(new_n423), .B2(new_n427), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n517), .B1(new_n530), .B2(new_n474), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n493), .B1(new_n516), .B2(new_n531), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n527), .A2(new_n529), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n471), .A2(new_n473), .ZN(new_n534));
  INV_X1    g333(.A(new_n467), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n391), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n537), .B(KEYINPUT91), .C1(new_n515), .C2(new_n506), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n532), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n480), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n540), .A2(KEYINPUT36), .A3(new_n478), .A4(new_n316), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT36), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT74), .B1(new_n317), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT74), .ZN(new_n544));
  AOI211_X1 g343(.A(new_n544), .B(KEYINPUT36), .C1(new_n313), .C2(new_n316), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n487), .A2(new_n474), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n541), .A2(new_n546), .B1(new_n547), .B2(new_n391), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n490), .A2(new_n492), .B1(new_n539), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT101), .ZN(new_n550));
  XNOR2_X1  g349(.A(G43gat), .B(G50gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT15), .ZN(new_n552));
  INV_X1    g351(.A(G43gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(KEYINPUT93), .A3(G50gat), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT15), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT93), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n556), .B1(new_n557), .B2(new_n551), .ZN(new_n558));
  INV_X1    g357(.A(G29gat), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n559), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT14), .B(G29gat), .ZN(new_n561));
  INV_X1    g360(.A(G36gat), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n552), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n563), .A2(new_n552), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT94), .B(KEYINPUT17), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT95), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G15gat), .B(G22gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT16), .ZN(new_n572));
  AOI21_X1  g371(.A(G1gat), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT96), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n573), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT97), .B(G8gat), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT97), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n576), .B1(new_n579), .B2(G8gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n566), .A2(KEYINPUT17), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n570), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G229gat), .A2(G233gat), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n564), .A2(new_n565), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n584), .A2(KEYINPUT18), .A3(new_n585), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT99), .ZN(new_n589));
  AOI22_X1  g388(.A1(new_n570), .A2(new_n583), .B1(new_n586), .B2(new_n581), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT99), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n590), .A2(new_n591), .A3(KEYINPUT18), .A4(new_n585), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n578), .A2(new_n566), .A3(new_n580), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n585), .B(KEYINPUT13), .Z(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(KEYINPUT100), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n595), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT100), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n589), .A2(new_n592), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G113gat), .B(G141gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(G197gat), .ZN(new_n602));
  XOR2_X1   g401(.A(KEYINPUT11), .B(G169gat), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n604), .B(KEYINPUT12), .Z(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT18), .B1(new_n607), .B2(KEYINPUT98), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT98), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n590), .A2(new_n609), .A3(new_n585), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n600), .A2(new_n606), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n606), .B1(new_n600), .B2(new_n611), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n550), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n600), .A2(new_n611), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(new_n605), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n606), .A3(new_n611), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(KEYINPUT101), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n549), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT107), .ZN(new_n621));
  XOR2_X1   g420(.A(G134gat), .B(G162gat), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT104), .ZN(new_n623));
  AND2_X1   g422(.A1(G232gat), .A2(G233gat), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n624), .A2(KEYINPUT41), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n623), .B(new_n625), .Z(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(KEYINPUT41), .ZN(new_n627));
  NAND2_X1  g426(.A1(G85gat), .A2(G92gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT7), .ZN(new_n629));
  NAND2_X1  g428(.A1(G99gat), .A2(G106gat), .ZN(new_n630));
  INV_X1    g429(.A(G85gat), .ZN(new_n631));
  INV_X1    g430(.A(G92gat), .ZN(new_n632));
  AOI22_X1  g431(.A1(KEYINPUT8), .A2(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G99gat), .B(G106gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n634), .B(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n627), .B1(new_n637), .B2(new_n566), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n634), .B(new_n635), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n582), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n638), .B1(new_n570), .B2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G190gat), .B(G218gat), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n641), .A2(KEYINPUT105), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT105), .B1(new_n641), .B2(new_n643), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n621), .B(new_n626), .C1(new_n647), .C2(KEYINPUT106), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n641), .A2(new_n643), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT105), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(KEYINPUT106), .B1(new_n651), .B2(new_n644), .ZN(new_n652));
  INV_X1    g451(.A(new_n626), .ZN(new_n653));
  OAI21_X1  g452(.A(KEYINPUT107), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  OAI22_X1  g454(.A1(new_n645), .A2(new_n646), .B1(new_n643), .B2(new_n641), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n656), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n648), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G71gat), .B(G78gat), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT9), .ZN(new_n662));
  INV_X1    g461(.A(G71gat), .ZN(new_n663));
  INV_X1    g462(.A(G78gat), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(G64gat), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n667));
  INV_X1    g466(.A(G57gat), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(KEYINPUT103), .A2(G57gat), .A3(G64gat), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n661), .A2(new_n665), .A3(new_n669), .A4(new_n670), .ZN(new_n671));
  XOR2_X1   g470(.A(G71gat), .B(G78gat), .Z(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n666), .ZN(new_n673));
  NAND2_X1  g472(.A1(G57gat), .A2(G64gat), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(KEYINPUT9), .A3(new_n674), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n672), .A2(new_n675), .A3(KEYINPUT102), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT102), .B1(new_n672), .B2(new_n675), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n671), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT21), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(G231gat), .A2(G233gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G127gat), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n578), .B(new_n580), .C1(new_n679), .C2(new_n678), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n683), .B(new_n684), .Z(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(G155gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(G183gat), .B(G211gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n685), .B(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT10), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n637), .A2(new_n678), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT109), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n636), .A2(KEYINPUT108), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n678), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n639), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n637), .B1(new_n678), .B2(new_n694), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n693), .B1(new_n698), .B2(KEYINPUT10), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n696), .A2(new_n697), .A3(KEYINPUT109), .A4(new_n691), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n692), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(G230gat), .A2(G233gat), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n698), .A2(new_n703), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(G120gat), .B(G148gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(G176gat), .B(G204gat), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n707), .B(new_n708), .Z(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n706), .A2(KEYINPUT111), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT111), .B1(new_n706), .B2(new_n710), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n705), .B(new_n709), .C1(new_n701), .C2(new_n703), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT110), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n660), .A2(new_n690), .A3(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n620), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n487), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G1gat), .ZN(G1324gat));
  INV_X1    g523(.A(G8gat), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(new_n721), .B2(new_n536), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT16), .B(G8gat), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n720), .A2(new_n474), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT42), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n729), .B1(KEYINPUT42), .B2(new_n728), .ZN(G1325gat));
  INV_X1    g529(.A(new_n543), .ZN(new_n731));
  INV_X1    g530(.A(new_n545), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n731), .A2(new_n732), .A3(new_n541), .ZN(new_n733));
  OAI21_X1  g532(.A(G15gat), .B1(new_n720), .B2(new_n733), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n317), .A2(G15gat), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n720), .B2(new_n735), .ZN(G1326gat));
  NAND3_X1  g535(.A1(new_n721), .A2(KEYINPUT112), .A3(new_n391), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT112), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n720), .B2(new_n517), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(KEYINPUT43), .B(G22gat), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1327gat));
  INV_X1    g541(.A(new_n690), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n717), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(new_n660), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n620), .A2(new_n559), .A3(new_n722), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT45), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n549), .B2(new_n660), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n648), .A2(new_n654), .A3(new_n658), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n658), .B1(new_n648), .B2(new_n654), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n488), .A2(new_n491), .A3(KEYINPUT35), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n491), .B1(new_n488), .B2(KEYINPUT35), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n753), .A2(new_n754), .A3(new_n476), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n547), .A2(new_n391), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n733), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n757), .B1(new_n532), .B2(new_n538), .ZN(new_n758));
  OAI211_X1 g557(.A(KEYINPUT44), .B(new_n752), .C1(new_n755), .C2(new_n758), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n749), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n612), .A2(new_n613), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n744), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(new_n722), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT113), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G29gat), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n763), .A2(KEYINPUT113), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n747), .B1(new_n765), .B2(new_n766), .ZN(G1328gat));
  NAND2_X1  g566(.A1(new_n620), .A2(new_n745), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n768), .A2(G36gat), .A3(new_n474), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT46), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n760), .A2(new_n536), .A3(new_n762), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n562), .B2(new_n771), .ZN(G1329gat));
  INV_X1    g571(.A(new_n733), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n760), .A2(G43gat), .A3(new_n773), .A4(new_n762), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n553), .B1(new_n768), .B2(new_n317), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g576(.A1(new_n749), .A2(new_n391), .A3(new_n759), .A4(new_n762), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(G50gat), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n768), .A2(KEYINPUT114), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n517), .A2(G50gat), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n768), .A2(KEYINPUT114), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n779), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT48), .B1(new_n779), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n784), .B(new_n786), .ZN(G1331gat));
  NAND2_X1  g586(.A1(new_n489), .A2(KEYINPUT92), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n788), .A2(new_n492), .A3(new_n475), .ZN(new_n789));
  AND4_X1   g588(.A1(new_n443), .A2(new_n446), .A3(new_n505), .A4(new_n447), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n511), .A2(new_n514), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT91), .B1(new_n792), .B2(new_n537), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n516), .A2(new_n493), .A3(new_n531), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n548), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n789), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n616), .A2(new_n617), .ZN(new_n797));
  NOR4_X1   g596(.A1(new_n752), .A2(new_n717), .A3(new_n797), .A4(new_n743), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(new_n487), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(new_n668), .ZN(G1332gat));
  NOR2_X1   g600(.A1(new_n799), .A2(new_n474), .ZN(new_n802));
  NOR2_X1   g601(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n803));
  AND2_X1   g602(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n805), .B1(new_n802), .B2(new_n803), .ZN(G1333gat));
  OAI21_X1  g605(.A(G71gat), .B1(new_n799), .B2(new_n733), .ZN(new_n807));
  INV_X1    g606(.A(new_n317), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n663), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n807), .B1(new_n799), .B2(new_n809), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n810), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g610(.A1(new_n799), .A2(new_n517), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(new_n664), .ZN(G1335gat));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n797), .B2(new_n690), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n743), .A2(new_n761), .A3(KEYINPUT116), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(new_n717), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n760), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(G85gat), .B1(new_n820), .B2(new_n487), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n796), .A2(new_n752), .A3(new_n817), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(KEYINPUT51), .ZN(new_n823));
  INV_X1    g622(.A(new_n717), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n824), .A2(new_n722), .A3(new_n631), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n821), .B1(new_n823), .B2(new_n825), .ZN(G1336gat));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n749), .A2(new_n536), .A3(new_n759), .A4(new_n819), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(G92gat), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n717), .A2(G92gat), .A3(new_n474), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n827), .B(new_n829), .C1(new_n823), .C2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n833));
  AOI211_X1 g632(.A(new_n660), .B(new_n818), .C1(new_n789), .C2(new_n795), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n822), .A2(KEYINPUT117), .A3(KEYINPUT51), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n838), .A2(new_n830), .B1(G92gat), .B2(new_n828), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n832), .B1(new_n839), .B2(new_n827), .ZN(G1337gat));
  NOR2_X1   g639(.A1(new_n820), .A2(new_n733), .ZN(new_n841));
  XNOR2_X1  g640(.A(KEYINPUT118), .B(G99gat), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n824), .A2(new_n808), .A3(new_n842), .ZN(new_n843));
  OAI22_X1  g642(.A1(new_n841), .A2(new_n842), .B1(new_n823), .B2(new_n843), .ZN(G1338gat));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n749), .A2(new_n391), .A3(new_n759), .A4(new_n819), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(G106gat), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n717), .A2(G106gat), .A3(new_n517), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n845), .B(new_n847), .C1(new_n823), .C2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n836), .A2(new_n837), .A3(new_n848), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n847), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT119), .B1(new_n852), .B2(KEYINPUT53), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT119), .ZN(new_n854));
  AOI211_X1 g653(.A(new_n854), .B(new_n845), .C1(new_n851), .C2(new_n847), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n850), .B1(new_n853), .B2(new_n855), .ZN(G1339gat));
  NAND2_X1  g655(.A1(new_n701), .A2(new_n703), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n704), .A2(KEYINPUT54), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n701), .A2(new_n703), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n709), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n858), .A2(new_n861), .A3(KEYINPUT55), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n715), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n858), .A2(new_n861), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT55), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n865), .A2(KEYINPUT120), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT120), .B1(new_n865), .B2(new_n866), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n797), .B(new_n864), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n594), .A2(new_n595), .ZN(new_n870));
  XOR2_X1   g669(.A(new_n870), .B(KEYINPUT121), .Z(new_n871));
  NOR2_X1   g670(.A1(new_n590), .A2(new_n585), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n604), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n873), .A2(new_n617), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n713), .B2(new_n716), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n752), .B1(new_n869), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n657), .A2(new_n659), .A3(new_n874), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n864), .B1(new_n867), .B2(new_n868), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n743), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n718), .A2(new_n797), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n487), .A2(new_n536), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n392), .ZN(new_n886));
  OAI21_X1  g685(.A(G113gat), .B1(new_n886), .B2(new_n619), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n481), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n797), .A2(new_n264), .A3(new_n265), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(G1340gat));
  OAI21_X1  g689(.A(G120gat), .B1(new_n886), .B2(new_n717), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n824), .A2(new_n260), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT122), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n891), .B1(new_n888), .B2(new_n893), .ZN(G1341gat));
  OAI21_X1  g693(.A(G127gat), .B1(new_n886), .B2(new_n743), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n690), .A2(new_n252), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n888), .B2(new_n896), .ZN(G1342gat));
  NAND2_X1  g696(.A1(new_n752), .A2(new_n250), .ZN(new_n898));
  OR3_X1    g697(.A1(new_n888), .A2(KEYINPUT56), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(G134gat), .B1(new_n886), .B2(new_n660), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT56), .B1(new_n888), .B2(new_n898), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(G1343gat));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n869), .A2(new_n875), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n660), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n877), .A2(new_n878), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n690), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n903), .B(new_n391), .C1(new_n907), .C2(new_n881), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n733), .A2(new_n884), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n865), .A2(new_n866), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n614), .A2(new_n618), .A3(new_n864), .A4(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n752), .B1(new_n912), .B2(new_n875), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n743), .B1(new_n913), .B2(new_n879), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n517), .B1(new_n914), .B2(new_n882), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n908), .B(new_n910), .C1(new_n903), .C2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT123), .B1(new_n916), .B2(new_n619), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n912), .A2(new_n875), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n660), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n690), .B1(new_n919), .B2(new_n906), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n391), .B1(new_n920), .B2(new_n881), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n909), .B1(new_n921), .B2(KEYINPUT57), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n923));
  INV_X1    g722(.A(new_n619), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n922), .A2(new_n923), .A3(new_n924), .A4(new_n908), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n917), .A2(new_n925), .A3(G141gat), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n773), .A2(new_n517), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n885), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n619), .A2(G141gat), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT58), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(G141gat), .B1(new_n916), .B2(new_n761), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n928), .A2(new_n929), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(KEYINPUT58), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n931), .A2(new_n935), .ZN(G1344gat));
  INV_X1    g735(.A(G148gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n928), .A2(new_n937), .A3(new_n824), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT59), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n718), .A2(new_n924), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n903), .B(new_n391), .C1(new_n920), .C2(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n517), .B1(new_n880), .B2(new_n882), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(new_n903), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n910), .A2(new_n824), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n939), .B1(new_n945), .B2(G148gat), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n939), .A2(G148gat), .ZN(new_n947));
  INV_X1    g746(.A(new_n916), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n948), .B2(new_n824), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n938), .B1(new_n946), .B2(new_n949), .ZN(G1345gat));
  NAND3_X1  g749(.A1(new_n928), .A2(KEYINPUT124), .A3(new_n690), .ZN(new_n951));
  INV_X1    g750(.A(G155gat), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n885), .A2(new_n690), .A3(new_n927), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT124), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n951), .A2(new_n952), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n948), .A2(G155gat), .A3(new_n690), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n956), .A2(new_n957), .ZN(G1346gat));
  AOI21_X1  g757(.A(G162gat), .B1(new_n928), .B2(new_n752), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n752), .A2(G162gat), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n959), .B1(new_n948), .B2(new_n960), .ZN(G1347gat));
  NOR2_X1   g760(.A1(new_n722), .A2(new_n474), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n883), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(new_n392), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n964), .A2(new_n202), .A3(new_n619), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n883), .A2(new_n481), .A3(new_n962), .ZN(new_n966));
  AOI21_X1  g765(.A(G169gat), .B1(new_n966), .B2(new_n797), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n965), .A2(new_n967), .ZN(G1348gat));
  OAI21_X1  g767(.A(G176gat), .B1(new_n964), .B2(new_n717), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n966), .A2(new_n203), .A3(new_n824), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(G1349gat));
  OAI21_X1  g770(.A(G183gat), .B1(new_n964), .B2(new_n743), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n966), .A2(new_n222), .A3(new_n690), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(KEYINPUT60), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT60), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n972), .A2(new_n976), .A3(new_n973), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(new_n977), .ZN(G1350gat));
  NAND3_X1  g777(.A1(new_n966), .A2(new_n221), .A3(new_n752), .ZN(new_n979));
  NAND4_X1  g778(.A1(new_n883), .A2(new_n392), .A3(new_n752), .A4(new_n962), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT61), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n980), .A2(new_n981), .A3(G190gat), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n981), .B1(new_n980), .B2(G190gat), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n979), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g783(.A(new_n984), .B(KEYINPUT125), .ZN(G1351gat));
  AND2_X1   g784(.A1(new_n962), .A2(new_n733), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n942), .A2(new_n986), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n987), .A2(G197gat), .A3(new_n761), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT126), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n943), .A2(KEYINPUT127), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT127), .ZN(new_n991));
  OAI211_X1 g790(.A(new_n941), .B(new_n991), .C1(new_n903), .C2(new_n942), .ZN(new_n992));
  AND4_X1   g791(.A1(new_n924), .A2(new_n990), .A3(new_n992), .A4(new_n986), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n989), .B1(new_n993), .B2(new_n344), .ZN(G1352gat));
  NOR3_X1   g793(.A1(new_n987), .A2(G204gat), .A3(new_n717), .ZN(new_n995));
  XNOR2_X1  g794(.A(new_n995), .B(KEYINPUT62), .ZN(new_n996));
  AND4_X1   g795(.A1(new_n824), .A2(new_n990), .A3(new_n992), .A4(new_n986), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n996), .B1(new_n997), .B2(new_n342), .ZN(G1353gat));
  OR4_X1    g797(.A1(new_n338), .A2(new_n987), .A3(new_n337), .A4(new_n743), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n986), .A2(new_n690), .ZN(new_n1000));
  OAI21_X1  g799(.A(G211gat), .B1(new_n943), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT63), .ZN(new_n1002));
  AND2_X1   g801(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n999), .B1(new_n1003), .B2(new_n1004), .ZN(G1354gat));
  INV_X1    g804(.A(G218gat), .ZN(new_n1006));
  NOR2_X1   g805(.A1(new_n660), .A2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g806(.A1(new_n990), .A2(new_n992), .A3(new_n986), .A4(new_n1007), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1006), .B1(new_n987), .B2(new_n660), .ZN(new_n1009));
  AND2_X1   g808(.A1(new_n1008), .A2(new_n1009), .ZN(G1355gat));
endmodule


