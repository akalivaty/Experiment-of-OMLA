

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U553 ( .A1(n694), .A2(G40), .ZN(n784) );
  NOR2_X2 U554 ( .A1(n575), .A2(n574), .ZN(n694) );
  NOR2_X1 U555 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U556 ( .A1(G168), .A2(n702), .ZN(n703) );
  XNOR2_X2 U557 ( .A(n698), .B(n697), .ZN(n747) );
  NOR2_X1 U558 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U559 ( .A(n566), .B(n565), .ZN(n570) );
  XNOR2_X2 U560 ( .A(n568), .B(n567), .ZN(n624) );
  OR2_X1 U561 ( .A1(n780), .A2(n776), .ZN(n520) );
  XNOR2_X1 U562 ( .A(n596), .B(KEYINPUT13), .ZN(n521) );
  AND2_X1 U563 ( .A1(G8), .A2(n742), .ZN(n522) );
  XOR2_X1 U564 ( .A(n771), .B(KEYINPUT100), .Z(n523) );
  BUF_X1 U565 ( .A(n709), .Z(n748) );
  INV_X1 U566 ( .A(KEYINPUT32), .ZN(n755) );
  XNOR2_X1 U567 ( .A(n756), .B(n755), .ZN(n757) );
  NAND2_X1 U568 ( .A1(n785), .A2(n696), .ZN(n709) );
  NAND2_X1 U569 ( .A1(n520), .A2(n781), .ZN(n782) );
  XNOR2_X1 U570 ( .A(n564), .B(KEYINPUT23), .ZN(n565) );
  NOR2_X2 U571 ( .A1(G2104), .A2(n571), .ZN(n894) );
  AND2_X2 U572 ( .A1(n571), .A2(G2104), .ZN(n888) );
  NOR2_X1 U573 ( .A1(G651), .A2(n662), .ZN(n657) );
  XOR2_X1 U574 ( .A(KEYINPUT1), .B(n525), .Z(n661) );
  NOR2_X2 U575 ( .A1(n600), .A2(n599), .ZN(n948) );
  XNOR2_X1 U576 ( .A(G543), .B(KEYINPUT0), .ZN(n524) );
  XOR2_X1 U577 ( .A(n524), .B(KEYINPUT68), .Z(n662) );
  NAND2_X1 U578 ( .A1(G51), .A2(n657), .ZN(n527) );
  INV_X1 U579 ( .A(G651), .ZN(n530) );
  NOR2_X1 U580 ( .A1(G543), .A2(n530), .ZN(n525) );
  NAND2_X1 U581 ( .A1(G63), .A2(n661), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U583 ( .A(KEYINPUT6), .B(n528), .ZN(n537) );
  NOR2_X1 U584 ( .A1(G543), .A2(G651), .ZN(n650) );
  NAND2_X1 U585 ( .A1(n650), .A2(G89), .ZN(n529) );
  XNOR2_X1 U586 ( .A(n529), .B(KEYINPUT4), .ZN(n533) );
  OR2_X1 U587 ( .A1(n530), .A2(n662), .ZN(n531) );
  XNOR2_X2 U588 ( .A(KEYINPUT69), .B(n531), .ZN(n649) );
  NAND2_X1 U589 ( .A1(G76), .A2(n649), .ZN(n532) );
  NAND2_X1 U590 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U591 ( .A(KEYINPUT74), .B(n534), .Z(n535) );
  XNOR2_X1 U592 ( .A(KEYINPUT5), .B(n535), .ZN(n536) );
  NOR2_X1 U593 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U594 ( .A(KEYINPUT7), .B(n538), .Z(G168) );
  XOR2_X1 U595 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U596 ( .A1(G91), .A2(n650), .ZN(n540) );
  NAND2_X1 U597 ( .A1(G78), .A2(n649), .ZN(n539) );
  NAND2_X1 U598 ( .A1(n540), .A2(n539), .ZN(n544) );
  NAND2_X1 U599 ( .A1(G53), .A2(n657), .ZN(n542) );
  NAND2_X1 U600 ( .A1(G65), .A2(n661), .ZN(n541) );
  NAND2_X1 U601 ( .A1(n542), .A2(n541), .ZN(n543) );
  OR2_X1 U602 ( .A1(n544), .A2(n543), .ZN(G299) );
  NAND2_X1 U603 ( .A1(G52), .A2(n657), .ZN(n546) );
  NAND2_X1 U604 ( .A1(G64), .A2(n661), .ZN(n545) );
  NAND2_X1 U605 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U606 ( .A(KEYINPUT70), .B(n547), .ZN(n553) );
  NAND2_X1 U607 ( .A1(G90), .A2(n650), .ZN(n549) );
  NAND2_X1 U608 ( .A1(G77), .A2(n649), .ZN(n548) );
  NAND2_X1 U609 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U610 ( .A(KEYINPUT9), .B(n550), .ZN(n551) );
  XNOR2_X1 U611 ( .A(KEYINPUT71), .B(n551), .ZN(n552) );
  NOR2_X1 U612 ( .A1(n553), .A2(n552), .ZN(G171) );
  XOR2_X1 U613 ( .A(G2446), .B(G2430), .Z(n555) );
  XNOR2_X1 U614 ( .A(G2451), .B(G2454), .ZN(n554) );
  XNOR2_X1 U615 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U616 ( .A(n556), .B(G2427), .Z(n558) );
  XNOR2_X1 U617 ( .A(G1348), .B(G1341), .ZN(n557) );
  XNOR2_X1 U618 ( .A(n558), .B(n557), .ZN(n562) );
  XOR2_X1 U619 ( .A(G2443), .B(KEYINPUT104), .Z(n560) );
  XNOR2_X1 U620 ( .A(G2438), .B(G2435), .ZN(n559) );
  XNOR2_X1 U621 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U622 ( .A(n562), .B(n561), .Z(n563) );
  AND2_X1 U623 ( .A1(G14), .A2(n563), .ZN(G401) );
  AND2_X1 U624 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U625 ( .A(G57), .ZN(G237) );
  INV_X1 U626 ( .A(G108), .ZN(G238) );
  INV_X1 U627 ( .A(G120), .ZN(G236) );
  NAND2_X1 U628 ( .A1(G101), .A2(n888), .ZN(n566) );
  INV_X1 U629 ( .A(KEYINPUT66), .ZN(n564) );
  XNOR2_X1 U630 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n568) );
  NOR2_X1 U631 ( .A1(G2104), .A2(G2105), .ZN(n567) );
  NAND2_X1 U632 ( .A1(G137), .A2(n624), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n575) );
  INV_X1 U634 ( .A(G2105), .ZN(n571) );
  AND2_X1 U635 ( .A1(G2104), .A2(G2105), .ZN(n892) );
  NAND2_X1 U636 ( .A1(G113), .A2(n892), .ZN(n573) );
  NAND2_X1 U637 ( .A1(G125), .A2(n894), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  BUF_X1 U639 ( .A(n694), .Z(G160) );
  NAND2_X1 U640 ( .A1(G88), .A2(n650), .ZN(n577) );
  NAND2_X1 U641 ( .A1(G75), .A2(n649), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(KEYINPUT78), .B(n578), .ZN(n582) );
  NAND2_X1 U644 ( .A1(G50), .A2(n657), .ZN(n580) );
  NAND2_X1 U645 ( .A1(G62), .A2(n661), .ZN(n579) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U647 ( .A1(n582), .A2(n581), .ZN(G166) );
  NAND2_X1 U648 ( .A1(G114), .A2(n892), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n583), .B(KEYINPUT84), .ZN(n586) );
  NAND2_X1 U650 ( .A1(G102), .A2(n888), .ZN(n584) );
  XOR2_X1 U651 ( .A(KEYINPUT85), .B(n584), .Z(n585) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n590) );
  NAND2_X1 U653 ( .A1(G126), .A2(n894), .ZN(n588) );
  NAND2_X1 U654 ( .A1(G138), .A2(n624), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U656 ( .A1(n590), .A2(n589), .ZN(G164) );
  NAND2_X1 U657 ( .A1(G7), .A2(G661), .ZN(n591) );
  XNOR2_X1 U658 ( .A(n591), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U659 ( .A(G223), .ZN(n835) );
  NAND2_X1 U660 ( .A1(n835), .A2(G567), .ZN(n592) );
  XOR2_X1 U661 ( .A(KEYINPUT11), .B(n592), .Z(G234) );
  NAND2_X1 U662 ( .A1(n650), .A2(G81), .ZN(n593) );
  XNOR2_X1 U663 ( .A(n593), .B(KEYINPUT12), .ZN(n595) );
  NAND2_X1 U664 ( .A1(G68), .A2(n649), .ZN(n594) );
  NAND2_X1 U665 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U666 ( .A1(G43), .A2(n657), .ZN(n597) );
  NAND2_X1 U667 ( .A1(n521), .A2(n597), .ZN(n600) );
  NAND2_X1 U668 ( .A1(n661), .A2(G56), .ZN(n598) );
  XOR2_X1 U669 ( .A(KEYINPUT14), .B(n598), .Z(n599) );
  NAND2_X1 U670 ( .A1(n948), .A2(G860), .ZN(G153) );
  NAND2_X1 U671 ( .A1(G868), .A2(G171), .ZN(n610) );
  NAND2_X1 U672 ( .A1(n657), .A2(G54), .ZN(n607) );
  NAND2_X1 U673 ( .A1(G92), .A2(n650), .ZN(n602) );
  NAND2_X1 U674 ( .A1(G79), .A2(n649), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n602), .A2(n601), .ZN(n605) );
  NAND2_X1 U676 ( .A1(n661), .A2(G66), .ZN(n603) );
  XOR2_X1 U677 ( .A(KEYINPUT72), .B(n603), .Z(n604) );
  NOR2_X1 U678 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X2 U680 ( .A(KEYINPUT15), .B(n608), .Z(n951) );
  INV_X1 U681 ( .A(n951), .ZN(n631) );
  INV_X1 U682 ( .A(G868), .ZN(n675) );
  NAND2_X1 U683 ( .A1(n631), .A2(n675), .ZN(n609) );
  NAND2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U685 ( .A(n611), .B(KEYINPUT73), .ZN(G284) );
  NOR2_X1 U686 ( .A1(G286), .A2(n675), .ZN(n613) );
  NOR2_X1 U687 ( .A1(G868), .A2(G299), .ZN(n612) );
  NOR2_X1 U688 ( .A1(n613), .A2(n612), .ZN(G297) );
  INV_X1 U689 ( .A(G860), .ZN(n633) );
  NAND2_X1 U690 ( .A1(G559), .A2(n633), .ZN(n614) );
  XOR2_X1 U691 ( .A(KEYINPUT75), .B(n614), .Z(n615) );
  NAND2_X1 U692 ( .A1(n615), .A2(n631), .ZN(n616) );
  XNOR2_X1 U693 ( .A(n616), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U694 ( .A1(n631), .A2(G868), .ZN(n617) );
  NOR2_X1 U695 ( .A1(G559), .A2(n617), .ZN(n619) );
  AND2_X1 U696 ( .A1(n675), .A2(n948), .ZN(n618) );
  NOR2_X1 U697 ( .A1(n619), .A2(n618), .ZN(G282) );
  NAND2_X1 U698 ( .A1(G123), .A2(n894), .ZN(n620) );
  XNOR2_X1 U699 ( .A(n620), .B(KEYINPUT76), .ZN(n621) );
  XNOR2_X1 U700 ( .A(n621), .B(KEYINPUT18), .ZN(n623) );
  NAND2_X1 U701 ( .A1(G111), .A2(n892), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n628) );
  NAND2_X1 U703 ( .A1(G99), .A2(n888), .ZN(n626) );
  NAND2_X1 U704 ( .A1(G135), .A2(n624), .ZN(n625) );
  NAND2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n997) );
  XNOR2_X1 U707 ( .A(G2096), .B(n997), .ZN(n630) );
  INV_X1 U708 ( .A(G2100), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n630), .A2(n629), .ZN(G156) );
  NAND2_X1 U710 ( .A1(G559), .A2(n631), .ZN(n632) );
  XNOR2_X1 U711 ( .A(n632), .B(n948), .ZN(n672) );
  NAND2_X1 U712 ( .A1(n633), .A2(n672), .ZN(n640) );
  NAND2_X1 U713 ( .A1(G55), .A2(n657), .ZN(n635) );
  NAND2_X1 U714 ( .A1(G67), .A2(n661), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U716 ( .A1(G93), .A2(n650), .ZN(n637) );
  NAND2_X1 U717 ( .A1(G80), .A2(n649), .ZN(n636) );
  NAND2_X1 U718 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U719 ( .A1(n639), .A2(n638), .ZN(n674) );
  XOR2_X1 U720 ( .A(n640), .B(n674), .Z(G145) );
  NAND2_X1 U721 ( .A1(G86), .A2(n650), .ZN(n642) );
  NAND2_X1 U722 ( .A1(G61), .A2(n661), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U724 ( .A1(G73), .A2(n649), .ZN(n643) );
  XNOR2_X1 U725 ( .A(n643), .B(KEYINPUT77), .ZN(n644) );
  XNOR2_X1 U726 ( .A(n644), .B(KEYINPUT2), .ZN(n645) );
  NOR2_X1 U727 ( .A1(n646), .A2(n645), .ZN(n648) );
  NAND2_X1 U728 ( .A1(n657), .A2(G48), .ZN(n647) );
  NAND2_X1 U729 ( .A1(n648), .A2(n647), .ZN(G305) );
  AND2_X1 U730 ( .A1(n649), .A2(G72), .ZN(n654) );
  NAND2_X1 U731 ( .A1(G85), .A2(n650), .ZN(n652) );
  NAND2_X1 U732 ( .A1(G47), .A2(n657), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U734 ( .A1(n654), .A2(n653), .ZN(n656) );
  NAND2_X1 U735 ( .A1(n661), .A2(G60), .ZN(n655) );
  NAND2_X1 U736 ( .A1(n656), .A2(n655), .ZN(G290) );
  NAND2_X1 U737 ( .A1(G49), .A2(n657), .ZN(n659) );
  NAND2_X1 U738 ( .A1(G74), .A2(G651), .ZN(n658) );
  NAND2_X1 U739 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U740 ( .A1(n661), .A2(n660), .ZN(n664) );
  NAND2_X1 U741 ( .A1(G87), .A2(n662), .ZN(n663) );
  NAND2_X1 U742 ( .A1(n664), .A2(n663), .ZN(G288) );
  XOR2_X1 U743 ( .A(G290), .B(G299), .Z(n665) );
  XNOR2_X1 U744 ( .A(G305), .B(n665), .ZN(n669) );
  XNOR2_X1 U745 ( .A(KEYINPUT79), .B(KEYINPUT80), .ZN(n667) );
  XNOR2_X1 U746 ( .A(G288), .B(KEYINPUT19), .ZN(n666) );
  XNOR2_X1 U747 ( .A(n667), .B(n666), .ZN(n668) );
  XOR2_X1 U748 ( .A(n669), .B(n668), .Z(n671) );
  XNOR2_X1 U749 ( .A(G166), .B(n674), .ZN(n670) );
  XNOR2_X1 U750 ( .A(n671), .B(n670), .ZN(n905) );
  XOR2_X1 U751 ( .A(n905), .B(n672), .Z(n673) );
  NOR2_X1 U752 ( .A1(n675), .A2(n673), .ZN(n677) );
  AND2_X1 U753 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U754 ( .A1(n677), .A2(n676), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2078), .A2(G2084), .ZN(n678) );
  XOR2_X1 U756 ( .A(KEYINPUT20), .B(n678), .Z(n679) );
  NAND2_X1 U757 ( .A1(G2090), .A2(n679), .ZN(n680) );
  XNOR2_X1 U758 ( .A(KEYINPUT21), .B(n680), .ZN(n681) );
  NAND2_X1 U759 ( .A1(n681), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U760 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U761 ( .A1(G236), .A2(G238), .ZN(n682) );
  NAND2_X1 U762 ( .A1(G69), .A2(n682), .ZN(n683) );
  NOR2_X1 U763 ( .A1(n683), .A2(G237), .ZN(n684) );
  XNOR2_X1 U764 ( .A(n684), .B(KEYINPUT83), .ZN(n839) );
  NAND2_X1 U765 ( .A1(n839), .A2(G567), .ZN(n691) );
  XOR2_X1 U766 ( .A(KEYINPUT22), .B(KEYINPUT81), .Z(n686) );
  NAND2_X1 U767 ( .A1(G132), .A2(G82), .ZN(n685) );
  XNOR2_X1 U768 ( .A(n686), .B(n685), .ZN(n687) );
  NOR2_X1 U769 ( .A1(n687), .A2(G218), .ZN(n688) );
  XNOR2_X1 U770 ( .A(KEYINPUT82), .B(n688), .ZN(n689) );
  NAND2_X1 U771 ( .A1(n689), .A2(G96), .ZN(n840) );
  NAND2_X1 U772 ( .A1(n840), .A2(G2106), .ZN(n690) );
  NAND2_X1 U773 ( .A1(n691), .A2(n690), .ZN(n841) );
  NAND2_X1 U774 ( .A1(G661), .A2(G483), .ZN(n692) );
  NOR2_X1 U775 ( .A1(n841), .A2(n692), .ZN(n838) );
  NAND2_X1 U776 ( .A1(n838), .A2(G36), .ZN(G176) );
  INV_X1 U777 ( .A(G166), .ZN(G303) );
  INV_X1 U778 ( .A(G171), .ZN(G301) );
  XOR2_X1 U779 ( .A(G1981), .B(KEYINPUT101), .Z(n693) );
  XNOR2_X1 U780 ( .A(G305), .B(n693), .ZN(n946) );
  NOR2_X1 U781 ( .A1(G164), .A2(G1384), .ZN(n785) );
  INV_X1 U782 ( .A(KEYINPUT90), .ZN(n695) );
  XNOR2_X1 U783 ( .A(n695), .B(n784), .ZN(n696) );
  NAND2_X1 U784 ( .A1(n709), .A2(G8), .ZN(n698) );
  INV_X1 U785 ( .A(KEYINPUT91), .ZN(n697) );
  NOR2_X1 U786 ( .A1(G1966), .A2(n747), .ZN(n743) );
  NOR2_X1 U787 ( .A1(G2084), .A2(n748), .ZN(n742) );
  NOR2_X1 U788 ( .A1(n743), .A2(n742), .ZN(n699) );
  XNOR2_X1 U789 ( .A(n699), .B(KEYINPUT96), .ZN(n700) );
  NAND2_X1 U790 ( .A1(n700), .A2(G8), .ZN(n701) );
  XNOR2_X1 U791 ( .A(n701), .B(KEYINPUT30), .ZN(n702) );
  XNOR2_X1 U792 ( .A(n703), .B(KEYINPUT97), .ZN(n707) );
  XOR2_X1 U793 ( .A(G2078), .B(KEYINPUT25), .Z(n926) );
  NOR2_X1 U794 ( .A1(n926), .A2(n748), .ZN(n705) );
  INV_X1 U795 ( .A(n709), .ZN(n721) );
  NOR2_X1 U796 ( .A1(n721), .A2(G1961), .ZN(n704) );
  NOR2_X1 U797 ( .A1(n705), .A2(n704), .ZN(n737) );
  NAND2_X1 U798 ( .A1(n737), .A2(G301), .ZN(n706) );
  NAND2_X1 U799 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U800 ( .A(n708), .B(KEYINPUT31), .ZN(n741) );
  INV_X1 U801 ( .A(G1996), .ZN(n923) );
  NOR2_X1 U802 ( .A1(n709), .A2(n923), .ZN(n711) );
  XOR2_X1 U803 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n710) );
  XNOR2_X1 U804 ( .A(n711), .B(n710), .ZN(n713) );
  NAND2_X1 U805 ( .A1(n748), .A2(G1341), .ZN(n712) );
  NAND2_X1 U806 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U807 ( .A(KEYINPUT93), .B(n714), .ZN(n715) );
  NAND2_X1 U808 ( .A1(n715), .A2(n948), .ZN(n716) );
  XNOR2_X1 U809 ( .A(n716), .B(KEYINPUT65), .ZN(n720) );
  NAND2_X1 U810 ( .A1(G1348), .A2(n748), .ZN(n718) );
  NAND2_X1 U811 ( .A1(G2067), .A2(n721), .ZN(n717) );
  NAND2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n726) );
  NAND2_X1 U813 ( .A1(n726), .A2(n951), .ZN(n719) );
  NAND2_X1 U814 ( .A1(n720), .A2(n719), .ZN(n730) );
  NAND2_X1 U815 ( .A1(n721), .A2(G2072), .ZN(n722) );
  XOR2_X1 U816 ( .A(KEYINPUT27), .B(n722), .Z(n724) );
  NAND2_X1 U817 ( .A1(G1956), .A2(n748), .ZN(n723) );
  NAND2_X1 U818 ( .A1(n724), .A2(n723), .ZN(n732) );
  NOR2_X1 U819 ( .A1(G299), .A2(n732), .ZN(n725) );
  XNOR2_X1 U820 ( .A(n725), .B(KEYINPUT94), .ZN(n728) );
  NOR2_X1 U821 ( .A1(n951), .A2(n726), .ZN(n727) );
  NOR2_X1 U822 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U823 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U824 ( .A(KEYINPUT95), .B(n731), .ZN(n735) );
  NAND2_X1 U825 ( .A1(G299), .A2(n732), .ZN(n733) );
  XOR2_X1 U826 ( .A(KEYINPUT28), .B(n733), .Z(n734) );
  XNOR2_X1 U827 ( .A(n736), .B(KEYINPUT29), .ZN(n739) );
  OR2_X1 U828 ( .A1(G301), .A2(n737), .ZN(n738) );
  NAND2_X1 U829 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U830 ( .A1(n741), .A2(n740), .ZN(n746) );
  NOR2_X1 U831 ( .A1(n743), .A2(n522), .ZN(n744) );
  NAND2_X1 U832 ( .A1(n746), .A2(n744), .ZN(n745) );
  XOR2_X1 U833 ( .A(KEYINPUT98), .B(n745), .Z(n758) );
  NAND2_X1 U834 ( .A1(n746), .A2(G286), .ZN(n753) );
  INV_X1 U835 ( .A(n747), .ZN(n780) );
  NOR2_X1 U836 ( .A1(G1971), .A2(n747), .ZN(n750) );
  NOR2_X1 U837 ( .A1(G2090), .A2(n748), .ZN(n749) );
  NOR2_X1 U838 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U839 ( .A1(n751), .A2(G303), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U841 ( .A1(G8), .A2(n754), .ZN(n756) );
  XNOR2_X1 U842 ( .A(n759), .B(KEYINPUT99), .ZN(n772) );
  NOR2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n761) );
  NOR2_X1 U844 ( .A1(G1971), .A2(G303), .ZN(n760) );
  NOR2_X1 U845 ( .A1(n761), .A2(n760), .ZN(n959) );
  NAND2_X1 U846 ( .A1(n761), .A2(n780), .ZN(n762) );
  NAND2_X1 U847 ( .A1(n762), .A2(KEYINPUT33), .ZN(n764) );
  AND2_X1 U848 ( .A1(n959), .A2(n764), .ZN(n763) );
  NAND2_X1 U849 ( .A1(n772), .A2(n763), .ZN(n770) );
  INV_X1 U850 ( .A(n764), .ZN(n768) );
  NAND2_X1 U851 ( .A1(G1976), .A2(G288), .ZN(n954) );
  INV_X1 U852 ( .A(KEYINPUT33), .ZN(n765) );
  NAND2_X1 U853 ( .A1(n954), .A2(n765), .ZN(n766) );
  NOR2_X1 U854 ( .A1(n766), .A2(n747), .ZN(n767) );
  OR2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n769) );
  AND2_X1 U856 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U857 ( .A1(n946), .A2(n523), .ZN(n783) );
  INV_X1 U858 ( .A(n772), .ZN(n775) );
  NAND2_X1 U859 ( .A1(G8), .A2(G166), .ZN(n773) );
  NOR2_X1 U860 ( .A1(G2090), .A2(n773), .ZN(n774) );
  NOR2_X1 U861 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U862 ( .A1(G1981), .A2(G305), .ZN(n777) );
  XNOR2_X1 U863 ( .A(n777), .B(KEYINPUT24), .ZN(n778) );
  XNOR2_X1 U864 ( .A(n778), .B(KEYINPUT92), .ZN(n779) );
  NAND2_X1 U865 ( .A1(n780), .A2(n779), .ZN(n781) );
  OR2_X1 U866 ( .A1(n783), .A2(n782), .ZN(n818) );
  XNOR2_X1 U867 ( .A(G1986), .B(G290), .ZN(n957) );
  NOR2_X1 U868 ( .A1(n785), .A2(n784), .ZN(n829) );
  NAND2_X1 U869 ( .A1(n957), .A2(n829), .ZN(n816) );
  NAND2_X1 U870 ( .A1(G95), .A2(n888), .ZN(n787) );
  NAND2_X1 U871 ( .A1(G131), .A2(n624), .ZN(n786) );
  NAND2_X1 U872 ( .A1(n787), .A2(n786), .ZN(n791) );
  NAND2_X1 U873 ( .A1(G107), .A2(n892), .ZN(n789) );
  NAND2_X1 U874 ( .A1(G119), .A2(n894), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U876 ( .A1(n791), .A2(n790), .ZN(n882) );
  INV_X1 U877 ( .A(G1991), .ZN(n920) );
  NOR2_X1 U878 ( .A1(n882), .A2(n920), .ZN(n801) );
  NAND2_X1 U879 ( .A1(G141), .A2(n624), .ZN(n792) );
  XNOR2_X1 U880 ( .A(n792), .B(KEYINPUT88), .ZN(n799) );
  NAND2_X1 U881 ( .A1(G117), .A2(n892), .ZN(n794) );
  NAND2_X1 U882 ( .A1(G129), .A2(n894), .ZN(n793) );
  NAND2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U884 ( .A1(n888), .A2(G105), .ZN(n795) );
  XOR2_X1 U885 ( .A(KEYINPUT38), .B(n795), .Z(n796) );
  NOR2_X1 U886 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U887 ( .A1(n799), .A2(n798), .ZN(n878) );
  AND2_X1 U888 ( .A1(n878), .A2(G1996), .ZN(n800) );
  NOR2_X1 U889 ( .A1(n801), .A2(n800), .ZN(n1003) );
  INV_X1 U890 ( .A(n829), .ZN(n802) );
  NOR2_X1 U891 ( .A1(n1003), .A2(n802), .ZN(n822) );
  XNOR2_X1 U892 ( .A(KEYINPUT89), .B(n822), .ZN(n814) );
  XNOR2_X1 U893 ( .A(G2067), .B(KEYINPUT37), .ZN(n803) );
  XNOR2_X1 U894 ( .A(n803), .B(KEYINPUT86), .ZN(n819) );
  NAND2_X1 U895 ( .A1(n624), .A2(G140), .ZN(n804) );
  XOR2_X1 U896 ( .A(KEYINPUT87), .B(n804), .Z(n806) );
  NAND2_X1 U897 ( .A1(n888), .A2(G104), .ZN(n805) );
  NAND2_X1 U898 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U899 ( .A(KEYINPUT34), .B(n807), .ZN(n812) );
  NAND2_X1 U900 ( .A1(G116), .A2(n892), .ZN(n809) );
  NAND2_X1 U901 ( .A1(G128), .A2(n894), .ZN(n808) );
  NAND2_X1 U902 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U903 ( .A(KEYINPUT35), .B(n810), .Z(n811) );
  NOR2_X1 U904 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U905 ( .A(KEYINPUT36), .B(n813), .ZN(n883) );
  NOR2_X1 U906 ( .A1(n819), .A2(n883), .ZN(n1019) );
  NAND2_X1 U907 ( .A1(n829), .A2(n1019), .ZN(n826) );
  AND2_X1 U908 ( .A1(n814), .A2(n826), .ZN(n815) );
  AND2_X1 U909 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U910 ( .A1(n818), .A2(n817), .ZN(n832) );
  NAND2_X1 U911 ( .A1(n819), .A2(n883), .ZN(n1016) );
  NOR2_X1 U912 ( .A1(G1996), .A2(n878), .ZN(n1000) );
  AND2_X1 U913 ( .A1(n920), .A2(n882), .ZN(n998) );
  NOR2_X1 U914 ( .A1(G1986), .A2(G290), .ZN(n820) );
  NOR2_X1 U915 ( .A1(n998), .A2(n820), .ZN(n821) );
  NOR2_X1 U916 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U917 ( .A1(n1000), .A2(n823), .ZN(n824) );
  XNOR2_X1 U918 ( .A(KEYINPUT102), .B(n824), .ZN(n825) );
  XNOR2_X1 U919 ( .A(n825), .B(KEYINPUT39), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U921 ( .A1(n1016), .A2(n828), .ZN(n830) );
  NAND2_X1 U922 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U923 ( .A1(n832), .A2(n831), .ZN(n834) );
  XOR2_X1 U924 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n833) );
  XNOR2_X1 U925 ( .A(n834), .B(n833), .ZN(G329) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n835), .ZN(G217) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n836) );
  NAND2_X1 U928 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U930 ( .A1(n838), .A2(n837), .ZN(G188) );
  INV_X1 U932 ( .A(G132), .ZN(G219) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  INV_X1 U934 ( .A(G82), .ZN(G220) );
  NOR2_X1 U935 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  INV_X1 U937 ( .A(n841), .ZN(G319) );
  XOR2_X1 U938 ( .A(G2678), .B(G2084), .Z(n843) );
  XNOR2_X1 U939 ( .A(G2090), .B(G2078), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U941 ( .A(n844), .B(G2096), .Z(n846) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2072), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U944 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n848) );
  XNOR2_X1 U945 ( .A(KEYINPUT42), .B(G2100), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U947 ( .A(n850), .B(n849), .Z(G227) );
  XOR2_X1 U948 ( .A(G1956), .B(G1986), .Z(n852) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n862) );
  XOR2_X1 U951 ( .A(KEYINPUT106), .B(KEYINPUT41), .Z(n854) );
  XNOR2_X1 U952 ( .A(G1981), .B(G2474), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U954 ( .A(G1976), .B(G1971), .Z(n856) );
  XNOR2_X1 U955 ( .A(G1966), .B(G1961), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U957 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U958 ( .A(KEYINPUT108), .B(KEYINPUT107), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(G229) );
  NAND2_X1 U961 ( .A1(G124), .A2(n894), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n863), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U963 ( .A1(n892), .A2(G112), .ZN(n864) );
  NAND2_X1 U964 ( .A1(n865), .A2(n864), .ZN(n869) );
  NAND2_X1 U965 ( .A1(G100), .A2(n888), .ZN(n867) );
  NAND2_X1 U966 ( .A1(G136), .A2(n624), .ZN(n866) );
  NAND2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U968 ( .A1(n869), .A2(n868), .ZN(G162) );
  NAND2_X1 U969 ( .A1(G115), .A2(n892), .ZN(n871) );
  NAND2_X1 U970 ( .A1(G127), .A2(n894), .ZN(n870) );
  NAND2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n872), .B(KEYINPUT47), .ZN(n874) );
  NAND2_X1 U973 ( .A1(G103), .A2(n888), .ZN(n873) );
  NAND2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n877) );
  NAND2_X1 U975 ( .A1(G139), .A2(n624), .ZN(n875) );
  XNOR2_X1 U976 ( .A(KEYINPUT111), .B(n875), .ZN(n876) );
  NOR2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n1010) );
  XOR2_X1 U978 ( .A(n878), .B(n1010), .Z(n887) );
  XOR2_X1 U979 ( .A(KEYINPUT48), .B(KEYINPUT112), .Z(n880) );
  XNOR2_X1 U980 ( .A(G160), .B(KEYINPUT46), .ZN(n879) );
  XNOR2_X1 U981 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U982 ( .A(n997), .B(n881), .ZN(n885) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n903) );
  NAND2_X1 U986 ( .A1(G106), .A2(n888), .ZN(n890) );
  NAND2_X1 U987 ( .A1(G142), .A2(n624), .ZN(n889) );
  NAND2_X1 U988 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U989 ( .A(n891), .B(KEYINPUT45), .ZN(n899) );
  NAND2_X1 U990 ( .A1(n892), .A2(G118), .ZN(n893) );
  XOR2_X1 U991 ( .A(KEYINPUT109), .B(n893), .Z(n896) );
  NAND2_X1 U992 ( .A1(n894), .A2(G130), .ZN(n895) );
  NAND2_X1 U993 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U994 ( .A(KEYINPUT110), .B(n897), .Z(n898) );
  NAND2_X1 U995 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n900), .B(G162), .ZN(n901) );
  XNOR2_X1 U997 ( .A(G164), .B(n901), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U999 ( .A1(G37), .A2(n904), .ZN(G395) );
  XNOR2_X1 U1000 ( .A(n948), .B(G286), .ZN(n906) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n908) );
  XOR2_X1 U1002 ( .A(n951), .B(G171), .Z(n907) );
  XNOR2_X1 U1003 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n909), .ZN(G397) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1008 ( .A(KEYINPUT49), .B(n912), .Z(n913) );
  NOR2_X1 U1009 ( .A1(G401), .A2(n913), .ZN(n914) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n914), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(KEYINPUT115), .B(n915), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1016 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n1027) );
  INV_X1 U1017 ( .A(KEYINPUT55), .ZN(n1021) );
  XOR2_X1 U1018 ( .A(KEYINPUT122), .B(G34), .Z(n919) );
  XNOR2_X1 U1019 ( .A(G2084), .B(KEYINPUT54), .ZN(n918) );
  XNOR2_X1 U1020 ( .A(n919), .B(n918), .ZN(n940) );
  XNOR2_X1 U1021 ( .A(n920), .B(G25), .ZN(n921) );
  NAND2_X1 U1022 ( .A1(n921), .A2(G28), .ZN(n922) );
  XNOR2_X1 U1023 ( .A(n922), .B(KEYINPUT119), .ZN(n930) );
  XOR2_X1 U1024 ( .A(G2067), .B(G26), .Z(n925) );
  XNOR2_X1 U1025 ( .A(n923), .B(G32), .ZN(n924) );
  NAND2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(G27), .B(n926), .ZN(n927) );
  NOR2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(KEYINPUT120), .B(G2072), .ZN(n931) );
  XNOR2_X1 U1031 ( .A(G33), .B(n931), .ZN(n932) );
  NOR2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1033 ( .A(n934), .B(KEYINPUT53), .Z(n935) );
  XNOR2_X1 U1034 ( .A(KEYINPUT121), .B(n935), .ZN(n938) );
  XNOR2_X1 U1035 ( .A(KEYINPUT118), .B(G2090), .ZN(n936) );
  XNOR2_X1 U1036 ( .A(G35), .B(n936), .ZN(n937) );
  NOR2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1039 ( .A(n1021), .B(n941), .ZN(n943) );
  INV_X1 U1040 ( .A(G29), .ZN(n942) );
  NAND2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1042 ( .A1(G11), .A2(n944), .ZN(n996) );
  XNOR2_X1 U1043 ( .A(G16), .B(KEYINPUT56), .ZN(n968) );
  XOR2_X1 U1044 ( .A(G168), .B(G1966), .Z(n945) );
  NOR2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1046 ( .A(KEYINPUT57), .B(n947), .Z(n966) );
  XOR2_X1 U1047 ( .A(n948), .B(G1341), .Z(n964) );
  XNOR2_X1 U1048 ( .A(G1961), .B(G171), .ZN(n950) );
  NAND2_X1 U1049 ( .A1(G1971), .A2(G303), .ZN(n949) );
  NAND2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n961) );
  XNOR2_X1 U1051 ( .A(n951), .B(G1348), .ZN(n953) );
  XNOR2_X1 U1052 ( .A(G299), .B(G1956), .ZN(n952) );
  NOR2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n955) );
  NAND2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1058 ( .A(KEYINPUT123), .B(n962), .ZN(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n994) );
  INV_X1 U1062 ( .A(G16), .ZN(n992) );
  XOR2_X1 U1063 ( .A(G1986), .B(KEYINPUT124), .Z(n969) );
  XNOR2_X1 U1064 ( .A(G24), .B(n969), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(G1971), .B(G22), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(G23), .B(G1976), .ZN(n970) );
  NOR2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(n974), .B(KEYINPUT58), .ZN(n975) );
  XNOR2_X1 U1070 ( .A(KEYINPUT125), .B(n975), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(G1966), .B(G21), .ZN(n977) );
  XNOR2_X1 U1072 ( .A(G5), .B(G1961), .ZN(n976) );
  NOR2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n989) );
  XOR2_X1 U1075 ( .A(G1348), .B(KEYINPUT59), .Z(n980) );
  XNOR2_X1 U1076 ( .A(G4), .B(n980), .ZN(n982) );
  XNOR2_X1 U1077 ( .A(G20), .B(G1956), .ZN(n981) );
  NOR2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(G1341), .B(G19), .ZN(n984) );
  XNOR2_X1 U1080 ( .A(G6), .B(G1981), .ZN(n983) );
  NOR2_X1 U1081 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1082 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1083 ( .A(KEYINPUT60), .B(n987), .ZN(n988) );
  NOR2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1085 ( .A(KEYINPUT61), .B(n990), .ZN(n991) );
  NAND2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n1025) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n1009) );
  XOR2_X1 U1090 ( .A(G2090), .B(G162), .Z(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(n1001), .B(KEYINPUT117), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(n1002), .B(KEYINPUT51), .ZN(n1004) );
  NAND2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1007) );
  XOR2_X1 U1095 ( .A(G2084), .B(G160), .Z(n1005) );
  XNOR2_X1 U1096 ( .A(KEYINPUT116), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1015) );
  XOR2_X1 U1099 ( .A(G2072), .B(n1010), .Z(n1012) );
  XOR2_X1 U1100 ( .A(G164), .B(G2078), .Z(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1102 ( .A(KEYINPUT50), .B(n1013), .Z(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1106 ( .A(KEYINPUT52), .B(n1020), .ZN(n1022) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(G29), .ZN(n1024) );
  NAND2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1110 ( .A(n1027), .B(n1026), .ZN(G311) );
  XNOR2_X1 U1111 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

