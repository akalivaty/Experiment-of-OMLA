

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742;

  XNOR2_X1 U376 ( .A(G146), .B(G125), .ZN(n465) );
  XNOR2_X1 U377 ( .A(n424), .B(G953), .ZN(n728) );
  XNOR2_X2 U378 ( .A(n578), .B(n577), .ZN(n739) );
  AND2_X1 U379 ( .A1(n419), .A2(n418), .ZN(n417) );
  OR2_X2 U380 ( .A1(n372), .A2(n371), .ZN(n593) );
  NAND2_X1 U381 ( .A1(n549), .A2(n548), .ZN(n644) );
  XNOR2_X1 U382 ( .A(n485), .B(n484), .ZN(n548) );
  XNOR2_X1 U383 ( .A(n474), .B(n355), .ZN(n594) );
  XNOR2_X1 U384 ( .A(n501), .B(n500), .ZN(n542) );
  XNOR2_X1 U385 ( .A(n698), .B(n697), .ZN(n699) );
  AND2_X1 U386 ( .A1(n728), .A2(G224), .ZN(n423) );
  INV_X2 U387 ( .A(KEYINPUT4), .ZN(n427) );
  XNOR2_X1 U388 ( .A(n726), .B(G146), .ZN(n370) );
  XNOR2_X1 U389 ( .A(n538), .B(KEYINPUT1), .ZN(n655) );
  XNOR2_X1 U390 ( .A(n506), .B(n507), .ZN(n726) );
  AND2_X1 U391 ( .A1(G227), .A2(n728), .ZN(n437) );
  NAND2_X1 U392 ( .A1(n610), .A2(G472), .ZN(n373) );
  OR2_X1 U393 ( .A1(n604), .A2(G902), .ZN(n518) );
  XNOR2_X1 U394 ( .A(n443), .B(G107), .ZN(n515) );
  XNOR2_X1 U395 ( .A(G104), .B(G110), .ZN(n443) );
  XNOR2_X1 U396 ( .A(n589), .B(KEYINPUT22), .ZN(n595) );
  INV_X1 U397 ( .A(KEYINPUT44), .ZN(n431) );
  AND2_X1 U398 ( .A1(n435), .A2(KEYINPUT44), .ZN(n433) );
  NOR2_X1 U399 ( .A1(n737), .A2(n391), .ZN(n390) );
  NOR2_X1 U400 ( .A1(G953), .A2(G237), .ZN(n508) );
  XNOR2_X1 U401 ( .A(n398), .B(n397), .ZN(n677) );
  INV_X1 U402 ( .A(KEYINPUT45), .ZN(n397) );
  NAND2_X1 U403 ( .A1(n402), .A2(n399), .ZN(n398) );
  OR2_X1 U404 ( .A1(n596), .A2(n380), .ZN(n558) );
  NAND2_X1 U405 ( .A1(n521), .A2(n381), .ZN(n380) );
  NOR2_X1 U406 ( .A1(n571), .A2(n361), .ZN(n415) );
  XNOR2_X1 U407 ( .A(n368), .B(n367), .ZN(n502) );
  XNOR2_X1 U408 ( .A(n369), .B(G119), .ZN(n367) );
  INV_X1 U409 ( .A(KEYINPUT3), .ZN(n369) );
  XNOR2_X1 U410 ( .A(n466), .B(KEYINPUT90), .ZN(n394) );
  XNOR2_X1 U411 ( .A(KEYINPUT91), .B(KEYINPUT24), .ZN(n466) );
  XOR2_X1 U412 ( .A(G137), .B(G128), .Z(n469) );
  XNOR2_X1 U413 ( .A(G119), .B(G110), .ZN(n467) );
  XNOR2_X1 U414 ( .A(G116), .B(G107), .ZN(n478) );
  XOR2_X1 U415 ( .A(KEYINPUT9), .B(G122), .Z(n479) );
  XOR2_X1 U416 ( .A(KEYINPUT101), .B(KEYINPUT7), .Z(n480) );
  XNOR2_X1 U417 ( .A(n483), .B(G134), .ZN(n506) );
  XNOR2_X1 U418 ( .A(n406), .B(n405), .ZN(n517) );
  XNOR2_X1 U419 ( .A(n437), .B(G101), .ZN(n405) );
  XNOR2_X1 U420 ( .A(n574), .B(n573), .ZN(n672) );
  XNOR2_X1 U421 ( .A(KEYINPUT86), .B(KEYINPUT33), .ZN(n573) );
  XNOR2_X1 U422 ( .A(n554), .B(n553), .ZN(n565) );
  BUF_X1 U423 ( .A(n655), .Z(n382) );
  NAND2_X1 U424 ( .A1(n373), .A2(n376), .ZN(n372) );
  NAND2_X1 U425 ( .A1(G902), .A2(G472), .ZN(n376) );
  NOR2_X1 U426 ( .A1(n705), .A2(G902), .ZN(n485) );
  AND2_X1 U427 ( .A1(n356), .A2(n430), .ZN(n429) );
  NAND2_X1 U428 ( .A1(KEYINPUT65), .A2(n431), .ZN(n430) );
  NOR2_X1 U429 ( .A1(n739), .A2(KEYINPUT44), .ZN(n599) );
  NOR2_X1 U430 ( .A1(G237), .A2(G902), .ZN(n448) );
  XNOR2_X1 U431 ( .A(n389), .B(KEYINPUT46), .ZN(n388) );
  NOR2_X1 U432 ( .A1(n742), .A2(n741), .ZN(n389) );
  XNOR2_X1 U433 ( .A(G101), .B(G116), .ZN(n366) );
  XOR2_X1 U434 ( .A(KEYINPUT23), .B(G140), .Z(n468) );
  XOR2_X1 U435 ( .A(G131), .B(G140), .Z(n514) );
  NAND2_X1 U436 ( .A1(G234), .A2(G237), .ZN(n453) );
  NAND2_X1 U437 ( .A1(n587), .A2(KEYINPUT104), .ZN(n411) );
  NOR2_X1 U438 ( .A1(n587), .A2(KEYINPUT104), .ZN(n412) );
  AND2_X1 U439 ( .A1(n594), .A2(n395), .ZN(n521) );
  AND2_X1 U440 ( .A1(n651), .A2(n396), .ZN(n395) );
  INV_X1 U441 ( .A(n539), .ZN(n396) );
  NAND2_X1 U442 ( .A1(n378), .A2(n375), .ZN(n374) );
  INV_X1 U443 ( .A(G472), .ZN(n375) );
  XNOR2_X1 U444 ( .A(n510), .B(n511), .ZN(n610) );
  XNOR2_X1 U445 ( .A(n370), .B(n509), .ZN(n510) );
  XNOR2_X1 U446 ( .A(G113), .B(G143), .ZN(n488) );
  XNOR2_X1 U447 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n490) );
  XOR2_X1 U448 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n491) );
  XOR2_X1 U449 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n495) );
  INV_X1 U450 ( .A(KEYINPUT64), .ZN(n424) );
  NOR2_X1 U451 ( .A1(n672), .A2(n583), .ZN(n386) );
  AND2_X1 U452 ( .A1(n593), .A2(n641), .ZN(n537) );
  XNOR2_X1 U453 ( .A(n499), .B(G475), .ZN(n500) );
  NOR2_X1 U454 ( .A1(G902), .A2(n698), .ZN(n501) );
  INV_X1 U455 ( .A(n593), .ZN(n654) );
  XOR2_X1 U456 ( .A(G122), .B(KEYINPUT16), .Z(n444) );
  NOR2_X1 U457 ( .A1(n678), .A2(G953), .ZN(n713) );
  XNOR2_X1 U458 ( .A(n392), .B(n473), .ZN(n707) );
  XNOR2_X1 U459 ( .A(n471), .B(n393), .ZN(n392) );
  XNOR2_X1 U460 ( .A(n486), .B(n394), .ZN(n393) );
  XNOR2_X1 U461 ( .A(n384), .B(n383), .ZN(n705) );
  XNOR2_X1 U462 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U463 ( .A(n604), .B(n603), .ZN(n605) );
  XNOR2_X1 U464 ( .A(n520), .B(KEYINPUT109), .ZN(n737) );
  NOR2_X1 U465 ( .A1(n551), .A2(n523), .ZN(n625) );
  XNOR2_X1 U466 ( .A(n592), .B(n422), .ZN(n421) );
  INV_X1 U467 ( .A(KEYINPUT105), .ZN(n422) );
  INV_X1 U468 ( .A(n632), .ZN(n381) );
  NAND2_X1 U469 ( .A1(n417), .A2(n414), .ZN(n588) );
  XOR2_X1 U470 ( .A(n464), .B(n463), .Z(n355) );
  AND2_X1 U471 ( .A1(n591), .A2(n618), .ZN(n356) );
  AND2_X1 U472 ( .A1(n593), .A2(n521), .ZN(n357) );
  NOR2_X2 U473 ( .A1(n595), .A2(n382), .ZN(n592) );
  XNOR2_X1 U474 ( .A(KEYINPUT28), .B(n357), .ZN(n358) );
  AND2_X1 U475 ( .A1(n644), .A2(KEYINPUT104), .ZN(n359) );
  NAND2_X1 U476 ( .A1(n529), .A2(KEYINPUT47), .ZN(n360) );
  XNOR2_X1 U477 ( .A(KEYINPUT85), .B(KEYINPUT0), .ZN(n361) );
  INV_X1 U478 ( .A(KEYINPUT65), .ZN(n435) );
  XNOR2_X2 U479 ( .A(n362), .B(KEYINPUT32), .ZN(n740) );
  OR2_X1 U480 ( .A1(n595), .A2(n363), .ZN(n362) );
  NAND2_X1 U481 ( .A1(n597), .A2(n594), .ZN(n363) );
  XNOR2_X2 U482 ( .A(n364), .B(n522), .ZN(n572) );
  NOR2_X1 U483 ( .A1(n512), .A2(n364), .ZN(n513) );
  NAND2_X1 U484 ( .A1(n535), .A2(n641), .ZN(n364) );
  NAND2_X1 U485 ( .A1(n365), .A2(n433), .ZN(n432) );
  NOR2_X1 U486 ( .A1(n365), .A2(n435), .ZN(n434) );
  XNOR2_X1 U487 ( .A(n365), .B(KEYINPUT81), .ZN(n400) );
  XNOR2_X2 U488 ( .A(n598), .B(KEYINPUT82), .ZN(n365) );
  XNOR2_X1 U489 ( .A(n442), .B(n366), .ZN(n368) );
  XNOR2_X1 U490 ( .A(n517), .B(n370), .ZN(n604) );
  NOR2_X1 U491 ( .A1(n610), .A2(n374), .ZN(n371) );
  XNOR2_X2 U492 ( .A(n593), .B(KEYINPUT6), .ZN(n596) );
  XNOR2_X1 U493 ( .A(n377), .B(n423), .ZN(n446) );
  XNOR2_X1 U494 ( .A(n425), .B(n441), .ZN(n377) );
  INV_X1 U495 ( .A(G902), .ZN(n378) );
  NAND2_X1 U496 ( .A1(n379), .A2(n411), .ZN(n410) );
  NAND2_X1 U497 ( .A1(n413), .A2(n412), .ZN(n379) );
  INV_X2 U498 ( .A(G143), .ZN(n426) );
  NAND2_X1 U499 ( .A1(n740), .A2(n624), .ZN(n598) );
  XNOR2_X1 U500 ( .A(n516), .B(n515), .ZN(n406) );
  NAND2_X1 U501 ( .A1(n477), .A2(G217), .ZN(n383) );
  XNOR2_X1 U502 ( .A(n506), .B(n482), .ZN(n384) );
  NAND2_X1 U503 ( .A1(n385), .A2(n575), .ZN(n578) );
  XNOR2_X1 U504 ( .A(n386), .B(KEYINPUT34), .ZN(n385) );
  NAND2_X1 U505 ( .A1(n678), .A2(n679), .ZN(n680) );
  NAND2_X1 U506 ( .A1(n678), .A2(n682), .ZN(n683) );
  XNOR2_X1 U507 ( .A(n387), .B(KEYINPUT48), .ZN(n564) );
  NAND2_X1 U508 ( .A1(n390), .A2(n388), .ZN(n387) );
  NAND2_X1 U509 ( .A1(n547), .A2(n360), .ZN(n391) );
  NAND2_X1 U510 ( .A1(n401), .A2(n400), .ZN(n399) );
  XNOR2_X1 U511 ( .A(n599), .B(KEYINPUT66), .ZN(n401) );
  AND2_X1 U512 ( .A1(n403), .A2(n404), .ZN(n402) );
  XNOR2_X1 U513 ( .A(n579), .B(KEYINPUT80), .ZN(n403) );
  NOR2_X1 U514 ( .A1(n428), .A2(n434), .ZN(n404) );
  AND2_X1 U515 ( .A1(n541), .A2(n540), .ZN(n408) );
  NAND2_X1 U516 ( .A1(n407), .A2(n541), .ZN(n554) );
  AND2_X1 U517 ( .A1(n540), .A2(n642), .ZN(n407) );
  NAND2_X1 U518 ( .A1(n408), .A2(n575), .ZN(n543) );
  NOR2_X1 U519 ( .A1(n712), .A2(n613), .ZN(n616) );
  NOR2_X1 U520 ( .A1(n712), .A2(n695), .ZN(n696) );
  NOR2_X1 U521 ( .A1(n712), .A2(n701), .ZN(n702) );
  XNOR2_X1 U522 ( .A(n600), .B(KEYINPUT2), .ZN(n602) );
  NAND2_X1 U523 ( .A1(n588), .A2(n409), .ZN(n589) );
  NOR2_X1 U524 ( .A1(n410), .A2(n359), .ZN(n409) );
  INV_X1 U525 ( .A(n644), .ZN(n413) );
  NAND2_X1 U526 ( .A1(n416), .A2(n415), .ZN(n414) );
  INV_X1 U527 ( .A(n572), .ZN(n416) );
  NAND2_X1 U528 ( .A1(n571), .A2(n361), .ZN(n418) );
  NAND2_X1 U529 ( .A1(n572), .A2(n361), .ZN(n419) );
  NAND2_X1 U530 ( .A1(n421), .A2(n420), .ZN(n624) );
  NOR2_X1 U531 ( .A1(n593), .A2(n650), .ZN(n420) );
  XNOR2_X1 U532 ( .A(n483), .B(n505), .ZN(n425) );
  XNOR2_X2 U533 ( .A(n426), .B(G128), .ZN(n483) );
  XNOR2_X2 U534 ( .A(n427), .B(KEYINPUT68), .ZN(n505) );
  NAND2_X1 U535 ( .A1(n432), .A2(n429), .ZN(n428) );
  NOR2_X1 U536 ( .A1(n607), .A2(n712), .ZN(n609) );
  BUF_X1 U537 ( .A(n703), .Z(n708) );
  XNOR2_X1 U538 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U539 ( .A(KEYINPUT110), .B(KEYINPUT62), .ZN(n436) );
  XOR2_X1 U540 ( .A(n693), .B(n692), .Z(n438) );
  INV_X1 U541 ( .A(KEYINPUT71), .ZN(n461) );
  XNOR2_X1 U542 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U543 ( .A(n514), .B(n487), .ZN(n724) );
  XNOR2_X1 U544 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U545 ( .A(n515), .B(n444), .ZN(n445) );
  XNOR2_X1 U546 ( .A(n502), .B(n445), .ZN(n720) );
  XNOR2_X1 U547 ( .A(n614), .B(KEYINPUT63), .ZN(n615) );
  NOR2_X1 U548 ( .A1(n728), .A2(G952), .ZN(n712) );
  XNOR2_X2 U549 ( .A(G902), .B(KEYINPUT15), .ZN(n439) );
  XNOR2_X2 U550 ( .A(n439), .B(KEYINPUT88), .ZN(n601) );
  INV_X1 U551 ( .A(n601), .ZN(n447) );
  XNOR2_X1 U552 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n440) );
  XNOR2_X1 U553 ( .A(n465), .B(n440), .ZN(n441) );
  XNOR2_X1 U554 ( .A(G113), .B(KEYINPUT69), .ZN(n442) );
  XNOR2_X1 U555 ( .A(n720), .B(n446), .ZN(n691) );
  NOR2_X1 U556 ( .A1(n447), .A2(n691), .ZN(n450) );
  XOR2_X1 U557 ( .A(KEYINPUT70), .B(n448), .Z(n451) );
  NAND2_X1 U558 ( .A1(n451), .A2(G210), .ZN(n449) );
  XNOR2_X1 U559 ( .A(n450), .B(n449), .ZN(n535) );
  NAND2_X1 U560 ( .A1(G214), .A2(n451), .ZN(n452) );
  XNOR2_X1 U561 ( .A(n452), .B(KEYINPUT89), .ZN(n559) );
  INV_X1 U562 ( .A(n559), .ZN(n641) );
  XNOR2_X1 U563 ( .A(n453), .B(KEYINPUT14), .ZN(n454) );
  NAND2_X1 U564 ( .A1(G952), .A2(n454), .ZN(n670) );
  NOR2_X1 U565 ( .A1(G953), .A2(n670), .ZN(n570) );
  NAND2_X1 U566 ( .A1(G902), .A2(n454), .ZN(n568) );
  NOR2_X1 U567 ( .A1(n728), .A2(n568), .ZN(n455) );
  XOR2_X1 U568 ( .A(KEYINPUT106), .B(n455), .Z(n456) );
  NOR2_X1 U569 ( .A1(G900), .A2(n456), .ZN(n457) );
  NOR2_X1 U570 ( .A1(n570), .A2(n457), .ZN(n539) );
  XOR2_X1 U571 ( .A(KEYINPUT25), .B(KEYINPUT93), .Z(n460) );
  NAND2_X1 U572 ( .A1(n601), .A2(G234), .ZN(n458) );
  XNOR2_X1 U573 ( .A(KEYINPUT20), .B(n458), .ZN(n475) );
  NAND2_X1 U574 ( .A1(n475), .A2(G217), .ZN(n459) );
  XNOR2_X1 U575 ( .A(n460), .B(n459), .ZN(n464) );
  XNOR2_X1 U576 ( .A(KEYINPUT92), .B(KEYINPUT94), .ZN(n462) );
  XNOR2_X1 U577 ( .A(KEYINPUT10), .B(n465), .ZN(n486) );
  XOR2_X1 U578 ( .A(n468), .B(n467), .Z(n470) );
  NAND2_X1 U579 ( .A1(n728), .A2(G234), .ZN(n472) );
  XOR2_X1 U580 ( .A(KEYINPUT8), .B(n472), .Z(n477) );
  NAND2_X1 U581 ( .A1(G221), .A2(n477), .ZN(n473) );
  NOR2_X1 U582 ( .A1(G902), .A2(n707), .ZN(n474) );
  NAND2_X1 U583 ( .A1(n475), .A2(G221), .ZN(n476) );
  XOR2_X1 U584 ( .A(KEYINPUT21), .B(n476), .Z(n651) );
  XNOR2_X1 U585 ( .A(n479), .B(n478), .ZN(n481) );
  XNOR2_X1 U586 ( .A(KEYINPUT102), .B(G478), .ZN(n484) );
  INV_X1 U587 ( .A(n486), .ZN(n487) );
  XOR2_X1 U588 ( .A(G122), .B(G104), .Z(n489) );
  XNOR2_X1 U589 ( .A(n489), .B(n488), .ZN(n493) );
  XNOR2_X1 U590 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U591 ( .A(n492), .B(n493), .ZN(n497) );
  NAND2_X1 U592 ( .A1(G214), .A2(n508), .ZN(n494) );
  XNOR2_X1 U593 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U594 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U595 ( .A(n724), .B(n498), .ZN(n698) );
  XNOR2_X1 U596 ( .A(KEYINPUT100), .B(KEYINPUT13), .ZN(n499) );
  NAND2_X1 U597 ( .A1(n548), .A2(n542), .ZN(n632) );
  XOR2_X1 U598 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n504) );
  XNOR2_X1 U599 ( .A(n502), .B(G131), .ZN(n503) );
  XNOR2_X1 U600 ( .A(n504), .B(n503), .ZN(n511) );
  XNOR2_X1 U601 ( .A(G137), .B(n505), .ZN(n507) );
  NAND2_X1 U602 ( .A1(n508), .A2(G210), .ZN(n509) );
  XNOR2_X1 U603 ( .A(n558), .B(KEYINPUT108), .ZN(n512) );
  XNOR2_X1 U604 ( .A(KEYINPUT36), .B(n513), .ZN(n519) );
  XOR2_X1 U605 ( .A(KEYINPUT72), .B(n514), .Z(n516) );
  XNOR2_X2 U606 ( .A(n518), .B(G469), .ZN(n538) );
  NAND2_X1 U607 ( .A1(n519), .A2(n382), .ZN(n520) );
  NAND2_X1 U608 ( .A1(n358), .A2(n538), .ZN(n551) );
  INV_X1 U609 ( .A(KEYINPUT19), .ZN(n522) );
  BUF_X1 U610 ( .A(n572), .Z(n523) );
  INV_X1 U611 ( .A(n625), .ZN(n526) );
  NOR2_X1 U612 ( .A1(n548), .A2(n542), .ZN(n524) );
  XNOR2_X1 U613 ( .A(KEYINPUT103), .B(n524), .ZN(n635) );
  NAND2_X1 U614 ( .A1(n632), .A2(n635), .ZN(n530) );
  NOR2_X1 U615 ( .A1(KEYINPUT75), .A2(n530), .ZN(n525) );
  NOR2_X1 U616 ( .A1(n526), .A2(n525), .ZN(n528) );
  XOR2_X1 U617 ( .A(KEYINPUT76), .B(n530), .Z(n532) );
  INV_X1 U618 ( .A(n532), .ZN(n585) );
  NAND2_X1 U619 ( .A1(KEYINPUT67), .A2(n585), .ZN(n527) );
  NAND2_X1 U620 ( .A1(n528), .A2(n527), .ZN(n529) );
  INV_X1 U621 ( .A(n530), .ZN(n646) );
  NAND2_X1 U622 ( .A1(KEYINPUT47), .A2(n646), .ZN(n531) );
  NAND2_X1 U623 ( .A1(n531), .A2(KEYINPUT75), .ZN(n546) );
  NOR2_X1 U624 ( .A1(KEYINPUT67), .A2(n532), .ZN(n533) );
  NAND2_X1 U625 ( .A1(n625), .A2(n533), .ZN(n534) );
  NOR2_X1 U626 ( .A1(n534), .A2(KEYINPUT47), .ZN(n544) );
  BUF_X1 U627 ( .A(n535), .Z(n536) );
  INV_X1 U628 ( .A(n536), .ZN(n557) );
  XNOR2_X1 U629 ( .A(n537), .B(KEYINPUT30), .ZN(n541) );
  INV_X1 U630 ( .A(n651), .ZN(n587) );
  NOR2_X1 U631 ( .A1(n594), .A2(n587), .ZN(n656) );
  NAND2_X1 U632 ( .A1(n538), .A2(n656), .ZN(n580) );
  NOR2_X1 U633 ( .A1(n580), .A2(n539), .ZN(n540) );
  INV_X1 U634 ( .A(n542), .ZN(n549) );
  NOR2_X1 U635 ( .A1(n548), .A2(n549), .ZN(n575) );
  NOR2_X1 U636 ( .A1(n557), .A2(n543), .ZN(n630) );
  NOR2_X1 U637 ( .A1(n544), .A2(n630), .ZN(n545) );
  AND2_X1 U638 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U639 ( .A(KEYINPUT38), .B(n557), .ZN(n642) );
  NAND2_X1 U640 ( .A1(n642), .A2(n641), .ZN(n645) );
  NOR2_X1 U641 ( .A1(n645), .A2(n644), .ZN(n550) );
  XNOR2_X1 U642 ( .A(KEYINPUT41), .B(n550), .ZN(n671) );
  NOR2_X1 U643 ( .A1(n671), .A2(n551), .ZN(n552) );
  XNOR2_X1 U644 ( .A(KEYINPUT42), .B(n552), .ZN(n742) );
  INV_X1 U645 ( .A(KEYINPUT40), .ZN(n556) );
  XOR2_X1 U646 ( .A(KEYINPUT79), .B(KEYINPUT39), .Z(n553) );
  NAND2_X1 U647 ( .A1(n565), .A2(n381), .ZN(n555) );
  XNOR2_X1 U648 ( .A(n556), .B(n555), .ZN(n741) );
  NOR2_X1 U649 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U650 ( .A(n560), .B(KEYINPUT107), .ZN(n561) );
  NOR2_X1 U651 ( .A1(n382), .A2(n561), .ZN(n562) );
  XNOR2_X1 U652 ( .A(n562), .B(KEYINPUT43), .ZN(n563) );
  NOR2_X1 U653 ( .A1(n536), .A2(n563), .ZN(n639) );
  NOR2_X1 U654 ( .A1(n564), .A2(n639), .ZN(n566) );
  INV_X1 U655 ( .A(n635), .ZN(n626) );
  NAND2_X1 U656 ( .A1(n565), .A2(n626), .ZN(n638) );
  NAND2_X1 U657 ( .A1(n566), .A2(n638), .ZN(n727) );
  INV_X1 U658 ( .A(G898), .ZN(n567) );
  NAND2_X1 U659 ( .A1(G953), .A2(n567), .ZN(n721) );
  NOR2_X1 U660 ( .A1(n568), .A2(n721), .ZN(n569) );
  NOR2_X1 U661 ( .A1(n570), .A2(n569), .ZN(n571) );
  INV_X1 U662 ( .A(n588), .ZN(n583) );
  NAND2_X1 U663 ( .A1(n656), .A2(n655), .ZN(n582) );
  NOR2_X1 U664 ( .A1(n596), .A2(n582), .ZN(n574) );
  XOR2_X1 U665 ( .A(KEYINPUT73), .B(KEYINPUT78), .Z(n576) );
  XNOR2_X1 U666 ( .A(KEYINPUT35), .B(n576), .ZN(n577) );
  NAND2_X1 U667 ( .A1(n739), .A2(KEYINPUT44), .ZN(n579) );
  NOR2_X1 U668 ( .A1(n583), .A2(n580), .ZN(n581) );
  NAND2_X1 U669 ( .A1(n581), .A2(n654), .ZN(n620) );
  OR2_X1 U670 ( .A1(n654), .A2(n582), .ZN(n661) );
  NOR2_X1 U671 ( .A1(n661), .A2(n583), .ZN(n584) );
  XNOR2_X1 U672 ( .A(n584), .B(KEYINPUT31), .ZN(n634) );
  NAND2_X1 U673 ( .A1(n620), .A2(n634), .ZN(n586) );
  NAND2_X1 U674 ( .A1(n586), .A2(n585), .ZN(n591) );
  INV_X1 U675 ( .A(n594), .ZN(n650) );
  AND2_X1 U676 ( .A1(n596), .A2(n650), .ZN(n590) );
  NAND2_X1 U677 ( .A1(n592), .A2(n590), .ZN(n618) );
  AND2_X1 U678 ( .A1(n382), .A2(n596), .ZN(n597) );
  NOR2_X1 U679 ( .A1(n727), .A2(n677), .ZN(n600) );
  NOR2_X4 U680 ( .A1(n602), .A2(n601), .ZN(n703) );
  NAND2_X1 U681 ( .A1(n703), .A2(G469), .ZN(n606) );
  XOR2_X1 U682 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n603) );
  XNOR2_X1 U683 ( .A(n606), .B(n605), .ZN(n607) );
  INV_X1 U684 ( .A(KEYINPUT119), .ZN(n608) );
  XNOR2_X1 U685 ( .A(n609), .B(n608), .ZN(G54) );
  NAND2_X1 U686 ( .A1(n703), .A2(G472), .ZN(n612) );
  XNOR2_X1 U687 ( .A(n610), .B(n436), .ZN(n611) );
  XNOR2_X1 U688 ( .A(n612), .B(n611), .ZN(n613) );
  XOR2_X1 U689 ( .A(KEYINPUT83), .B(KEYINPUT87), .Z(n614) );
  XNOR2_X1 U690 ( .A(n616), .B(n615), .ZN(G57) );
  XOR2_X1 U691 ( .A(G101), .B(KEYINPUT111), .Z(n617) );
  XNOR2_X1 U692 ( .A(n618), .B(n617), .ZN(G3) );
  NOR2_X1 U693 ( .A1(n632), .A2(n620), .ZN(n619) );
  XOR2_X1 U694 ( .A(G104), .B(n619), .Z(G6) );
  NOR2_X1 U695 ( .A1(n635), .A2(n620), .ZN(n622) );
  XNOR2_X1 U696 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n621) );
  XNOR2_X1 U697 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U698 ( .A(G107), .B(n623), .ZN(G9) );
  XNOR2_X1 U699 ( .A(G110), .B(n624), .ZN(G12) );
  XOR2_X1 U700 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n628) );
  NAND2_X1 U701 ( .A1(n625), .A2(n626), .ZN(n627) );
  XNOR2_X1 U702 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U703 ( .A(G128), .B(n629), .ZN(G30) );
  XOR2_X1 U704 ( .A(G143), .B(n630), .Z(G45) );
  NAND2_X1 U705 ( .A1(n625), .A2(n381), .ZN(n631) );
  XNOR2_X1 U706 ( .A(n631), .B(G146), .ZN(G48) );
  NOR2_X1 U707 ( .A1(n632), .A2(n634), .ZN(n633) );
  XOR2_X1 U708 ( .A(G113), .B(n633), .Z(G15) );
  NOR2_X1 U709 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U710 ( .A(G116), .B(n636), .Z(G18) );
  XOR2_X1 U711 ( .A(G134), .B(KEYINPUT113), .Z(n637) );
  XNOR2_X1 U712 ( .A(n638), .B(n637), .ZN(G36) );
  XOR2_X1 U713 ( .A(G140), .B(n639), .Z(n640) );
  XNOR2_X1 U714 ( .A(KEYINPUT114), .B(n640), .ZN(G42) );
  XOR2_X1 U715 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n690) );
  NOR2_X1 U716 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U717 ( .A1(n644), .A2(n643), .ZN(n648) );
  NOR2_X1 U718 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U719 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U720 ( .A1(n672), .A2(n649), .ZN(n667) );
  NOR2_X1 U721 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U722 ( .A(n652), .B(KEYINPUT49), .ZN(n653) );
  NAND2_X1 U723 ( .A1(n654), .A2(n653), .ZN(n659) );
  NOR2_X1 U724 ( .A1(n656), .A2(n382), .ZN(n657) );
  XNOR2_X1 U725 ( .A(n657), .B(KEYINPUT50), .ZN(n658) );
  NOR2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U727 ( .A(n660), .B(KEYINPUT115), .ZN(n662) );
  NAND2_X1 U728 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U729 ( .A(KEYINPUT51), .B(n663), .ZN(n664) );
  NOR2_X1 U730 ( .A1(n671), .A2(n664), .ZN(n665) );
  XNOR2_X1 U731 ( .A(n665), .B(KEYINPUT116), .ZN(n666) );
  NOR2_X1 U732 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U733 ( .A(n668), .B(KEYINPUT52), .ZN(n669) );
  NOR2_X1 U734 ( .A1(n670), .A2(n669), .ZN(n674) );
  NOR2_X1 U735 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U736 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U737 ( .A(n675), .B(KEYINPUT117), .ZN(n676) );
  NOR2_X1 U738 ( .A1(G953), .A2(n676), .ZN(n688) );
  XOR2_X1 U739 ( .A(KEYINPUT2), .B(KEYINPUT74), .Z(n679) );
  BUF_X1 U740 ( .A(n677), .Z(n678) );
  XOR2_X1 U741 ( .A(KEYINPUT77), .B(n680), .Z(n686) );
  NAND2_X1 U742 ( .A1(n727), .A2(KEYINPUT74), .ZN(n681) );
  XNOR2_X1 U743 ( .A(n681), .B(KEYINPUT2), .ZN(n684) );
  INV_X1 U744 ( .A(n727), .ZN(n682) );
  NAND2_X1 U745 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U746 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U748 ( .A(n690), .B(n689), .ZN(G75) );
  NAND2_X1 U749 ( .A1(n703), .A2(G210), .ZN(n694) );
  XNOR2_X1 U750 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n693) );
  XNOR2_X1 U751 ( .A(n691), .B(KEYINPUT84), .ZN(n692) );
  XNOR2_X1 U752 ( .A(n694), .B(n438), .ZN(n695) );
  XNOR2_X1 U753 ( .A(KEYINPUT56), .B(n696), .ZN(G51) );
  NAND2_X1 U754 ( .A1(n703), .A2(G475), .ZN(n700) );
  XOR2_X1 U755 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n697) );
  XNOR2_X1 U756 ( .A(KEYINPUT60), .B(n702), .ZN(G60) );
  NAND2_X1 U757 ( .A1(G478), .A2(n708), .ZN(n704) );
  XNOR2_X1 U758 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U759 ( .A1(n712), .A2(n706), .ZN(G63) );
  XOR2_X1 U760 ( .A(n707), .B(KEYINPUT121), .Z(n710) );
  NAND2_X1 U761 ( .A1(n708), .A2(G217), .ZN(n709) );
  XNOR2_X1 U762 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U763 ( .A1(n712), .A2(n711), .ZN(G66) );
  XNOR2_X1 U764 ( .A(KEYINPUT123), .B(n713), .ZN(n718) );
  NAND2_X1 U765 ( .A1(G224), .A2(G953), .ZN(n714) );
  XNOR2_X1 U766 ( .A(n714), .B(KEYINPUT61), .ZN(n715) );
  XNOR2_X1 U767 ( .A(KEYINPUT122), .B(n715), .ZN(n716) );
  NAND2_X1 U768 ( .A1(n716), .A2(G898), .ZN(n717) );
  NAND2_X1 U769 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U770 ( .A(n719), .B(KEYINPUT124), .ZN(n723) );
  NAND2_X1 U771 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U772 ( .A(n723), .B(n722), .Z(G69) );
  XOR2_X1 U773 ( .A(n724), .B(KEYINPUT125), .Z(n725) );
  XOR2_X1 U774 ( .A(n726), .B(n725), .Z(n731) );
  XNOR2_X1 U775 ( .A(n727), .B(n731), .ZN(n729) );
  NAND2_X1 U776 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U777 ( .A(n730), .B(KEYINPUT126), .ZN(n736) );
  XNOR2_X1 U778 ( .A(G227), .B(n731), .ZN(n732) );
  NAND2_X1 U779 ( .A1(n732), .A2(G900), .ZN(n733) );
  XOR2_X1 U780 ( .A(KEYINPUT127), .B(n733), .Z(n734) );
  NAND2_X1 U781 ( .A1(G953), .A2(n734), .ZN(n735) );
  NAND2_X1 U782 ( .A1(n736), .A2(n735), .ZN(G72) );
  XNOR2_X1 U783 ( .A(G125), .B(n737), .ZN(n738) );
  XNOR2_X1 U784 ( .A(n738), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U785 ( .A(n739), .B(G122), .Z(G24) );
  XNOR2_X1 U786 ( .A(n740), .B(G119), .ZN(G21) );
  XOR2_X1 U787 ( .A(n741), .B(G131), .Z(G33) );
  XOR2_X1 U788 ( .A(G137), .B(n742), .Z(G39) );
endmodule

