//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1185, new_n1186, new_n1187, new_n1188, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n212), .B(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G87), .A2(G250), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(KEYINPUT66), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT65), .B(G238), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n220), .B1(G68), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G116), .A2(G270), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n219), .A2(KEYINPUT66), .ZN(new_n225));
  AND3_X1   g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G226), .ZN(new_n227));
  INV_X1    g0027(.A(G77), .ZN(new_n228));
  INV_X1    g0028(.A(G244), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n226), .B1(new_n201), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(new_n210), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT1), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n233), .A2(new_n208), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n202), .A2(new_n203), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n235), .A2(G50), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  AOI211_X1 g0037(.A(new_n214), .B(new_n232), .C1(new_n234), .C2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G250), .B(G257), .Z(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G68), .B(G77), .Z(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G58), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n254), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n222), .A2(new_n259), .B1(G107), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n257), .A2(new_n258), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(G232), .A3(new_n254), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G41), .ZN(new_n267));
  OAI211_X1 g0067(.A(G1), .B(G13), .C1(new_n256), .C2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G179), .ZN(new_n271));
  INV_X1    g0071(.A(G45), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT67), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT67), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G45), .ZN(new_n275));
  AOI21_X1  g0075(.A(G41), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n207), .A2(G274), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n268), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G244), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n270), .A2(new_n271), .A3(new_n279), .A4(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT71), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n278), .B1(new_n266), .B2(new_n269), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n287), .A2(KEYINPUT71), .A3(new_n271), .A4(new_n283), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT8), .B(G58), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n290), .A2(new_n292), .B1(new_n208), .B2(new_n228), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n293), .A2(KEYINPUT69), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(KEYINPUT69), .ZN(new_n295));
  XOR2_X1   g0095(.A(KEYINPUT15), .B(G87), .Z(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n208), .A2(G33), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n294), .B(new_n295), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n233), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT70), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(G77), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n207), .A2(G20), .ZN(new_n307));
  INV_X1    g0107(.A(new_n301), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n304), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n302), .B(new_n306), .C1(new_n228), .C2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n287), .A2(new_n283), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n289), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT13), .ZN(new_n315));
  OAI211_X1 g0115(.A(G226), .B(new_n254), .C1(new_n260), .C2(new_n261), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT72), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n264), .A2(KEYINPUT72), .A3(G226), .A4(new_n254), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G33), .A2(G97), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n264), .A2(G232), .A3(G1698), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n318), .A2(new_n319), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n269), .ZN(new_n323));
  INV_X1    g0123(.A(G238), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n281), .A2(new_n324), .B1(new_n276), .B2(new_n277), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n315), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  AOI211_X1 g0127(.A(KEYINPUT13), .B(new_n325), .C1(new_n322), .C2(new_n269), .ZN(new_n328));
  OAI21_X1  g0128(.A(G169), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT14), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n327), .A2(new_n328), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G179), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT14), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n333), .B(G169), .C1(new_n327), .C2(new_n328), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n330), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n298), .A2(new_n228), .B1(new_n208), .B2(G68), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT73), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI221_X1 g0138(.A(KEYINPUT73), .B1(new_n208), .B2(G68), .C1(new_n298), .C2(new_n228), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n338), .B(new_n339), .C1(new_n201), .C2(new_n292), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n301), .ZN(new_n341));
  XOR2_X1   g0141(.A(new_n341), .B(KEYINPUT11), .Z(new_n342));
  INV_X1    g0142(.A(new_n303), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT70), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT70), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n303), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(KEYINPUT12), .A3(new_n203), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n309), .A2(KEYINPUT12), .ZN(new_n349));
  OAI221_X1 g0149(.A(new_n348), .B1(KEYINPUT12), .B2(new_n343), .C1(new_n349), .C2(new_n203), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n342), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n335), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n331), .A2(G190), .ZN(new_n354));
  INV_X1    g0154(.A(G200), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n351), .B(new_n354), .C1(new_n331), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n314), .B1(new_n357), .B2(KEYINPUT74), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G58), .A2(G68), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT76), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(KEYINPUT76), .A2(G58), .A3(G68), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(new_n235), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n208), .A2(new_n256), .A3(G159), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT77), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n291), .A2(KEYINPUT77), .A3(G159), .ZN(new_n368));
  AOI22_X1  g0168(.A1(G20), .A2(new_n364), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n257), .A2(new_n208), .A3(new_n258), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT7), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n258), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT75), .B1(new_n374), .B2(G68), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT75), .ZN(new_n376));
  AOI211_X1 g0176(.A(new_n376), .B(new_n203), .C1(new_n372), .C2(new_n373), .ZN(new_n377));
  OAI211_X1 g0177(.A(KEYINPUT16), .B(new_n369), .C1(new_n375), .C2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT7), .B1(new_n262), .B2(new_n208), .ZN(new_n379));
  INV_X1    g0179(.A(new_n373), .ZN(new_n380));
  OAI21_X1  g0180(.A(G68), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n369), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT16), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n308), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n378), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n290), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n307), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n387), .A2(new_n301), .B1(new_n303), .B2(new_n386), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G223), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n254), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n227), .A2(G1698), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n392), .B(new_n393), .C1(new_n260), .C2(new_n261), .ZN(new_n394));
  NAND2_X1  g0194(.A1(G33), .A2(G87), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT78), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT78), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n394), .A2(new_n398), .A3(new_n395), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n269), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n278), .B1(G232), .B2(new_n282), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G169), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n400), .A2(G179), .A3(new_n401), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT18), .B1(new_n390), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n388), .B1(new_n378), .B2(new_n384), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n400), .A2(G179), .A3(new_n401), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n312), .B1(new_n400), .B2(new_n401), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT18), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n407), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT79), .B1(new_n406), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n400), .A2(G190), .A3(new_n401), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n402), .A2(G200), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n385), .A2(new_n414), .A3(new_n389), .A4(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT17), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n407), .A2(KEYINPUT17), .A3(new_n414), .A4(new_n415), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n203), .B1(new_n372), .B2(new_n373), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n364), .A2(G20), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n367), .A2(new_n368), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n383), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n301), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n381), .A2(new_n376), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n421), .A2(KEYINPUT75), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n424), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n426), .B1(new_n429), .B2(KEYINPUT16), .ZN(new_n430));
  OAI211_X1 g0230(.A(KEYINPUT18), .B(new_n405), .C1(new_n430), .C2(new_n388), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n411), .B1(new_n407), .B2(new_n410), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT79), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n413), .A2(new_n420), .A3(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n309), .A2(new_n228), .ZN(new_n436));
  AOI211_X1 g0236(.A(new_n305), .B(new_n436), .C1(new_n299), .C2(new_n301), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n311), .A2(G200), .ZN(new_n438));
  INV_X1    g0238(.A(G190), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n437), .B(new_n438), .C1(new_n439), .C2(new_n311), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n435), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n254), .A2(G222), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n264), .B(new_n443), .C1(new_n391), .C2(new_n254), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n444), .B(new_n269), .C1(G77), .C2(new_n264), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n445), .B(new_n279), .C1(new_n227), .C2(new_n281), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n312), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n308), .A2(G50), .A3(new_n307), .ZN(new_n448));
  INV_X1    g0248(.A(G150), .ZN(new_n449));
  OAI22_X1  g0249(.A1(new_n290), .A2(new_n298), .B1(new_n449), .B2(new_n292), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n450), .B1(G20), .B2(new_n204), .ZN(new_n451));
  OAI221_X1 g0251(.A(new_n448), .B1(G50), .B2(new_n303), .C1(new_n451), .C2(new_n308), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n447), .B(new_n452), .C1(G179), .C2(new_n446), .ZN(new_n453));
  XOR2_X1   g0253(.A(new_n453), .B(KEYINPUT68), .Z(new_n454));
  AOI21_X1  g0254(.A(new_n454), .B1(new_n357), .B2(KEYINPUT74), .ZN(new_n455));
  XNOR2_X1  g0255(.A(new_n452), .B(KEYINPUT9), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n446), .A2(G200), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n456), .B(new_n457), .C1(new_n439), .C2(new_n446), .ZN(new_n458));
  XNOR2_X1  g0258(.A(new_n458), .B(KEYINPUT10), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n359), .A2(new_n442), .A3(new_n455), .A4(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(G250), .B(new_n254), .C1(new_n260), .C2(new_n261), .ZN(new_n461));
  OAI211_X1 g0261(.A(G257), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G294), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n269), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT84), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n272), .A2(G1), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n267), .A2(KEYINPUT5), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT5), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G41), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n468), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G274), .ZN(new_n473));
  OR2_X1    g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(G264), .A3(new_n268), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n464), .A2(KEYINPUT84), .A3(new_n269), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n467), .A2(new_n474), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G169), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n465), .A2(new_n475), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(G179), .A3(new_n474), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n256), .A2(G20), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G116), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n208), .A2(G107), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n484), .B(KEYINPUT23), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n208), .B(G87), .C1(new_n260), .C2(new_n261), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n486), .A2(KEYINPUT22), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n486), .A2(KEYINPUT22), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n483), .B(new_n485), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT24), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n486), .B(KEYINPUT22), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n492), .A2(KEYINPUT24), .A3(new_n483), .A4(new_n485), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(new_n301), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n207), .A2(G33), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n308), .A2(new_n303), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G107), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n303), .A2(G107), .ZN(new_n499));
  XNOR2_X1  g0299(.A(new_n499), .B(KEYINPUT25), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n494), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n481), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n465), .A2(new_n475), .A3(new_n474), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n355), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(new_n477), .B2(G190), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n505), .A2(new_n498), .A3(new_n500), .A4(new_n494), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n304), .A2(new_n296), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT19), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n482), .A2(new_n509), .A3(G97), .ZN(new_n510));
  NOR2_X1   g0310(.A1(G97), .A2(G107), .ZN(new_n511));
  INV_X1    g0311(.A(G87), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n511), .A2(new_n512), .B1(new_n320), .B2(new_n208), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n510), .B1(new_n513), .B2(new_n509), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n208), .B(G68), .C1(new_n260), .C2(new_n261), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT83), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n264), .A2(KEYINPUT83), .A3(new_n208), .A4(G68), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n514), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n508), .B1(new_n519), .B2(new_n301), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n497), .A2(new_n296), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n324), .A2(new_n254), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n229), .A2(G1698), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n522), .B(new_n523), .C1(new_n260), .C2(new_n261), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G116), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n268), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n207), .A2(G45), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n527), .A2(new_n473), .ZN(new_n528));
  AND2_X1   g0328(.A1(G33), .A2(G41), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n527), .B(G250), .C1(new_n529), .C2(new_n233), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n526), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n520), .A2(new_n521), .B1(new_n271), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n528), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n524), .A2(new_n525), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n534), .B(new_n530), .C1(new_n535), .C2(new_n268), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n312), .ZN(new_n537));
  NOR4_X1   g0337(.A1(new_n526), .A2(new_n439), .A3(new_n531), .A4(new_n528), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(G200), .B2(new_n536), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n496), .A2(new_n512), .ZN(new_n540));
  AOI211_X1 g0340(.A(new_n540), .B(new_n508), .C1(new_n301), .C2(new_n519), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n533), .A2(new_n537), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n259), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n543));
  OAI211_X1 g0343(.A(G244), .B(new_n254), .C1(new_n260), .C2(new_n261), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT82), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT4), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n546), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n545), .A2(new_n546), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n264), .A2(G244), .A3(new_n254), .A4(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n543), .A2(new_n547), .A3(new_n548), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n269), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n472), .A2(new_n268), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n474), .B1(new_n218), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n312), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n374), .A2(G107), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT6), .ZN(new_n559));
  INV_X1    g0359(.A(G107), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n217), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n559), .B1(new_n561), .B2(new_n511), .ZN(new_n562));
  NAND2_X1  g0362(.A1(KEYINPUT6), .A2(G97), .ZN(new_n563));
  OAI21_X1  g0363(.A(KEYINPUT81), .B1(new_n563), .B2(G107), .ZN(new_n564));
  OR3_X1    g0364(.A1(new_n563), .A2(KEYINPUT81), .A3(G107), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n562), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G20), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n291), .A2(G77), .ZN(new_n568));
  XNOR2_X1  g0368(.A(new_n568), .B(KEYINPUT80), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n558), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n301), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n303), .A2(G97), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n496), .B2(new_n217), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n554), .B1(new_n551), .B2(new_n269), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n271), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n557), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(G190), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n574), .B1(new_n570), .B2(new_n301), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n580), .B(new_n581), .C1(new_n355), .C2(new_n577), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n542), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n304), .A2(G116), .A3(new_n308), .A4(new_n495), .ZN(new_n584));
  NAND2_X1  g0384(.A1(G33), .A2(G283), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n585), .B(new_n208), .C1(G33), .C2(new_n217), .ZN(new_n586));
  INV_X1    g0386(.A(G116), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G20), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n301), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT20), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n586), .A2(KEYINPUT20), .A3(new_n301), .A4(new_n588), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n347), .A2(new_n587), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n584), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n472), .A2(G270), .A3(new_n268), .ZN(new_n596));
  OAI211_X1 g0396(.A(G264), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n597));
  OAI211_X1 g0397(.A(G257), .B(new_n254), .C1(new_n260), .C2(new_n261), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n257), .A2(G303), .A3(new_n258), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n474), .B(new_n596), .C1(new_n600), .C2(new_n268), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n595), .A2(G169), .A3(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT21), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n601), .A2(new_n271), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n595), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n595), .A2(KEYINPUT21), .A3(new_n601), .A4(G169), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n604), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n595), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n601), .A2(new_n439), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(G200), .B2(new_n601), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n608), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n507), .A2(new_n583), .A3(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n460), .A2(new_n613), .ZN(G372));
  NAND2_X1  g0414(.A1(new_n353), .A2(new_n314), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n615), .A2(new_n356), .A3(new_n420), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n431), .A2(new_n432), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n454), .B1(new_n619), .B2(new_n459), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n533), .A2(new_n537), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n506), .A2(new_n579), .A3(new_n542), .A4(new_n582), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n608), .B1(new_n481), .B2(new_n501), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n539), .A2(new_n541), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n626), .A2(new_n579), .A3(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n557), .A2(new_n576), .A3(new_n578), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT26), .B1(new_n629), .B2(new_n542), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n624), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n620), .B1(new_n460), .B2(new_n632), .ZN(G369));
  INV_X1    g0433(.A(G13), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(G20), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n207), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(G213), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(G343), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n501), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n507), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n641), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n643), .B1(new_n502), .B2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n608), .A2(new_n644), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(G330), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n612), .B1(new_n609), .B2(new_n644), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n608), .A2(new_n595), .A3(new_n641), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n481), .A2(new_n501), .A3(new_n644), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n507), .A2(new_n646), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(G399));
  INV_X1    g0455(.A(new_n211), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(G41), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NOR4_X1   g0458(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(G1), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n236), .B2(new_n658), .ZN(new_n661));
  XOR2_X1   g0461(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n662));
  XNOR2_X1  g0462(.A(new_n661), .B(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n644), .B1(new_n624), .B2(new_n631), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT29), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n601), .A2(new_n271), .A3(new_n536), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT86), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n601), .A2(new_n536), .A3(KEYINPUT86), .A4(new_n271), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n669), .A2(new_n556), .A3(new_n503), .A4(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT30), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n552), .A2(new_n479), .A3(new_n555), .A4(new_n532), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n601), .A2(new_n271), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n479), .A2(new_n532), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n676), .A2(KEYINPUT30), .A3(new_n605), .A4(new_n577), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n671), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n678), .A2(KEYINPUT31), .A3(new_n641), .ZN(new_n679));
  AOI21_X1  g0479(.A(KEYINPUT31), .B1(new_n678), .B2(new_n641), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n507), .A2(new_n583), .A3(new_n612), .A4(new_n644), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n648), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n666), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n663), .B1(new_n685), .B2(G1), .ZN(G364));
  XNOR2_X1  g0486(.A(new_n651), .B(KEYINPUT87), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n635), .A2(G45), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT88), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT88), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G1), .A3(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n657), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n649), .A2(new_n650), .ZN(new_n694));
  OAI211_X1 g0494(.A(new_n687), .B(new_n693), .C1(G330), .C2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n208), .A2(new_n439), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n271), .A2(new_n355), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n271), .A2(G200), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n208), .A2(G190), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI22_X1  g0501(.A1(new_n698), .A2(new_n201), .B1(new_n701), .B2(new_n228), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n696), .A2(new_n699), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n702), .B1(G58), .B2(new_n704), .ZN(new_n705));
  XOR2_X1   g0505(.A(new_n705), .B(KEYINPUT89), .Z(new_n706));
  NOR2_X1   g0506(.A1(new_n355), .A2(G179), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n696), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(new_n512), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n707), .A2(new_n700), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT90), .Z(new_n712));
  NAND2_X1  g0512(.A1(new_n697), .A2(new_n700), .ZN(new_n713));
  OAI22_X1  g0513(.A1(new_n712), .A2(new_n560), .B1(new_n203), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(G179), .A2(G200), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n700), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(G159), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n262), .B1(new_n719), .B2(KEYINPUT32), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n715), .A2(G190), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G20), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n720), .B1(new_n217), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n714), .A2(new_n724), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n710), .B(new_n725), .C1(KEYINPUT32), .C2(new_n719), .ZN(new_n726));
  INV_X1    g0526(.A(G322), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n703), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(G326), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n262), .B1(new_n698), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(G303), .ZN(new_n731));
  INV_X1    g0531(.A(G329), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n708), .A2(new_n731), .B1(new_n716), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n701), .ZN(new_n734));
  AOI211_X1 g0534(.A(new_n730), .B(new_n733), .C1(G311), .C2(new_n734), .ZN(new_n735));
  XNOR2_X1  g0535(.A(KEYINPUT91), .B(KEYINPUT33), .ZN(new_n736));
  INV_X1    g0536(.A(G317), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n736), .B(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n713), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n738), .A2(new_n739), .B1(G294), .B2(new_n722), .ZN(new_n740));
  INV_X1    g0540(.A(G283), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n735), .B(new_n740), .C1(new_n741), .C2(new_n712), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n726), .B1(new_n728), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n233), .B1(G20), .B2(new_n312), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n656), .A2(new_n264), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n273), .A2(new_n275), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n747), .B1(new_n237), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n749), .B1(new_n272), .B2(new_n252), .ZN(new_n750));
  INV_X1    g0550(.A(G355), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n211), .A2(new_n264), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n750), .B1(G116), .B2(new_n211), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n744), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n756), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n745), .B(new_n758), .C1(new_n694), .C2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n695), .B1(new_n693), .B2(new_n760), .ZN(G396));
  AND4_X1   g0561(.A1(new_n310), .A2(new_n289), .A3(new_n313), .A4(new_n644), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT93), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n310), .A2(new_n763), .A3(new_n641), .ZN(new_n764));
  OAI21_X1  g0564(.A(KEYINPUT93), .B1(new_n437), .B2(new_n644), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n440), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n762), .B1(new_n766), .B2(new_n314), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n754), .ZN(new_n769));
  INV_X1    g0569(.A(new_n712), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n264), .B1(new_n770), .B2(G87), .ZN(new_n771));
  INV_X1    g0571(.A(new_n698), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G303), .ZN(new_n773));
  INV_X1    g0573(.A(new_n716), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n774), .A2(G311), .B1(new_n722), .B2(G97), .ZN(new_n775));
  INV_X1    g0575(.A(G294), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n560), .A2(new_n708), .B1(new_n703), .B2(new_n776), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n713), .A2(new_n741), .B1(new_n701), .B2(new_n587), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n771), .A2(new_n773), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n774), .A2(G132), .ZN(new_n781));
  AOI22_X1  g0581(.A1(G143), .A2(new_n704), .B1(new_n739), .B2(G150), .ZN(new_n782));
  INV_X1    g0582(.A(G137), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n782), .B1(new_n783), .B2(new_n698), .C1(new_n717), .C2(new_n701), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT34), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n262), .B(new_n781), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n722), .A2(G58), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n784), .A2(new_n785), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n712), .A2(new_n203), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n786), .A2(new_n787), .A3(new_n788), .A4(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n708), .A2(new_n201), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n780), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n744), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n744), .A2(new_n754), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT92), .Z(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n228), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n769), .A2(new_n692), .A3(new_n794), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n664), .A2(new_n768), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n767), .B(new_n644), .C1(new_n624), .C2(new_n631), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(new_n684), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n798), .B1(new_n802), .B2(new_n692), .ZN(G384));
  NOR2_X1   g0603(.A1(new_n353), .A2(new_n641), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT38), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n403), .A2(new_n404), .A3(new_n639), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n390), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT37), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n808), .A2(new_n809), .A3(new_n416), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n369), .B1(new_n375), .B2(new_n377), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n383), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n812), .A2(new_n301), .A3(new_n378), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n813), .A2(new_n389), .B1(new_n410), .B2(new_n639), .ZN(new_n814));
  INV_X1    g0614(.A(new_n416), .ZN(new_n815));
  OAI21_X1  g0615(.A(KEYINPUT37), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n639), .B1(new_n813), .B2(new_n389), .ZN(new_n817));
  AOI221_X4 g0617(.A(new_n806), .B1(new_n810), .B2(new_n816), .C1(new_n435), .C2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n435), .A2(new_n817), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n816), .A2(new_n810), .ZN(new_n820));
  AOI21_X1  g0620(.A(KEYINPUT38), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(KEYINPUT39), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n639), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n418), .A2(new_n419), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n390), .B(new_n823), .C1(new_n617), .C2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT94), .ZN(new_n826));
  AND3_X1   g0626(.A1(new_n808), .A2(new_n809), .A3(new_n416), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n809), .B1(new_n808), .B2(new_n416), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n808), .A2(new_n416), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT37), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n831), .A2(KEYINPUT94), .A3(new_n810), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n825), .A2(new_n829), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n806), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT39), .ZN(new_n835));
  AND3_X1   g0635(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n433), .B1(new_n431), .B2(new_n432), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n836), .A2(new_n837), .A3(new_n824), .ZN(new_n838));
  INV_X1    g0638(.A(new_n817), .ZN(new_n839));
  OAI211_X1 g0639(.A(KEYINPUT38), .B(new_n820), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n834), .A2(new_n835), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n805), .B1(new_n822), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n818), .A2(new_n821), .ZN(new_n843));
  INV_X1    g0643(.A(new_n762), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n800), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n352), .A2(new_n641), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n353), .A2(new_n846), .A3(new_n356), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n335), .A2(new_n352), .A3(new_n641), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n843), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n618), .A2(new_n823), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n842), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n620), .B1(new_n666), .B2(new_n460), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n853), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g0655(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n834), .A2(new_n840), .ZN(new_n858));
  INV_X1    g0658(.A(new_n680), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n678), .A2(KEYINPUT31), .A3(new_n641), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n682), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n861), .A2(new_n849), .A3(new_n767), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n858), .A2(KEYINPUT40), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n820), .B1(new_n838), .B2(new_n839), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n806), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n862), .B1(new_n866), .B2(new_n840), .ZN(new_n867));
  XNOR2_X1  g0667(.A(KEYINPUT97), .B(KEYINPUT40), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n864), .B(G330), .C1(new_n867), .C2(new_n869), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n358), .A2(new_n441), .A3(new_n435), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n871), .A2(new_n455), .A3(new_n459), .A4(new_n683), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n863), .B1(new_n818), .B2(new_n821), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT40), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n834), .B2(new_n840), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n874), .A2(new_n868), .B1(new_n876), .B2(new_n863), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n861), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n873), .B1(new_n878), .B2(new_n460), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n857), .B(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n207), .B2(new_n635), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n587), .B1(new_n566), .B2(KEYINPUT35), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n882), .B(new_n234), .C1(KEYINPUT35), .C2(new_n566), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT36), .ZN(new_n884));
  AND4_X1   g0684(.A1(G77), .A2(new_n237), .A3(new_n362), .A4(new_n363), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n203), .A2(G50), .ZN(new_n886));
  OAI211_X1 g0686(.A(G1), .B(new_n634), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n881), .A2(new_n884), .A3(new_n887), .ZN(G367));
  OAI211_X1 g0688(.A(new_n579), .B(new_n582), .C1(new_n581), .C2(new_n644), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n629), .A2(new_n641), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n891), .A2(new_n654), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n892), .B(KEYINPUT42), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n579), .B1(new_n889), .B2(new_n502), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n644), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n896), .A2(KEYINPUT98), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(KEYINPUT98), .ZN(new_n898));
  OR3_X1    g0698(.A1(new_n621), .A2(new_n541), .A3(new_n644), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n542), .B1(new_n541), .B2(new_n644), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n901), .A2(KEYINPUT43), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n897), .A2(new_n898), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(KEYINPUT43), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n897), .B2(new_n898), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n652), .A2(new_n891), .ZN(new_n907));
  OR3_X1    g0707(.A1(new_n903), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n907), .B1(new_n903), .B2(new_n906), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n691), .B(KEYINPUT99), .Z(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n652), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n647), .A2(new_n654), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n913), .B1(new_n687), .B2(new_n914), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n915), .A2(new_n685), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n654), .A2(new_n653), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n891), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT44), .Z(new_n919));
  NOR2_X1   g0719(.A1(new_n917), .A2(new_n891), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT45), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n916), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n685), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n657), .B(KEYINPUT41), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n912), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n901), .A2(new_n759), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n701), .A2(new_n741), .B1(new_n716), .B2(new_n737), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n264), .B(new_n928), .C1(G294), .C2(new_n739), .ZN(new_n929));
  INV_X1    g0729(.A(new_n708), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT46), .B1(new_n930), .B2(G116), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n703), .A2(new_n731), .ZN(new_n932));
  INV_X1    g0732(.A(G311), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n698), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n711), .A2(new_n217), .ZN(new_n935));
  NOR4_X1   g0735(.A1(new_n931), .A2(new_n932), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n722), .A2(G107), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n930), .A2(KEYINPUT46), .A3(G116), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n929), .A2(new_n936), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(G143), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n698), .A2(new_n940), .B1(new_n703), .B2(new_n449), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(G68), .B2(new_n722), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n202), .B2(new_n708), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n264), .B1(new_n716), .B2(new_n783), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n713), .A2(new_n717), .B1(new_n711), .B2(new_n228), .ZN(new_n945));
  OR3_X1    g0745(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n701), .A2(new_n201), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n939), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT47), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n744), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n757), .B1(new_n211), .B2(new_n297), .C1(new_n747), .C2(new_n245), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n950), .A2(new_n692), .A3(new_n951), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n910), .A2(new_n926), .B1(new_n927), .B2(new_n952), .ZN(G387));
  NAND2_X1  g0753(.A1(new_n915), .A2(new_n912), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n704), .A2(G50), .B1(new_n722), .B2(new_n296), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n264), .B1(new_n955), .B2(KEYINPUT102), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(KEYINPUT102), .B2(new_n955), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n930), .A2(G77), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n449), .B2(new_n716), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n770), .A2(G97), .B1(KEYINPUT101), .B2(new_n959), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n957), .B(new_n960), .C1(KEYINPUT101), .C2(new_n959), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(G159), .B2(new_n772), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n962), .B1(new_n203), .B2(new_n701), .C1(new_n290), .C2(new_n713), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n703), .A2(new_n737), .B1(new_n701), .B2(new_n731), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT103), .Z(new_n965));
  OAI221_X1 g0765(.A(new_n965), .B1(new_n933), .B2(new_n713), .C1(new_n727), .C2(new_n698), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT48), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n967), .B1(new_n741), .B2(new_n723), .C1(new_n776), .C2(new_n708), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT49), .Z(new_n969));
  OAI221_X1 g0769(.A(new_n262), .B1(new_n716), .B2(new_n729), .C1(new_n587), .C2(new_n711), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n963), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n744), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n645), .A2(new_n759), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n659), .B(new_n272), .C1(new_n203), .C2(new_n228), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT100), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n386), .A2(new_n201), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT50), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n746), .B1(new_n975), .B2(new_n977), .C1(new_n242), .C2(new_n748), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(G107), .B2(new_n211), .C1(new_n659), .C2(new_n752), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n757), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n972), .A2(new_n692), .A3(new_n973), .A4(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n657), .B1(new_n915), .B2(new_n685), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n954), .B(new_n981), .C1(new_n916), .C2(new_n982), .ZN(G393));
  NOR2_X1   g0783(.A1(new_n716), .A2(new_n727), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n262), .B1(new_n708), .B2(new_n741), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n698), .A2(new_n737), .B1(new_n703), .B2(new_n933), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT104), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT52), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n713), .A2(new_n731), .B1(new_n701), .B2(new_n776), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(new_n770), .B2(G107), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n989), .B(new_n991), .C1(new_n988), .C2(new_n987), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n984), .B(new_n992), .C1(G116), .C2(new_n722), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n770), .A2(G87), .B1(G50), .B2(new_n739), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n994), .B(new_n264), .C1(new_n203), .C2(new_n708), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n723), .A2(new_n228), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n698), .A2(new_n449), .B1(new_n703), .B2(new_n717), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT51), .Z(new_n998));
  OAI22_X1  g0798(.A1(new_n701), .A2(new_n290), .B1(new_n716), .B2(new_n940), .ZN(new_n999));
  NOR4_X1   g0799(.A1(new_n995), .A2(new_n996), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n993), .A2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT105), .Z(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n744), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n757), .B1(new_n217), .B2(new_n211), .C1(new_n747), .C2(new_n249), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1003), .A2(new_n692), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n756), .B2(new_n891), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n922), .A2(new_n913), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n919), .A2(new_n652), .A3(new_n921), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n915), .A2(new_n685), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n658), .B1(new_n1012), .B2(KEYINPUT106), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n923), .A2(KEYINPUT106), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n1011), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1006), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1007), .A2(new_n912), .A3(new_n1008), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(G390));
  NAND4_X1  g0818(.A1(new_n861), .A2(new_n849), .A3(G330), .A4(new_n767), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n804), .B1(new_n845), .B2(new_n849), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n822), .B2(new_n841), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n850), .A2(new_n805), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1023), .A2(new_n858), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1020), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n835), .B1(new_n866), .B2(new_n840), .ZN(new_n1026));
  AND3_X1   g0826(.A1(new_n834), .A2(new_n835), .A3(new_n840), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1023), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1021), .A2(new_n840), .A3(new_n834), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT107), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1019), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n683), .A2(KEYINPUT107), .A3(new_n767), .A4(new_n849), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1028), .A2(new_n1029), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1025), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n912), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n822), .A2(new_n754), .A3(new_n841), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n262), .B1(new_n701), .B2(new_n217), .C1(new_n560), .C2(new_n713), .ZN(new_n1038));
  OR3_X1    g0838(.A1(new_n789), .A2(new_n709), .A3(new_n996), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(G294), .C2(new_n774), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n587), .B2(new_n703), .C1(new_n741), .C2(new_n698), .ZN(new_n1041));
  XOR2_X1   g0841(.A(KEYINPUT54), .B(G143), .Z(new_n1042));
  AOI22_X1  g0842(.A1(G132), .A2(new_n704), .B1(new_n734), .B2(new_n1042), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n201), .B2(new_n711), .C1(new_n783), .C2(new_n713), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n262), .B(new_n1044), .C1(G125), .C2(new_n774), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n772), .A2(G128), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(new_n717), .C2(new_n723), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n708), .A2(new_n449), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT111), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT53), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1041), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT112), .Z(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n744), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n796), .A2(new_n290), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1037), .A2(new_n1053), .A3(new_n692), .A4(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1036), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n861), .A2(G330), .A3(new_n767), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n849), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1031), .A2(new_n1032), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n845), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n849), .B1(KEYINPUT108), .B2(new_n767), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1062), .A2(new_n1057), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n845), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1062), .A2(new_n1057), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1061), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n872), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n854), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n1025), .B2(new_n1034), .ZN(new_n1071));
  OAI21_X1  g0871(.A(KEYINPUT109), .B1(new_n1071), .B2(new_n658), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1070), .A2(new_n1025), .A3(new_n1034), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n872), .B(new_n620), .C1(new_n460), .C2(new_n666), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n1061), .B2(new_n1066), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1035), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT109), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1076), .A2(new_n1077), .A3(new_n657), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1072), .A2(new_n1073), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT110), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1072), .A2(KEYINPUT110), .A3(new_n1078), .A4(new_n1073), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1056), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(G378));
  INV_X1    g0884(.A(KEYINPUT57), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1069), .A2(KEYINPUT117), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT117), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1074), .A2(new_n1087), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1086), .B(new_n1088), .C1(new_n1035), .C2(new_n1075), .ZN(new_n1089));
  XOR2_X1   g0889(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n452), .A2(new_n823), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(KEYINPUT115), .B(KEYINPUT116), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1092), .B(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n459), .A2(new_n453), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1095), .B1(new_n459), .B2(new_n453), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1091), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1098), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1100), .A2(new_n1090), .A3(new_n1096), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n877), .A2(G330), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1102), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n870), .A2(new_n1104), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n853), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n842), .A2(new_n852), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n851), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1105), .A2(new_n1103), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1085), .B1(new_n1089), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1086), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1088), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1076), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1105), .A2(new_n1103), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n853), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n853), .A2(new_n1105), .A3(new_n1103), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1114), .A2(KEYINPUT57), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1111), .A2(new_n657), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n912), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n693), .B1(new_n1104), .B2(new_n754), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n201), .B1(new_n260), .B2(G41), .ZN(new_n1124));
  INV_X1    g0924(.A(G125), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n723), .A2(new_n449), .B1(new_n698), .B2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(G128), .A2(new_n704), .B1(new_n739), .B2(G132), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n783), .B2(new_n701), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1126), .B(new_n1128), .C1(new_n930), .C2(new_n1042), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT59), .ZN(new_n1130));
  AOI21_X1  g0930(.A(G33), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(G41), .B1(new_n774), .B2(G124), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1131), .B(new_n1132), .C1(new_n717), .C2(new_n711), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1124), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n703), .A2(new_n560), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT114), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n264), .A2(G41), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n739), .A2(G97), .B1(new_n774), .B2(G283), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1137), .A2(new_n958), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n711), .A2(new_n202), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT113), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1142), .B1(new_n587), .B2(new_n698), .C1(new_n297), .C2(new_n701), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n1140), .B(new_n1143), .C1(G68), .C2(new_n722), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT58), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n744), .B1(new_n1135), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n796), .A2(new_n201), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1123), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1122), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1121), .A2(new_n1149), .ZN(G375));
  NAND2_X1  g0950(.A1(new_n1058), .A2(new_n754), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(G97), .A2(new_n930), .B1(new_n774), .B2(G303), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n776), .B2(new_n698), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n262), .B1(new_n712), .B2(new_n228), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT118), .Z(new_n1155));
  AOI22_X1  g0955(.A1(new_n704), .A2(G283), .B1(new_n722), .B2(new_n296), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1155), .B(new_n1156), .C1(new_n560), .C2(new_n701), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1153), .B(new_n1157), .C1(G116), .C2(new_n739), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(G159), .A2(new_n930), .B1(new_n774), .B2(G128), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1159), .B(KEYINPUT119), .Z(new_n1160));
  AOI22_X1  g0960(.A1(new_n739), .A2(new_n1042), .B1(new_n734), .B2(G150), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n772), .A2(G132), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1142), .B1(new_n201), .B2(new_n723), .C1(new_n783), .C2(new_n703), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n1163), .A2(new_n262), .A3(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n744), .B1(new_n1158), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n796), .A2(new_n203), .ZN(new_n1167));
  AND4_X1   g0967(.A1(new_n692), .A2(new_n1151), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n1067), .B2(new_n912), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1074), .A2(new_n1061), .A3(new_n1066), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n925), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1169), .B1(new_n1171), .B2(new_n1075), .ZN(G381));
  XNOR2_X1  g0972(.A(G375), .B(KEYINPUT120), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1056), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1079), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n952), .A2(new_n927), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n908), .A2(new_n909), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n924), .A2(new_n925), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n911), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1177), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1181), .A2(new_n1017), .A3(new_n1016), .ZN(new_n1182));
  OR3_X1    g0982(.A1(new_n1182), .A2(G396), .A3(G393), .ZN(new_n1183));
  OR4_X1    g0983(.A1(G384), .A2(new_n1176), .A3(G381), .A4(new_n1183), .ZN(G407));
  NAND2_X1  g0984(.A1(new_n640), .A2(G213), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1176), .A2(new_n1185), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1186), .A2(KEYINPUT121), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(KEYINPUT121), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1187), .A2(G213), .A3(G407), .A4(new_n1188), .ZN(G409));
  NAND2_X1  g0989(.A1(G390), .A2(G387), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(G393), .B(G396), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1182), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1191), .B1(new_n1182), .B2(new_n1190), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT122), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1119), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1117), .A2(KEYINPUT122), .A3(new_n1118), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(new_n912), .A3(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1114), .A2(new_n925), .A3(new_n1119), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1198), .A2(new_n1148), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n1175), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n1083), .B2(G375), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(KEYINPUT123), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT60), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1170), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1170), .A2(new_n1204), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1205), .A2(new_n657), .A3(new_n1070), .A4(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n1169), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(G384), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT123), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1201), .B(new_n1210), .C1(new_n1083), .C2(G375), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1203), .A2(new_n1185), .A3(new_n1209), .A4(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1212), .A2(KEYINPUT62), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1202), .A2(new_n1185), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1209), .ZN(new_n1215));
  OAI21_X1  g1015(.A(KEYINPUT62), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n640), .A2(G213), .A3(G2897), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1209), .B(new_n1217), .Z(new_n1218));
  AOI21_X1  g1018(.A(KEYINPUT61), .B1(new_n1214), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1216), .A2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1194), .B1(new_n1213), .B2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1203), .A2(new_n1185), .A3(new_n1211), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(KEYINPUT124), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT124), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1203), .A2(new_n1224), .A3(new_n1185), .A4(new_n1211), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1223), .A2(new_n1218), .A3(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT125), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1202), .A2(KEYINPUT63), .A3(new_n1185), .A4(new_n1209), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1192), .A2(new_n1193), .A3(KEYINPUT61), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT63), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1230), .B1(new_n1231), .B2(new_n1212), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1226), .A2(new_n1227), .A3(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1227), .B1(new_n1226), .B2(new_n1232), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1221), .B1(new_n1233), .B2(new_n1234), .ZN(G405));
  XOR2_X1   g1035(.A(new_n1194), .B(KEYINPUT127), .Z(new_n1236));
  NOR2_X1   g1036(.A1(new_n1194), .A2(KEYINPUT127), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(G375), .A2(new_n1175), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1083), .A2(G375), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1215), .A2(KEYINPUT126), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1241), .B(new_n1242), .ZN(new_n1243));
  MUX2_X1   g1043(.A(new_n1236), .B(new_n1237), .S(new_n1243), .Z(G402));
endmodule


