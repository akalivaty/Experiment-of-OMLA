

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593;

  NOR2_X2 U327 ( .A1(n515), .A2(n483), .ZN(n484) );
  XNOR2_X1 U328 ( .A(n369), .B(n582), .ZN(n560) );
  XNOR2_X1 U329 ( .A(n295), .B(n296), .ZN(n357) );
  XNOR2_X1 U330 ( .A(n356), .B(n355), .ZN(n433) );
  NOR2_X1 U331 ( .A1(n483), .A2(n460), .ZN(n554) );
  NOR2_X2 U332 ( .A1(n542), .A2(n454), .ZN(n551) );
  NOR2_X1 U333 ( .A1(n474), .A2(n473), .ZN(n505) );
  XNOR2_X1 U334 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U335 ( .A(n368), .B(n367), .Z(n582) );
  XOR2_X1 U336 ( .A(G78GAT), .B(G148GAT), .Z(n295) );
  NOR2_X1 U337 ( .A1(n582), .A2(n397), .ZN(n398) );
  INV_X1 U338 ( .A(KEYINPUT11), .ZN(n380) );
  XNOR2_X1 U339 ( .A(n381), .B(n380), .ZN(n386) );
  XNOR2_X1 U340 ( .A(n446), .B(n445), .ZN(n447) );
  INV_X1 U341 ( .A(KEYINPUT80), .ZN(n421) );
  XNOR2_X1 U342 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U343 ( .A(n448), .B(n447), .ZN(n450) );
  NOR2_X1 U344 ( .A1(n532), .A2(n496), .ZN(n478) );
  XNOR2_X1 U345 ( .A(n424), .B(n423), .ZN(n439) );
  XOR2_X1 U346 ( .A(n390), .B(n389), .Z(n565) );
  INV_X1 U347 ( .A(G78GAT), .ZN(n479) );
  XNOR2_X1 U348 ( .A(n452), .B(n451), .ZN(n540) );
  XNOR2_X1 U349 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n489) );
  XNOR2_X1 U350 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U351 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U352 ( .A(n490), .B(n489), .ZN(G1351GAT) );
  XNOR2_X1 U353 ( .A(n482), .B(n481), .ZN(G1335GAT) );
  XNOR2_X1 U354 ( .A(G106GAT), .B(KEYINPUT76), .ZN(n296) );
  XOR2_X1 U355 ( .A(G204GAT), .B(n357), .Z(n298) );
  NAND2_X1 U356 ( .A1(G228GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U357 ( .A(n298), .B(n297), .ZN(n315) );
  XOR2_X1 U358 ( .A(KEYINPUT86), .B(KEYINPUT82), .Z(n300) );
  XNOR2_X1 U359 ( .A(G50GAT), .B(KEYINPUT24), .ZN(n299) );
  XNOR2_X1 U360 ( .A(n300), .B(n299), .ZN(n303) );
  XOR2_X1 U361 ( .A(KEYINPUT83), .B(KEYINPUT21), .Z(n302) );
  XNOR2_X1 U362 ( .A(G197GAT), .B(G218GAT), .ZN(n301) );
  XNOR2_X1 U363 ( .A(n302), .B(n301), .ZN(n425) );
  XOR2_X1 U364 ( .A(n303), .B(n425), .Z(n313) );
  XOR2_X1 U365 ( .A(KEYINPUT84), .B(KEYINPUT2), .Z(n305) );
  XNOR2_X1 U366 ( .A(G162GAT), .B(KEYINPUT85), .ZN(n304) );
  XNOR2_X1 U367 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U368 ( .A(n306), .B(KEYINPUT3), .Z(n308) );
  XNOR2_X1 U369 ( .A(G141GAT), .B(G155GAT), .ZN(n307) );
  XNOR2_X1 U370 ( .A(n308), .B(n307), .ZN(n406) );
  XOR2_X1 U371 ( .A(G211GAT), .B(KEYINPUT23), .Z(n310) );
  XNOR2_X1 U372 ( .A(G22GAT), .B(KEYINPUT22), .ZN(n309) );
  XNOR2_X1 U373 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U374 ( .A(n406), .B(n311), .ZN(n312) );
  XNOR2_X1 U375 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U376 ( .A(n315), .B(n314), .ZN(n486) );
  XOR2_X1 U377 ( .A(KEYINPUT28), .B(n486), .Z(n521) );
  INV_X1 U378 ( .A(n521), .ZN(n542) );
  XNOR2_X1 U379 ( .A(G155GAT), .B(G78GAT), .ZN(n316) );
  XOR2_X1 U380 ( .A(G1GAT), .B(G127GAT), .Z(n407) );
  XOR2_X1 U381 ( .A(n316), .B(n407), .Z(n329) );
  XNOR2_X1 U382 ( .A(G22GAT), .B(G15GAT), .ZN(n317) );
  XNOR2_X1 U383 ( .A(n317), .B(KEYINPUT72), .ZN(n336) );
  XOR2_X1 U384 ( .A(KEYINPUT77), .B(n336), .Z(n319) );
  NAND2_X1 U385 ( .A1(G231GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U386 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U387 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n321) );
  XNOR2_X1 U388 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n320) );
  XNOR2_X1 U389 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U390 ( .A(n323), .B(n322), .Z(n327) );
  XOR2_X1 U391 ( .A(G71GAT), .B(G57GAT), .Z(n324) );
  XOR2_X1 U392 ( .A(KEYINPUT13), .B(n324), .Z(n368) );
  XNOR2_X1 U393 ( .A(G8GAT), .B(G183GAT), .ZN(n325) );
  XNOR2_X1 U394 ( .A(n325), .B(G211GAT), .ZN(n432) );
  XNOR2_X1 U395 ( .A(n368), .B(n432), .ZN(n326) );
  XNOR2_X1 U396 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U397 ( .A(n329), .B(n328), .Z(n587) );
  INV_X1 U398 ( .A(n587), .ZN(n507) );
  XOR2_X1 U399 ( .A(KEYINPUT110), .B(n507), .Z(n570) );
  INV_X1 U400 ( .A(KEYINPUT46), .ZN(n371) );
  XOR2_X1 U401 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n331) );
  XNOR2_X1 U402 ( .A(KEYINPUT30), .B(G8GAT), .ZN(n330) );
  XNOR2_X1 U403 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U404 ( .A(KEYINPUT29), .B(KEYINPUT70), .Z(n333) );
  XNOR2_X1 U405 ( .A(G1GAT), .B(KEYINPUT73), .ZN(n332) );
  XNOR2_X1 U406 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U407 ( .A(n335), .B(n334), .ZN(n343) );
  XOR2_X1 U408 ( .A(n336), .B(KEYINPUT69), .Z(n341) );
  XOR2_X1 U409 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n338) );
  XNOR2_X1 U410 ( .A(G50GAT), .B(G43GAT), .ZN(n337) );
  XNOR2_X1 U411 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U412 ( .A(KEYINPUT71), .B(n339), .Z(n390) );
  XNOR2_X1 U413 ( .A(n390), .B(KEYINPUT74), .ZN(n340) );
  XNOR2_X1 U414 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U415 ( .A(n343), .B(n342), .ZN(n349) );
  XOR2_X1 U416 ( .A(G113GAT), .B(G197GAT), .Z(n345) );
  XNOR2_X1 U417 ( .A(G169GAT), .B(G141GAT), .ZN(n344) );
  XNOR2_X1 U418 ( .A(n345), .B(n344), .ZN(n347) );
  XOR2_X1 U419 ( .A(G29GAT), .B(G36GAT), .Z(n346) );
  XNOR2_X1 U420 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U421 ( .A(n349), .B(n348), .ZN(n351) );
  AND2_X1 U422 ( .A1(G229GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U423 ( .A(n351), .B(n350), .ZN(n495) );
  INV_X1 U424 ( .A(n495), .ZN(n579) );
  INV_X1 U425 ( .A(KEYINPUT41), .ZN(n369) );
  XNOR2_X1 U426 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n353) );
  AND2_X1 U427 ( .A1(G230GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U428 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U429 ( .A(n354), .B(KEYINPUT33), .Z(n359) );
  XOR2_X1 U430 ( .A(G64GAT), .B(G92GAT), .Z(n356) );
  XNOR2_X1 U431 ( .A(G176GAT), .B(G204GAT), .ZN(n355) );
  XNOR2_X1 U432 ( .A(n357), .B(n433), .ZN(n358) );
  XNOR2_X1 U433 ( .A(n359), .B(n358), .ZN(n361) );
  INV_X1 U434 ( .A(KEYINPUT75), .ZN(n360) );
  NAND2_X1 U435 ( .A1(n361), .A2(n360), .ZN(n364) );
  INV_X1 U436 ( .A(n361), .ZN(n362) );
  NAND2_X1 U437 ( .A1(n362), .A2(KEYINPUT75), .ZN(n363) );
  NAND2_X1 U438 ( .A1(n364), .A2(n363), .ZN(n366) );
  XOR2_X1 U439 ( .A(G99GAT), .B(G85GAT), .Z(n382) );
  XNOR2_X1 U440 ( .A(G120GAT), .B(n382), .ZN(n365) );
  XNOR2_X1 U441 ( .A(n366), .B(n365), .ZN(n367) );
  NAND2_X1 U442 ( .A1(n579), .A2(n560), .ZN(n370) );
  XNOR2_X1 U443 ( .A(n371), .B(n370), .ZN(n372) );
  NOR2_X1 U444 ( .A1(n570), .A2(n372), .ZN(n373) );
  XNOR2_X1 U445 ( .A(n373), .B(KEYINPUT111), .ZN(n391) );
  XOR2_X1 U446 ( .A(G29GAT), .B(G134GAT), .Z(n408) );
  XOR2_X1 U447 ( .A(G92GAT), .B(G106GAT), .Z(n375) );
  NAND2_X1 U448 ( .A1(G232GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U449 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U450 ( .A(n408), .B(n376), .ZN(n388) );
  XOR2_X1 U451 ( .A(KEYINPUT9), .B(KEYINPUT64), .Z(n378) );
  XNOR2_X1 U452 ( .A(G162GAT), .B(KEYINPUT66), .ZN(n377) );
  XNOR2_X1 U453 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U454 ( .A(G218GAT), .B(n379), .ZN(n381) );
  XOR2_X1 U455 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n384) );
  XOR2_X1 U456 ( .A(G36GAT), .B(G190GAT), .Z(n428) );
  XNOR2_X1 U457 ( .A(n382), .B(n428), .ZN(n383) );
  XNOR2_X1 U458 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U459 ( .A(n388), .B(n387), .ZN(n389) );
  NOR2_X1 U460 ( .A1(n391), .A2(n565), .ZN(n392) );
  XNOR2_X1 U461 ( .A(n392), .B(KEYINPUT112), .ZN(n394) );
  INV_X1 U462 ( .A(KEYINPUT47), .ZN(n393) );
  XNOR2_X1 U463 ( .A(n394), .B(n393), .ZN(n401) );
  XNOR2_X1 U464 ( .A(KEYINPUT36), .B(KEYINPUT98), .ZN(n395) );
  XOR2_X1 U465 ( .A(n395), .B(n565), .Z(n590) );
  NOR2_X1 U466 ( .A1(n507), .A2(n590), .ZN(n396) );
  XOR2_X1 U467 ( .A(KEYINPUT45), .B(n396), .Z(n397) );
  XNOR2_X1 U468 ( .A(n398), .B(KEYINPUT113), .ZN(n399) );
  NOR2_X1 U469 ( .A1(n399), .A2(n579), .ZN(n400) );
  NOR2_X1 U470 ( .A1(n401), .A2(n400), .ZN(n402) );
  XNOR2_X1 U471 ( .A(n402), .B(KEYINPUT48), .ZN(n483) );
  XOR2_X1 U472 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n404) );
  XNOR2_X1 U473 ( .A(KEYINPUT87), .B(KEYINPUT5), .ZN(n403) );
  XNOR2_X1 U474 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U475 ( .A(n406), .B(n405), .ZN(n419) );
  XOR2_X1 U476 ( .A(KEYINPUT88), .B(G57GAT), .Z(n410) );
  XNOR2_X1 U477 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U478 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U479 ( .A(n411), .B(G85GAT), .Z(n417) );
  XNOR2_X1 U480 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n412) );
  XNOR2_X1 U481 ( .A(n412), .B(G120GAT), .ZN(n440) );
  XOR2_X1 U482 ( .A(n440), .B(KEYINPUT4), .Z(n414) );
  NAND2_X1 U483 ( .A1(G225GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U484 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U485 ( .A(G148GAT), .B(n415), .ZN(n416) );
  XNOR2_X1 U486 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U487 ( .A(n419), .B(n418), .ZN(n472) );
  XOR2_X1 U488 ( .A(KEYINPUT89), .B(n472), .Z(n533) );
  XNOR2_X1 U489 ( .A(KEYINPUT81), .B(KEYINPUT19), .ZN(n420) );
  XNOR2_X1 U490 ( .A(n420), .B(KEYINPUT17), .ZN(n424) );
  XNOR2_X1 U491 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n422) );
  XOR2_X1 U492 ( .A(n425), .B(KEYINPUT92), .Z(n427) );
  NAND2_X1 U493 ( .A1(G226GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U494 ( .A(n427), .B(n426), .ZN(n431) );
  XNOR2_X1 U495 ( .A(n428), .B(KEYINPUT91), .ZN(n429) );
  XNOR2_X1 U496 ( .A(n429), .B(KEYINPUT90), .ZN(n430) );
  XOR2_X1 U497 ( .A(n431), .B(n430), .Z(n435) );
  XNOR2_X1 U498 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U499 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U500 ( .A(n439), .B(n436), .Z(n537) );
  XNOR2_X1 U501 ( .A(KEYINPUT27), .B(n537), .ZN(n464) );
  NAND2_X1 U502 ( .A1(n533), .A2(n464), .ZN(n460) );
  XOR2_X1 U503 ( .A(G176GAT), .B(G127GAT), .Z(n438) );
  XNOR2_X1 U504 ( .A(KEYINPUT78), .B(KEYINPUT79), .ZN(n437) );
  XNOR2_X1 U505 ( .A(n438), .B(n437), .ZN(n452) );
  XNOR2_X1 U506 ( .A(G15GAT), .B(n439), .ZN(n448) );
  XOR2_X1 U507 ( .A(G71GAT), .B(n440), .Z(n446) );
  XOR2_X1 U508 ( .A(G183GAT), .B(KEYINPUT20), .Z(n442) );
  XNOR2_X1 U509 ( .A(G43GAT), .B(G190GAT), .ZN(n441) );
  XNOR2_X1 U510 ( .A(n442), .B(n441), .ZN(n444) );
  XOR2_X1 U511 ( .A(G134GAT), .B(G99GAT), .Z(n443) );
  XNOR2_X1 U512 ( .A(n444), .B(n443), .ZN(n445) );
  NAND2_X1 U513 ( .A1(G227GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U514 ( .A(n450), .B(n449), .ZN(n451) );
  NAND2_X1 U515 ( .A1(n554), .A2(n540), .ZN(n453) );
  XNOR2_X1 U516 ( .A(KEYINPUT114), .B(n453), .ZN(n454) );
  NAND2_X1 U517 ( .A1(n551), .A2(n570), .ZN(n458) );
  XOR2_X1 U518 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n456) );
  INV_X1 U519 ( .A(G127GAT), .ZN(n455) );
  XNOR2_X1 U520 ( .A(n458), .B(n457), .ZN(G1342GAT) );
  NAND2_X1 U521 ( .A1(n495), .A2(n560), .ZN(n459) );
  XNOR2_X1 U522 ( .A(n459), .B(KEYINPUT102), .ZN(n532) );
  NOR2_X1 U523 ( .A1(n542), .A2(n460), .ZN(n461) );
  XNOR2_X1 U524 ( .A(n461), .B(KEYINPUT93), .ZN(n462) );
  NOR2_X1 U525 ( .A1(n540), .A2(n462), .ZN(n474) );
  INV_X1 U526 ( .A(n540), .ZN(n517) );
  NAND2_X1 U527 ( .A1(n486), .A2(n517), .ZN(n463) );
  XOR2_X1 U528 ( .A(n463), .B(KEYINPUT26), .Z(n578) );
  NAND2_X1 U529 ( .A1(n578), .A2(n464), .ZN(n469) );
  XNOR2_X1 U530 ( .A(KEYINPUT25), .B(KEYINPUT94), .ZN(n467) );
  INV_X1 U531 ( .A(n537), .ZN(n515) );
  NOR2_X1 U532 ( .A1(n517), .A2(n515), .ZN(n465) );
  NOR2_X1 U533 ( .A1(n486), .A2(n465), .ZN(n466) );
  XNOR2_X1 U534 ( .A(n467), .B(n466), .ZN(n468) );
  NAND2_X1 U535 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U536 ( .A(n470), .B(KEYINPUT95), .ZN(n471) );
  NOR2_X1 U537 ( .A1(n472), .A2(n471), .ZN(n473) );
  NOR2_X1 U538 ( .A1(n565), .A2(n507), .ZN(n475) );
  XOR2_X1 U539 ( .A(KEYINPUT16), .B(n475), .Z(n476) );
  NOR2_X1 U540 ( .A1(n505), .A2(n476), .ZN(n477) );
  XOR2_X1 U541 ( .A(KEYINPUT96), .B(n477), .Z(n496) );
  XOR2_X1 U542 ( .A(KEYINPUT103), .B(n478), .Z(n528) );
  NAND2_X1 U543 ( .A1(n528), .A2(n542), .ZN(n482) );
  XOR2_X1 U544 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n480) );
  XNOR2_X1 U545 ( .A(n484), .B(KEYINPUT54), .ZN(n485) );
  INV_X1 U546 ( .A(n533), .ZN(n512) );
  NAND2_X1 U547 ( .A1(n485), .A2(n512), .ZN(n576) );
  NOR2_X1 U548 ( .A1(n486), .A2(n576), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n487), .B(KEYINPUT55), .ZN(n488) );
  NOR2_X2 U550 ( .A1(n517), .A2(n488), .ZN(n571) );
  NAND2_X1 U551 ( .A1(n571), .A2(n565), .ZN(n490) );
  NAND2_X1 U552 ( .A1(n571), .A2(n560), .ZN(n494) );
  XOR2_X1 U553 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n492) );
  XNOR2_X1 U554 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(G1349GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT34), .B(KEYINPUT97), .Z(n498) );
  OR2_X1 U558 ( .A1(n495), .A2(n582), .ZN(n509) );
  NOR2_X1 U559 ( .A1(n496), .A2(n509), .ZN(n503) );
  NAND2_X1 U560 ( .A1(n503), .A2(n533), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U562 ( .A(G1GAT), .B(n499), .ZN(G1324GAT) );
  NAND2_X1 U563 ( .A1(n503), .A2(n537), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n500), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U565 ( .A(G15GAT), .B(KEYINPUT35), .Z(n502) );
  NAND2_X1 U566 ( .A1(n503), .A2(n540), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n502), .B(n501), .ZN(G1326GAT) );
  NAND2_X1 U568 ( .A1(n503), .A2(n542), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n504), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U570 ( .A1(n505), .A2(n590), .ZN(n506) );
  NAND2_X1 U571 ( .A1(n507), .A2(n506), .ZN(n508) );
  XOR2_X1 U572 ( .A(KEYINPUT37), .B(n508), .Z(n531) );
  NOR2_X1 U573 ( .A1(n531), .A2(n509), .ZN(n511) );
  XNOR2_X1 U574 ( .A(KEYINPUT99), .B(KEYINPUT38), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(n522) );
  NOR2_X1 U576 ( .A1(n522), .A2(n512), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n513), .B(KEYINPUT39), .ZN(n514) );
  XNOR2_X1 U578 ( .A(G29GAT), .B(n514), .ZN(G1328GAT) );
  NOR2_X1 U579 ( .A1(n522), .A2(n515), .ZN(n516) );
  XOR2_X1 U580 ( .A(G36GAT), .B(n516), .Z(G1329GAT) );
  XNOR2_X1 U581 ( .A(KEYINPUT100), .B(KEYINPUT40), .ZN(n519) );
  NOR2_X1 U582 ( .A1(n517), .A2(n522), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U584 ( .A(G43GAT), .B(n520), .Z(G1330GAT) );
  NOR2_X1 U585 ( .A1(n522), .A2(n521), .ZN(n524) );
  XNOR2_X1 U586 ( .A(G50GAT), .B(KEYINPUT101), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n524), .B(n523), .ZN(G1331GAT) );
  NAND2_X1 U588 ( .A1(n528), .A2(n533), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n525), .B(KEYINPUT42), .ZN(n526) );
  XNOR2_X1 U590 ( .A(G57GAT), .B(n526), .ZN(G1332GAT) );
  NAND2_X1 U591 ( .A1(n537), .A2(n528), .ZN(n527) );
  XNOR2_X1 U592 ( .A(G64GAT), .B(n527), .ZN(G1333GAT) );
  NAND2_X1 U593 ( .A1(n540), .A2(n528), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n529), .B(KEYINPUT104), .ZN(n530) );
  XNOR2_X1 U595 ( .A(G71GAT), .B(n530), .ZN(G1334GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n535) );
  NOR2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n543), .A2(n533), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U600 ( .A(G85GAT), .B(n536), .ZN(G1336GAT) );
  NAND2_X1 U601 ( .A1(n543), .A2(n537), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n538), .B(KEYINPUT108), .ZN(n539) );
  XNOR2_X1 U603 ( .A(G92GAT), .B(n539), .ZN(G1337GAT) );
  NAND2_X1 U604 ( .A1(n540), .A2(n543), .ZN(n541) );
  XNOR2_X1 U605 ( .A(n541), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n545) );
  NAND2_X1 U607 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U609 ( .A(G106GAT), .B(n546), .ZN(G1339GAT) );
  NAND2_X1 U610 ( .A1(n579), .A2(n551), .ZN(n547) );
  XNOR2_X1 U611 ( .A(G113GAT), .B(n547), .ZN(G1340GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n549) );
  NAND2_X1 U613 ( .A1(n551), .A2(n560), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U615 ( .A(G120GAT), .B(n550), .Z(G1341GAT) );
  XOR2_X1 U616 ( .A(G134GAT), .B(KEYINPUT51), .Z(n553) );
  NAND2_X1 U617 ( .A1(n551), .A2(n565), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  XOR2_X1 U619 ( .A(G141GAT), .B(KEYINPUT117), .Z(n556) );
  AND2_X1 U620 ( .A1(n578), .A2(n554), .ZN(n566) );
  NAND2_X1 U621 ( .A1(n566), .A2(n579), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1344GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n558) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U626 ( .A(KEYINPUT53), .B(n559), .Z(n562) );
  NAND2_X1 U627 ( .A1(n566), .A2(n560), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1345GAT) );
  NAND2_X1 U629 ( .A1(n587), .A2(n566), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(KEYINPUT120), .ZN(n564) );
  XNOR2_X1 U631 ( .A(G155GAT), .B(n564), .ZN(G1346GAT) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U634 ( .A(G169GAT), .B(KEYINPUT121), .Z(n569) );
  NAND2_X1 U635 ( .A1(n571), .A2(n579), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G1348GAT) );
  XOR2_X1 U637 ( .A(G183GAT), .B(KEYINPUT123), .Z(n573) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1350GAT) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n574), .B(KEYINPUT59), .ZN(n575) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(n575), .Z(n581) );
  INV_X1 U643 ( .A(n576), .ZN(n577) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n589) );
  INV_X1 U645 ( .A(n589), .ZN(n586) );
  NAND2_X1 U646 ( .A1(n586), .A2(n579), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n584) );
  NAND2_X1 U649 ( .A1(n586), .A2(n582), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n585) );
  XOR2_X1 U651 ( .A(G204GAT), .B(n585), .Z(G1353GAT) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n592) );
  XNOR2_X1 U655 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n592), .B(n591), .ZN(n593) );
  XOR2_X1 U657 ( .A(G218GAT), .B(n593), .Z(G1355GAT) );
endmodule

