//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 0 1 0 0 1 1 1 0 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n553, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n605, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT65), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(new_n461), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n463), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n461), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(G160));
  INV_X1    g045(.A(new_n464), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G136), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n463), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  NOR2_X1   g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI21_X1  g050(.A(G2104), .B1(new_n461), .B2(G112), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n472), .B(new_n474), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  XOR2_X1   g052(.A(new_n477), .B(KEYINPUT67), .Z(G162));
  AND2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  OAI211_X1 g055(.A(G138), .B(new_n461), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n463), .A2(KEYINPUT69), .A3(G138), .A4(new_n461), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT70), .A4(KEYINPUT4), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n463), .A2(G126), .A3(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT68), .B1(new_n461), .B2(G114), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT68), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n488), .A2(new_n489), .A3(G2105), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n487), .A2(new_n490), .A3(G2104), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AND3_X1   g069(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n481), .B2(KEYINPUT4), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n485), .B(new_n494), .C1(new_n495), .C2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G651), .ZN(new_n501));
  XNOR2_X1  g076(.A(new_n501), .B(KEYINPUT71), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(G50), .A2(new_n507), .B1(new_n512), .B2(G88), .ZN(new_n513));
  INV_X1    g088(.A(G62), .ZN(new_n514));
  OR3_X1    g089(.A1(new_n511), .A2(KEYINPUT72), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  OAI21_X1  g091(.A(KEYINPUT72), .B1(new_n511), .B2(new_n514), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n513), .A2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  NAND2_X1  g096(.A1(new_n507), .A2(G51), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n512), .A2(G89), .ZN(new_n523));
  XOR2_X1   g098(.A(KEYINPUT73), .B(KEYINPUT7), .Z(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n524), .B(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n511), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n527), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n522), .A2(new_n523), .A3(new_n526), .A4(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(G168));
  AOI22_X1  g105(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(new_n503), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n507), .A2(G52), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n512), .A2(G90), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n535), .B1(new_n533), .B2(new_n534), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n532), .B1(new_n537), .B2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n511), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT75), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT76), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n512), .A2(G81), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n507), .A2(G43), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  XOR2_X1   g130(.A(new_n555), .B(KEYINPUT77), .Z(G188));
  NAND4_X1  g131(.A1(new_n502), .A2(G53), .A3(G543), .A4(new_n504), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n502), .A2(G91), .A3(new_n527), .A4(new_n504), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT78), .ZN(new_n562));
  OR2_X1    g137(.A1(KEYINPUT79), .A2(G65), .ZN(new_n563));
  NAND2_X1  g138(.A1(KEYINPUT79), .A2(G65), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n527), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT80), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT80), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n565), .A2(new_n569), .A3(new_n566), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(G651), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n560), .A2(new_n562), .A3(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT81), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n560), .A2(new_n562), .A3(KEYINPUT81), .A4(new_n571), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(G299));
  XNOR2_X1  g151(.A(new_n529), .B(KEYINPUT82), .ZN(G286));
  NAND2_X1  g152(.A1(new_n507), .A2(G49), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n512), .A2(G87), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  AND2_X1   g156(.A1(new_n527), .A2(G61), .ZN(new_n582));
  AND2_X1   g157(.A1(G73), .A2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  XOR2_X1   g159(.A(new_n584), .B(KEYINPUT83), .Z(new_n585));
  AOI22_X1  g160(.A1(G48), .A2(new_n507), .B1(new_n512), .B2(G86), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(new_n512), .A2(G85), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n507), .A2(G47), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n527), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n588), .B(new_n589), .C1(new_n503), .C2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n512), .A2(G92), .ZN(new_n593));
  XOR2_X1   g168(.A(new_n593), .B(KEYINPUT10), .Z(new_n594));
  NAND2_X1  g169(.A1(new_n507), .A2(G54), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n527), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(new_n503), .ZN(new_n597));
  AND3_X1   g172(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n592), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n592), .B1(new_n598), .B2(G868), .ZN(G321));
  NAND2_X1  g175(.A1(G286), .A2(G868), .ZN(new_n601));
  INV_X1    g176(.A(G299), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G297));
  OAI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n598), .B1(new_n605), .B2(G860), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT84), .ZN(G148));
  NAND2_X1  g182(.A1(new_n598), .A2(new_n605), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n473), .A2(G123), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT86), .Z(new_n613));
  NAND2_X1  g188(.A1(new_n471), .A2(G135), .ZN(new_n614));
  NOR2_X1   g189(.A1(G99), .A2(G2105), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(new_n461), .B2(G111), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n613), .B(new_n614), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G2096), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT85), .B(KEYINPUT12), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n620), .B(new_n621), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2100), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT87), .ZN(G156));
  XNOR2_X1  g201(.A(G2451), .B(G2454), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT16), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2443), .B(G2446), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G1341), .B(G1348), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2435), .ZN(new_n634));
  XOR2_X1   g209(.A(G2427), .B(G2438), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(KEYINPUT14), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n632), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G14), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT88), .Z(G401));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT89), .ZN(new_n642));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  XNOR2_X1  g218(.A(G2072), .B(G2078), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT18), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n642), .B(KEYINPUT90), .ZN(new_n647));
  INV_X1    g222(.A(new_n643), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT17), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(new_n644), .Z(new_n651));
  NOR2_X1   g226(.A1(new_n647), .A2(new_n648), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n646), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(new_n618), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(G2100), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n653), .B(G2096), .ZN(new_n656));
  INV_X1    g231(.A(G2100), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G227));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1956), .B(G2474), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT91), .ZN(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n661), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n663), .A2(new_n664), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n670), .A2(new_n667), .A3(new_n665), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n665), .A2(new_n661), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n672), .A2(new_n669), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n668), .B(new_n671), .C1(new_n673), .C2(new_n667), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT92), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(G229));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G24), .ZN(new_n685));
  XOR2_X1   g260(.A(G290), .B(KEYINPUT95), .Z(new_n686));
  OAI21_X1  g261(.A(new_n685), .B1(new_n686), .B2(new_n684), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT96), .B(G1986), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n684), .A2(G6), .ZN(new_n690));
  INV_X1    g265(.A(G305), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(new_n684), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT97), .B(KEYINPUT32), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1981), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n684), .A2(G23), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT98), .ZN(new_n697));
  NAND2_X1  g272(.A1(G288), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g273(.A1(new_n578), .A2(new_n579), .A3(KEYINPUT98), .A4(new_n580), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n696), .B1(new_n700), .B2(new_n684), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT33), .B(G1976), .Z(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n684), .A2(G22), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G166), .B2(new_n684), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(G1971), .Z(new_n707));
  NAND4_X1  g282(.A1(new_n695), .A2(new_n703), .A3(new_n704), .A4(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n689), .B1(new_n708), .B2(KEYINPUT34), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n473), .A2(G119), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT93), .Z(new_n711));
  OR2_X1    g286(.A1(G95), .A2(G2105), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n712), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n471), .A2(G131), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n711), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  MUX2_X1   g290(.A(G25), .B(new_n715), .S(G29), .Z(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT35), .B(G1991), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT94), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n716), .B(new_n718), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n709), .B(new_n719), .C1(KEYINPUT34), .C2(new_n708), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT36), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT101), .B(KEYINPUT24), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G34), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(G29), .ZN(new_n724));
  INV_X1    g299(.A(G160), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(G29), .ZN(new_n726));
  INV_X1    g301(.A(G2084), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n684), .A2(G4), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n598), .B2(new_n684), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n730), .A2(G1348), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n730), .A2(G1348), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G33), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n735), .A2(new_n461), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G139), .B2(new_n471), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT25), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n734), .B1(new_n741), .B2(new_n733), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G2072), .ZN(new_n743));
  INV_X1    g318(.A(G28), .ZN(new_n744));
  AOI21_X1  g319(.A(G29), .B1(new_n744), .B2(KEYINPUT30), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(KEYINPUT30), .B2(new_n744), .ZN(new_n746));
  OR2_X1    g321(.A1(G29), .A2(G32), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT102), .B(KEYINPUT26), .Z(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n471), .A2(G141), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n473), .A2(G129), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n750), .A2(new_n751), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n747), .B1(new_n754), .B2(new_n733), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT27), .B(G1996), .ZN(new_n756));
  OAI221_X1 g331(.A(new_n746), .B1(new_n755), .B2(new_n756), .C1(new_n617), .C2(new_n733), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT100), .B(KEYINPUT28), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n733), .A2(G26), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  AOI22_X1  g335(.A1(G140), .A2(new_n471), .B1(new_n473), .B2(G128), .ZN(new_n761));
  INV_X1    g336(.A(G2104), .ZN(new_n762));
  OR2_X1    g337(.A1(G104), .A2(G2105), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT99), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI221_X1 g340(.A(new_n765), .B1(new_n764), .B2(new_n763), .C1(G116), .C2(new_n461), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n761), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n760), .B1(new_n767), .B2(G29), .ZN(new_n768));
  INV_X1    g343(.A(G2067), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n757), .A2(new_n770), .ZN(new_n771));
  NOR4_X1   g346(.A1(new_n731), .A2(new_n732), .A3(new_n743), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n755), .A2(new_n756), .ZN(new_n773));
  NAND2_X1  g348(.A1(G168), .A2(G16), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G16), .B2(G21), .ZN(new_n775));
  INV_X1    g350(.A(G1966), .ZN(new_n776));
  OAI221_X1 g351(.A(new_n773), .B1(new_n727), .B2(new_n726), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G5), .A2(G16), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G171), .B2(G16), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n779), .A2(G1961), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n777), .B(new_n780), .C1(new_n776), .C2(new_n775), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n733), .A2(G35), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G162), .B2(new_n733), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT29), .B(G2090), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n779), .B2(G1961), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT31), .B(G11), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n772), .A2(new_n781), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT103), .B(KEYINPUT23), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n684), .A2(G20), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G299), .B2(G16), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(G1956), .Z(new_n793));
  NOR2_X1   g368(.A1(new_n549), .A2(new_n684), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n684), .B2(G19), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n796), .A2(G1341), .ZN(new_n797));
  NOR2_X1   g372(.A1(G164), .A2(new_n733), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G27), .B2(new_n733), .ZN(new_n799));
  INV_X1    g374(.A(G2078), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  INV_X1    g377(.A(G1341), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n801), .B(new_n802), .C1(new_n795), .C2(new_n803), .ZN(new_n804));
  NOR4_X1   g379(.A1(new_n788), .A2(new_n793), .A3(new_n797), .A4(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n721), .A2(new_n728), .A3(new_n805), .ZN(G150));
  XOR2_X1   g381(.A(G150), .B(KEYINPUT104), .Z(G311));
  NAND2_X1  g382(.A1(new_n512), .A2(G93), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n507), .A2(G55), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n527), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n808), .B(new_n809), .C1(new_n503), .C2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT105), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(G860), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT37), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n598), .A2(G559), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT38), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n546), .A2(new_n547), .A3(new_n548), .A4(new_n811), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n549), .B2(new_n812), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n816), .B(new_n818), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n820), .A2(KEYINPUT106), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n820), .A2(KEYINPUT106), .ZN(new_n822));
  OR3_X1    g397(.A1(new_n821), .A2(new_n822), .A3(G860), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n814), .B1(new_n823), .B2(new_n824), .ZN(G145));
  XNOR2_X1  g400(.A(new_n617), .B(G160), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G162), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n498), .B(new_n754), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n767), .ZN(new_n829));
  INV_X1    g404(.A(new_n741), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n471), .A2(G142), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n473), .A2(G130), .ZN(new_n834));
  NOR2_X1   g409(.A1(G106), .A2(G2105), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n833), .B(new_n834), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n715), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n622), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(KEYINPUT107), .B1(new_n832), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n840), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n831), .A2(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n829), .A2(new_n830), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n829), .A2(new_n830), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n840), .A2(new_n844), .A3(KEYINPUT107), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n827), .B1(new_n841), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G37), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n827), .B1(new_n832), .B2(new_n840), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(new_n843), .ZN(new_n851));
  AND3_X1   g426(.A1(new_n848), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g428(.A(new_n818), .B(new_n608), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT108), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(new_n574), .B2(new_n575), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n574), .A2(new_n855), .A3(new_n575), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n602), .A2(new_n598), .A3(new_n855), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n854), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n865), .A2(KEYINPUT41), .A3(new_n861), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(KEYINPUT41), .B1(new_n865), .B2(new_n861), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n854), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n864), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT42), .ZN(new_n871));
  XNOR2_X1  g446(.A(G303), .B(G290), .ZN(new_n872));
  INV_X1    g447(.A(new_n700), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n691), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n875), .A2(KEYINPUT109), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT42), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n864), .A2(new_n869), .A3(new_n877), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n871), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n876), .B1(new_n871), .B2(new_n878), .ZN(new_n880));
  OAI21_X1  g455(.A(G868), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n812), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n881), .B1(G868), .B2(new_n882), .ZN(G295));
  XNOR2_X1  g458(.A(G295), .B(KEYINPUT110), .ZN(G331));
  INV_X1    g459(.A(new_n875), .ZN(new_n885));
  NAND2_X1  g460(.A1(G171), .A2(G286), .ZN(new_n886));
  NAND2_X1  g461(.A1(G301), .A2(G168), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n818), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n882), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT82), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n529), .B(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n887), .B1(new_n892), .B2(G301), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n890), .A2(new_n893), .A3(new_n817), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(new_n860), .B2(new_n862), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n895), .B1(new_n897), .B2(new_n866), .ZN(new_n898));
  AOI22_X1  g473(.A1(new_n888), .A2(new_n894), .B1(new_n865), .B2(new_n861), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n885), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n888), .A2(new_n894), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n867), .B2(new_n868), .ZN(new_n902));
  INV_X1    g477(.A(new_n899), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n902), .A2(new_n875), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n900), .A2(new_n904), .A3(new_n849), .ZN(new_n905));
  XOR2_X1   g480(.A(KEYINPUT111), .B(KEYINPUT43), .Z(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n906), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n900), .A2(new_n904), .A3(new_n849), .A4(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n911), .A2(new_n909), .ZN(new_n912));
  MUX2_X1   g487(.A(new_n910), .B(new_n912), .S(KEYINPUT44), .Z(G397));
  INV_X1    g488(.A(G1384), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT45), .B1(new_n498), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  XOR2_X1   g491(.A(KEYINPUT112), .B(G40), .Z(new_n917));
  NOR2_X1   g492(.A1(new_n725), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n767), .A2(G2067), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n761), .A2(new_n769), .A3(new_n766), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G1996), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n754), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n715), .A2(new_n717), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n715), .A2(new_n717), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g505(.A1(G290), .A2(G1986), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(G290), .A2(G1986), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n920), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT4), .ZN(new_n936));
  INV_X1    g511(.A(new_n497), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n493), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI211_X1 g513(.A(new_n935), .B(G1384), .C1(new_n938), .C2(new_n485), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n939), .A2(new_n915), .A3(new_n919), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n800), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT53), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT50), .ZN(new_n944));
  AOI211_X1 g519(.A(new_n944), .B(G1384), .C1(new_n938), .C2(new_n485), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT50), .B1(new_n498), .B2(new_n914), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n918), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(KEYINPUT121), .A2(G1961), .ZN(new_n948));
  AND2_X1   g523(.A1(KEYINPUT121), .A2(G1961), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n939), .A2(new_n915), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n725), .A2(new_n942), .A3(G2078), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(G40), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n943), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(G171), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n950), .B1(new_n941), .B2(new_n942), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT122), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI211_X1 g533(.A(KEYINPUT122), .B(new_n950), .C1(new_n941), .C2(new_n942), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n943), .A3(new_n959), .ZN(new_n960));
  OAI211_X1 g535(.A(KEYINPUT54), .B(new_n955), .C1(new_n960), .C2(G171), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT114), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n700), .A2(new_n962), .A3(G1976), .ZN(new_n963));
  AOI21_X1  g538(.A(G1384), .B1(new_n938), .B2(new_n485), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n918), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G8), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n963), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n962), .B1(new_n700), .B2(G1976), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT52), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n970), .ZN(new_n972));
  INV_X1    g547(.A(G1976), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT52), .B1(G288), .B2(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n972), .A2(new_n968), .A3(new_n963), .A4(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G1981), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n585), .A2(new_n976), .A3(new_n586), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT49), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n586), .A2(new_n584), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(G1981), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n978), .B1(new_n977), .B2(new_n980), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n968), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n971), .A2(new_n975), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(G303), .A2(G8), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n985), .B(KEYINPUT55), .Z(new_n986));
  XNOR2_X1  g561(.A(KEYINPUT113), .B(G1971), .ZN(new_n987));
  OAI22_X1  g562(.A1(new_n940), .A2(new_n987), .B1(new_n947), .B2(G2090), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n986), .A2(new_n988), .A3(G8), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n986), .B1(new_n988), .B2(G8), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n984), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n961), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n960), .A2(G171), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n954), .A2(G171), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT54), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(G1966), .B1(new_n951), .B2(new_n918), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n727), .B(new_n918), .C1(new_n945), .C2(new_n946), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT117), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT117), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n1001), .B(new_n998), .C1(new_n940), .C2(G1966), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1000), .A2(G168), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1003), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT118), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT119), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n997), .A2(new_n999), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1006), .B1(new_n1007), .B2(new_n967), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n1009));
  NOR2_X1   g584(.A1(G168), .A2(new_n967), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(KEYINPUT119), .B(G8), .C1(new_n997), .C2(new_n999), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT118), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1003), .A2(new_n1014), .A3(KEYINPUT51), .A4(G8), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1005), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT120), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n1010), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1017), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n996), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT123), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n964), .A2(KEYINPUT45), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n916), .A2(new_n1025), .A3(new_n918), .ZN(new_n1026));
  XNOR2_X1  g601(.A(KEYINPUT58), .B(G1341), .ZN(new_n1027));
  OAI22_X1  g602(.A1(new_n1026), .A2(G1996), .B1(new_n966), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n549), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(KEYINPUT59), .ZN(new_n1030));
  INV_X1    g605(.A(new_n947), .ZN(new_n1031));
  XOR2_X1   g606(.A(KEYINPUT56), .B(G2072), .Z(new_n1032));
  OAI22_X1  g607(.A1(new_n1031), .A2(G1956), .B1(new_n1026), .B2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n572), .B(KEYINPUT57), .ZN(new_n1034));
  OR2_X1    g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT61), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1036), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1030), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI22_X1  g617(.A1(new_n1031), .A2(G1348), .B1(G2067), .B2(new_n965), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1043), .A2(new_n598), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1043), .A2(new_n598), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT60), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(KEYINPUT116), .B(new_n1030), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1047));
  OR3_X1    g622(.A1(new_n1043), .A2(KEYINPUT60), .A3(new_n858), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1042), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1035), .A2(new_n1044), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(new_n1050), .A3(new_n1037), .ZN(new_n1051));
  OAI211_X1 g626(.A(KEYINPUT123), .B(new_n996), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1024), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT62), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT120), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT62), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n993), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1054), .A2(new_n1059), .A3(new_n1060), .A4(new_n991), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1007), .A2(new_n967), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n991), .A2(new_n892), .A3(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(KEYINPUT63), .ZN(new_n1064));
  INV_X1    g639(.A(new_n989), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(new_n984), .ZN(new_n1066));
  NOR2_X1   g641(.A1(G288), .A2(G1976), .ZN(new_n1067));
  XOR2_X1   g642(.A(new_n1067), .B(KEYINPUT115), .Z(new_n1068));
  OR3_X1    g643(.A1(new_n1068), .A2(new_n981), .A3(new_n982), .ZN(new_n1069));
  AOI211_X1 g644(.A(new_n967), .B(new_n966), .C1(new_n1069), .C2(new_n977), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1064), .A2(new_n1066), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1061), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n934), .B1(new_n1053), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n920), .A2(new_n933), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT124), .B(KEYINPUT48), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1074), .B(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n920), .B2(new_n930), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT46), .ZN(new_n1078));
  INV_X1    g653(.A(new_n920), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1078), .B1(new_n1079), .B2(G1996), .ZN(new_n1080));
  INV_X1    g655(.A(new_n923), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n920), .B1(new_n754), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n920), .A2(KEYINPUT46), .A3(new_n924), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1080), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  XOR2_X1   g659(.A(new_n1084), .B(KEYINPUT47), .Z(new_n1085));
  OAI21_X1  g660(.A(new_n922), .B1(new_n929), .B2(new_n926), .ZN(new_n1086));
  AOI211_X1 g661(.A(new_n1077), .B(new_n1085), .C1(new_n920), .C2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1073), .A2(new_n1087), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g663(.A(new_n852), .ZN(new_n1090));
  INV_X1    g664(.A(KEYINPUT125), .ZN(new_n1091));
  NAND2_X1  g665(.A1(new_n639), .A2(G319), .ZN(new_n1092));
  INV_X1    g666(.A(new_n1092), .ZN(new_n1093));
  NAND4_X1  g667(.A1(new_n659), .A2(new_n1091), .A3(new_n682), .A4(new_n1093), .ZN(new_n1094));
  NAND3_X1  g668(.A1(new_n682), .A2(new_n655), .A3(new_n658), .ZN(new_n1095));
  OAI21_X1  g669(.A(KEYINPUT125), .B1(new_n1095), .B2(new_n1092), .ZN(new_n1096));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  AND4_X1   g671(.A1(KEYINPUT126), .A2(new_n910), .A3(new_n1090), .A4(new_n1097), .ZN(new_n1098));
  AOI21_X1  g672(.A(new_n852), .B1(new_n907), .B2(new_n909), .ZN(new_n1099));
  AOI21_X1  g673(.A(KEYINPUT126), .B1(new_n1099), .B2(new_n1097), .ZN(new_n1100));
  OAI21_X1  g674(.A(KEYINPUT127), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g675(.A1(new_n910), .A2(new_n1090), .A3(new_n1097), .ZN(new_n1102));
  INV_X1    g676(.A(KEYINPUT126), .ZN(new_n1103));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g678(.A(KEYINPUT127), .ZN(new_n1105));
  NAND3_X1  g679(.A1(new_n1099), .A2(KEYINPUT126), .A3(new_n1097), .ZN(new_n1106));
  NAND3_X1  g680(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g681(.A1(new_n1101), .A2(new_n1107), .ZN(G308));
  NAND2_X1  g682(.A1(new_n1104), .A2(new_n1106), .ZN(G225));
endmodule


