

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592;

  XOR2_X1 U320 ( .A(G36GAT), .B(G190GAT), .Z(n354) );
  NOR2_X2 U321 ( .A1(n484), .A2(n530), .ZN(n573) );
  NOR2_X1 U322 ( .A1(n373), .A2(n372), .ZN(n375) );
  INV_X1 U323 ( .A(G176GAT), .ZN(n314) );
  XNOR2_X1 U324 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U325 ( .A(n423), .B(n422), .ZN(n424) );
  NOR2_X1 U326 ( .A1(n401), .A2(n400), .ZN(n402) );
  XNOR2_X1 U327 ( .A(n392), .B(n316), .ZN(n317) );
  XNOR2_X1 U328 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U329 ( .A(n351), .B(KEYINPUT96), .ZN(n352) );
  XNOR2_X1 U330 ( .A(n312), .B(n311), .ZN(n319) );
  XNOR2_X1 U331 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U332 ( .A(n353), .B(n352), .ZN(n571) );
  XNOR2_X1 U333 ( .A(n319), .B(n318), .ZN(n324) );
  XNOR2_X1 U334 ( .A(n436), .B(n435), .ZN(n580) );
  NOR2_X1 U335 ( .A1(n507), .A2(n518), .ZN(n456) );
  XNOR2_X1 U336 ( .A(n456), .B(n455), .ZN(n533) );
  XNOR2_X1 U337 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U338 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U339 ( .A(n457), .B(G99GAT), .ZN(n458) );
  XNOR2_X1 U340 ( .A(n492), .B(n491), .ZN(G1351GAT) );
  XNOR2_X1 U341 ( .A(n459), .B(n458), .ZN(G1338GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT11), .B(KEYINPUT77), .Z(n289) );
  XOR2_X1 U343 ( .A(G99GAT), .B(G85GAT), .Z(n427) );
  XNOR2_X1 U344 ( .A(n427), .B(n354), .ZN(n288) );
  XNOR2_X1 U345 ( .A(n289), .B(n288), .ZN(n290) );
  XOR2_X1 U346 ( .A(n290), .B(KEYINPUT65), .Z(n295) );
  XOR2_X1 U347 ( .A(KEYINPUT76), .B(KEYINPUT9), .Z(n292) );
  XNOR2_X1 U348 ( .A(G134GAT), .B(KEYINPUT10), .ZN(n291) );
  XNOR2_X1 U349 ( .A(n292), .B(n291), .ZN(n293) );
  XNOR2_X1 U350 ( .A(G218GAT), .B(n293), .ZN(n294) );
  XNOR2_X1 U351 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U352 ( .A(G92GAT), .B(G106GAT), .Z(n297) );
  NAND2_X1 U353 ( .A1(G232GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U354 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U355 ( .A(n299), .B(n298), .Z(n305) );
  XNOR2_X1 U356 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n300), .B(G29GAT), .ZN(n301) );
  XOR2_X1 U358 ( .A(n301), .B(KEYINPUT8), .Z(n303) );
  XNOR2_X1 U359 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n303), .B(n302), .ZN(n452) );
  XOR2_X1 U361 ( .A(G50GAT), .B(G162GAT), .Z(n347) );
  XNOR2_X1 U362 ( .A(n452), .B(n347), .ZN(n304) );
  XNOR2_X1 U363 ( .A(n305), .B(n304), .ZN(n558) );
  XOR2_X1 U364 ( .A(KEYINPUT36), .B(n558), .Z(n590) );
  XOR2_X1 U365 ( .A(KEYINPUT86), .B(G99GAT), .Z(n307) );
  XOR2_X1 U366 ( .A(G15GAT), .B(G127GAT), .Z(n403) );
  XOR2_X1 U367 ( .A(G120GAT), .B(G71GAT), .Z(n429) );
  XNOR2_X1 U368 ( .A(n403), .B(n429), .ZN(n306) );
  XNOR2_X1 U369 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U370 ( .A(n308), .B(G190GAT), .Z(n312) );
  XOR2_X1 U371 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n310) );
  XNOR2_X1 U372 ( .A(KEYINPUT84), .B(KEYINPUT82), .ZN(n309) );
  XNOR2_X1 U373 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U374 ( .A(G113GAT), .B(G134GAT), .ZN(n313) );
  XNOR2_X1 U375 ( .A(n313), .B(KEYINPUT0), .ZN(n392) );
  NAND2_X1 U376 ( .A1(G227GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U377 ( .A(G43GAT), .B(n317), .ZN(n318) );
  XOR2_X1 U378 ( .A(KEYINPUT85), .B(G183GAT), .Z(n321) );
  XNOR2_X1 U379 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n320) );
  XNOR2_X1 U380 ( .A(n321), .B(n320), .ZN(n323) );
  XOR2_X1 U381 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n322) );
  XNOR2_X1 U382 ( .A(n323), .B(n322), .ZN(n368) );
  XNOR2_X1 U383 ( .A(n324), .B(n368), .ZN(n487) );
  INV_X1 U384 ( .A(n487), .ZN(n535) );
  XOR2_X1 U385 ( .A(KEYINPUT89), .B(G218GAT), .Z(n326) );
  XNOR2_X1 U386 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n325) );
  XNOR2_X1 U387 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U388 ( .A(G197GAT), .B(n327), .Z(n365) );
  INV_X1 U389 ( .A(KEYINPUT87), .ZN(n331) );
  XOR2_X1 U390 ( .A(G204GAT), .B(KEYINPUT22), .Z(n329) );
  XNOR2_X1 U391 ( .A(KEYINPUT92), .B(KEYINPUT24), .ZN(n328) );
  XNOR2_X1 U392 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U393 ( .A(n331), .B(n330), .ZN(n333) );
  NAND2_X1 U394 ( .A1(G228GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U395 ( .A(n333), .B(n332), .ZN(n336) );
  INV_X1 U396 ( .A(n336), .ZN(n334) );
  NAND2_X1 U397 ( .A1(n334), .A2(KEYINPUT88), .ZN(n338) );
  INV_X1 U398 ( .A(KEYINPUT88), .ZN(n335) );
  NAND2_X1 U399 ( .A1(n336), .A2(n335), .ZN(n337) );
  NAND2_X1 U400 ( .A1(n338), .A2(n337), .ZN(n343) );
  XOR2_X1 U401 ( .A(KEYINPUT91), .B(KEYINPUT2), .Z(n340) );
  XNOR2_X1 U402 ( .A(KEYINPUT90), .B(G155GAT), .ZN(n339) );
  XNOR2_X1 U403 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U404 ( .A(KEYINPUT3), .B(n341), .Z(n391) );
  XNOR2_X1 U405 ( .A(n391), .B(KEYINPUT23), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n343), .B(n342), .ZN(n346) );
  XOR2_X1 U407 ( .A(G78GAT), .B(G148GAT), .Z(n345) );
  XNOR2_X1 U408 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n344) );
  XNOR2_X1 U409 ( .A(n345), .B(n344), .ZN(n428) );
  XOR2_X1 U410 ( .A(n346), .B(n428), .Z(n349) );
  XOR2_X1 U411 ( .A(G141GAT), .B(G22GAT), .Z(n439) );
  XNOR2_X1 U412 ( .A(n439), .B(n347), .ZN(n348) );
  XNOR2_X1 U413 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U414 ( .A(n365), .B(n350), .ZN(n398) );
  NOR2_X1 U415 ( .A1(n535), .A2(n398), .ZN(n353) );
  INV_X1 U416 ( .A(KEYINPUT26), .ZN(n351) );
  XOR2_X1 U417 ( .A(n354), .B(KEYINPUT95), .Z(n356) );
  NAND2_X1 U418 ( .A1(G226GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U419 ( .A(n356), .B(n355), .ZN(n364) );
  INV_X1 U420 ( .A(KEYINPUT74), .ZN(n357) );
  NAND2_X1 U421 ( .A1(G92GAT), .A2(n357), .ZN(n360) );
  INV_X1 U422 ( .A(G92GAT), .ZN(n358) );
  NAND2_X1 U423 ( .A1(n358), .A2(KEYINPUT74), .ZN(n359) );
  NAND2_X1 U424 ( .A1(n360), .A2(n359), .ZN(n362) );
  XNOR2_X1 U425 ( .A(G176GAT), .B(G64GAT), .ZN(n361) );
  XNOR2_X1 U426 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U427 ( .A(G204GAT), .B(n363), .Z(n425) );
  XOR2_X1 U428 ( .A(n364), .B(n425), .Z(n367) );
  XNOR2_X1 U429 ( .A(G8GAT), .B(n365), .ZN(n366) );
  XNOR2_X1 U430 ( .A(n367), .B(n366), .ZN(n369) );
  XNOR2_X1 U431 ( .A(n369), .B(n368), .ZN(n532) );
  XOR2_X1 U432 ( .A(n532), .B(KEYINPUT27), .Z(n397) );
  NOR2_X1 U433 ( .A1(n571), .A2(n397), .ZN(n373) );
  NAND2_X1 U434 ( .A1(n535), .A2(n532), .ZN(n370) );
  NAND2_X1 U435 ( .A1(n398), .A2(n370), .ZN(n371) );
  XNOR2_X1 U436 ( .A(n371), .B(KEYINPUT25), .ZN(n372) );
  INV_X1 U437 ( .A(KEYINPUT97), .ZN(n374) );
  XNOR2_X1 U438 ( .A(n375), .B(n374), .ZN(n395) );
  XOR2_X1 U439 ( .A(G148GAT), .B(G120GAT), .Z(n377) );
  XNOR2_X1 U440 ( .A(G141GAT), .B(G1GAT), .ZN(n376) );
  XNOR2_X1 U441 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U442 ( .A(KEYINPUT93), .B(KEYINPUT6), .Z(n379) );
  XNOR2_X1 U443 ( .A(G57GAT), .B(KEYINPUT1), .ZN(n378) );
  XNOR2_X1 U444 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U445 ( .A(n381), .B(n380), .Z(n386) );
  XOR2_X1 U446 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n383) );
  NAND2_X1 U447 ( .A1(G225GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U448 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U449 ( .A(KEYINPUT4), .B(n384), .ZN(n385) );
  XNOR2_X1 U450 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U451 ( .A(G85GAT), .B(G162GAT), .Z(n388) );
  XNOR2_X1 U452 ( .A(G29GAT), .B(G127GAT), .ZN(n387) );
  XNOR2_X1 U453 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U454 ( .A(n390), .B(n389), .Z(n394) );
  XNOR2_X1 U455 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n394), .B(n393), .ZN(n530) );
  NOR2_X1 U457 ( .A1(n395), .A2(n530), .ZN(n401) );
  INV_X1 U458 ( .A(n530), .ZN(n396) );
  NOR2_X1 U459 ( .A1(n397), .A2(n396), .ZN(n549) );
  XNOR2_X1 U460 ( .A(KEYINPUT28), .B(KEYINPUT66), .ZN(n399) );
  XNOR2_X1 U461 ( .A(n399), .B(n398), .ZN(n460) );
  NAND2_X1 U462 ( .A1(n549), .A2(n460), .ZN(n537) );
  NOR2_X1 U463 ( .A1(n535), .A2(n537), .ZN(n400) );
  XNOR2_X1 U464 ( .A(KEYINPUT98), .B(n402), .ZN(n495) );
  NOR2_X1 U465 ( .A1(n590), .A2(n495), .ZN(n420) );
  XOR2_X1 U466 ( .A(KEYINPUT13), .B(G57GAT), .Z(n423) );
  XOR2_X1 U467 ( .A(n423), .B(G71GAT), .Z(n405) );
  XNOR2_X1 U468 ( .A(G183GAT), .B(n403), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U470 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n407) );
  NAND2_X1 U471 ( .A1(G231GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U473 ( .A(n409), .B(n408), .Z(n411) );
  XOR2_X1 U474 ( .A(G8GAT), .B(G1GAT), .Z(n438) );
  XNOR2_X1 U475 ( .A(n438), .B(KEYINPUT12), .ZN(n410) );
  XNOR2_X1 U476 ( .A(n411), .B(n410), .ZN(n419) );
  XOR2_X1 U477 ( .A(G78GAT), .B(G155GAT), .Z(n413) );
  XNOR2_X1 U478 ( .A(G22GAT), .B(G211GAT), .ZN(n412) );
  XNOR2_X1 U479 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U480 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n415) );
  XNOR2_X1 U481 ( .A(G64GAT), .B(KEYINPUT78), .ZN(n414) );
  XNOR2_X1 U482 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U483 ( .A(n417), .B(n416), .Z(n418) );
  XNOR2_X1 U484 ( .A(n419), .B(n418), .ZN(n584) );
  NAND2_X1 U485 ( .A1(n420), .A2(n584), .ZN(n421) );
  XOR2_X1 U486 ( .A(KEYINPUT37), .B(n421), .Z(n507) );
  XOR2_X1 U487 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n422) );
  XOR2_X1 U488 ( .A(n427), .B(n426), .Z(n436) );
  XNOR2_X1 U489 ( .A(n429), .B(n428), .ZN(n434) );
  XOR2_X1 U490 ( .A(KEYINPUT31), .B(KEYINPUT72), .Z(n431) );
  NAND2_X1 U491 ( .A1(G230GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U492 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U493 ( .A(KEYINPUT75), .B(n432), .ZN(n433) );
  XNOR2_X1 U494 ( .A(n580), .B(KEYINPUT64), .ZN(n437) );
  XNOR2_X1 U495 ( .A(n437), .B(KEYINPUT41), .ZN(n563) );
  XOR2_X1 U496 ( .A(G15GAT), .B(G113GAT), .Z(n441) );
  XNOR2_X1 U497 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U499 ( .A(n442), .B(G36GAT), .Z(n447) );
  XOR2_X1 U500 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n444) );
  XNOR2_X1 U501 ( .A(G169GAT), .B(G197GAT), .ZN(n443) );
  XNOR2_X1 U502 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U503 ( .A(n445), .B(G50GAT), .ZN(n446) );
  XNOR2_X1 U504 ( .A(n447), .B(n446), .ZN(n451) );
  XOR2_X1 U505 ( .A(KEYINPUT71), .B(KEYINPUT68), .Z(n449) );
  NAND2_X1 U506 ( .A1(G229GAT), .A2(G233GAT), .ZN(n448) );
  XNOR2_X1 U507 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U508 ( .A(n451), .B(n450), .Z(n454) );
  XNOR2_X1 U509 ( .A(n452), .B(KEYINPUT29), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n454), .B(n453), .ZN(n561) );
  INV_X1 U511 ( .A(n561), .ZN(n574) );
  NAND2_X1 U512 ( .A1(n563), .A2(n574), .ZN(n518) );
  INV_X1 U513 ( .A(KEYINPUT105), .ZN(n455) );
  NAND2_X1 U514 ( .A1(n533), .A2(n535), .ZN(n459) );
  XOR2_X1 U515 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n457) );
  INV_X1 U516 ( .A(n460), .ZN(n526) );
  NAND2_X1 U517 ( .A1(n533), .A2(n526), .ZN(n464) );
  XOR2_X1 U518 ( .A(KEYINPUT109), .B(KEYINPUT44), .Z(n462) );
  XNOR2_X1 U519 ( .A(G106GAT), .B(KEYINPUT108), .ZN(n461) );
  XNOR2_X1 U520 ( .A(n464), .B(n463), .ZN(G1339GAT) );
  XOR2_X1 U521 ( .A(KEYINPUT118), .B(KEYINPUT55), .Z(n486) );
  XNOR2_X1 U522 ( .A(KEYINPUT54), .B(KEYINPUT117), .ZN(n483) );
  XNOR2_X1 U523 ( .A(KEYINPUT112), .B(KEYINPUT48), .ZN(n481) );
  NAND2_X1 U524 ( .A1(n563), .A2(n561), .ZN(n466) );
  XNOR2_X1 U525 ( .A(KEYINPUT46), .B(KEYINPUT110), .ZN(n465) );
  XNOR2_X1 U526 ( .A(n466), .B(n465), .ZN(n468) );
  INV_X1 U527 ( .A(n584), .ZN(n567) );
  NOR2_X1 U528 ( .A1(n558), .A2(n567), .ZN(n467) );
  AND2_X1 U529 ( .A1(n468), .A2(n467), .ZN(n471) );
  INV_X1 U530 ( .A(n471), .ZN(n470) );
  INV_X1 U531 ( .A(KEYINPUT47), .ZN(n469) );
  NAND2_X1 U532 ( .A1(n470), .A2(n469), .ZN(n473) );
  NAND2_X1 U533 ( .A1(KEYINPUT47), .A2(n471), .ZN(n472) );
  NAND2_X1 U534 ( .A1(n473), .A2(n472), .ZN(n479) );
  NOR2_X1 U535 ( .A1(n590), .A2(n584), .ZN(n474) );
  XNOR2_X1 U536 ( .A(KEYINPUT45), .B(n474), .ZN(n475) );
  NAND2_X1 U537 ( .A1(n475), .A2(n580), .ZN(n476) );
  NOR2_X1 U538 ( .A1(n561), .A2(n476), .ZN(n477) );
  XNOR2_X1 U539 ( .A(KEYINPUT111), .B(n477), .ZN(n478) );
  NAND2_X1 U540 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n481), .B(n480), .ZN(n548) );
  AND2_X1 U542 ( .A1(n532), .A2(n548), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n483), .B(n482), .ZN(n484) );
  NAND2_X1 U544 ( .A1(n573), .A2(n398), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(n488) );
  NOR2_X2 U546 ( .A1(n488), .A2(n487), .ZN(n568) );
  NAND2_X1 U547 ( .A1(n568), .A2(n558), .ZN(n492) );
  XOR2_X1 U548 ( .A(KEYINPUT121), .B(KEYINPUT58), .Z(n490) );
  XNOR2_X1 U549 ( .A(G190GAT), .B(KEYINPUT120), .ZN(n489) );
  NAND2_X1 U550 ( .A1(n561), .A2(n580), .ZN(n508) );
  NOR2_X1 U551 ( .A1(n558), .A2(n584), .ZN(n494) );
  XNOR2_X1 U552 ( .A(KEYINPUT16), .B(KEYINPUT81), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(n496) );
  NOR2_X1 U554 ( .A1(n496), .A2(n495), .ZN(n497) );
  XNOR2_X1 U555 ( .A(KEYINPUT99), .B(n497), .ZN(n519) );
  NOR2_X1 U556 ( .A1(n508), .A2(n519), .ZN(n498) );
  XNOR2_X1 U557 ( .A(n498), .B(KEYINPUT100), .ZN(n505) );
  NAND2_X1 U558 ( .A1(n530), .A2(n505), .ZN(n500) );
  XOR2_X1 U559 ( .A(KEYINPUT34), .B(KEYINPUT101), .Z(n499) );
  XNOR2_X1 U560 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U561 ( .A(G1GAT), .B(n501), .ZN(G1324GAT) );
  NAND2_X1 U562 ( .A1(n505), .A2(n532), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n502), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U564 ( .A(G15GAT), .B(KEYINPUT35), .Z(n504) );
  NAND2_X1 U565 ( .A1(n535), .A2(n505), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n504), .B(n503), .ZN(G1326GAT) );
  NAND2_X1 U567 ( .A1(n526), .A2(n505), .ZN(n506) );
  XNOR2_X1 U568 ( .A(G22GAT), .B(n506), .ZN(G1327GAT) );
  XOR2_X1 U569 ( .A(G29GAT), .B(KEYINPUT39), .Z(n512) );
  NOR2_X1 U570 ( .A1(n508), .A2(n507), .ZN(n510) );
  XNOR2_X1 U571 ( .A(KEYINPUT102), .B(KEYINPUT38), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n510), .B(n509), .ZN(n514) );
  NAND2_X1 U573 ( .A1(n514), .A2(n530), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n512), .B(n511), .ZN(G1328GAT) );
  NAND2_X1 U575 ( .A1(n514), .A2(n532), .ZN(n513) );
  XNOR2_X1 U576 ( .A(n513), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U577 ( .A1(n514), .A2(n535), .ZN(n515) );
  XNOR2_X1 U578 ( .A(n515), .B(KEYINPUT40), .ZN(n516) );
  XNOR2_X1 U579 ( .A(G43GAT), .B(n516), .ZN(G1330GAT) );
  NAND2_X1 U580 ( .A1(n514), .A2(n526), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n517), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U582 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n521) );
  NOR2_X1 U583 ( .A1(n519), .A2(n518), .ZN(n527) );
  NAND2_X1 U584 ( .A1(n530), .A2(n527), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n521), .B(n520), .ZN(G1332GAT) );
  XOR2_X1 U586 ( .A(G64GAT), .B(KEYINPUT103), .Z(n523) );
  NAND2_X1 U587 ( .A1(n527), .A2(n532), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(G1333GAT) );
  NAND2_X1 U589 ( .A1(n527), .A2(n535), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n524), .B(KEYINPUT104), .ZN(n525) );
  XNOR2_X1 U591 ( .A(G71GAT), .B(n525), .ZN(G1334GAT) );
  XOR2_X1 U592 ( .A(G78GAT), .B(KEYINPUT43), .Z(n529) );
  NAND2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n529), .B(n528), .ZN(G1335GAT) );
  NAND2_X1 U595 ( .A1(n533), .A2(n530), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n531), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n534), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U599 ( .A(G113GAT), .B(KEYINPUT113), .Z(n539) );
  NAND2_X1 U600 ( .A1(n535), .A2(n548), .ZN(n536) );
  NOR2_X1 U601 ( .A1(n537), .A2(n536), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n545), .A2(n561), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(G120GAT), .B(KEYINPUT49), .Z(n541) );
  NAND2_X1 U605 ( .A1(n545), .A2(n563), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n543) );
  NAND2_X1 U608 ( .A1(n545), .A2(n567), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U610 ( .A(G127GAT), .B(n544), .Z(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U612 ( .A1(n545), .A2(n558), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U614 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U615 ( .A1(n571), .A2(n550), .ZN(n551) );
  XOR2_X1 U616 ( .A(KEYINPUT115), .B(n551), .Z(n559) );
  NAND2_X1 U617 ( .A1(n561), .A2(n559), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G141GAT), .B(n552), .ZN(G1344GAT) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n556) );
  XOR2_X1 U620 ( .A(KEYINPUT116), .B(KEYINPUT52), .Z(n554) );
  NAND2_X1 U621 ( .A1(n559), .A2(n563), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(G1345GAT) );
  NAND2_X1 U624 ( .A1(n559), .A2(n567), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n557), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n568), .A2(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n565) );
  NAND2_X1 U631 ( .A1(n568), .A2(n563), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(G176GAT), .B(n566), .ZN(G1349GAT) );
  XOR2_X1 U634 ( .A(G183GAT), .B(KEYINPUT119), .Z(n570) );
  NAND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1350GAT) );
  INV_X1 U637 ( .A(n571), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n589) );
  NOR2_X1 U639 ( .A1(n574), .A2(n589), .ZN(n579) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(KEYINPUT59), .B(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n589), .ZN(n582) );
  XNOR2_X1 U646 ( .A(KEYINPUT61), .B(KEYINPUT124), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(n583), .ZN(G1353GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n589), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1354GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n588) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n587) );
  XNOR2_X1 U654 ( .A(n588), .B(n587), .ZN(n592) );
  NOR2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U656 ( .A(n592), .B(n591), .Z(G1355GAT) );
endmodule

