//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069;
  NOR2_X1   g000(.A1(G475), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT75), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT75), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G125), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n188), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  NOR2_X1   g007(.A1(G125), .A2(G140), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT16), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT16), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(new_n188), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n197), .B1(new_n190), .B2(new_n192), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n195), .A2(G146), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  XNOR2_X1  g015(.A(G125), .B(G140), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT19), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n194), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT75), .B(G125), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(new_n188), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n201), .B(new_n204), .C1(new_n207), .C2(new_n203), .ZN(new_n208));
  NOR2_X1   g022(.A1(G237), .A2(G953), .ZN(new_n209));
  AND3_X1   g023(.A1(new_n209), .A2(G143), .A3(G214), .ZN(new_n210));
  AOI21_X1  g024(.A(G143), .B1(new_n209), .B2(G214), .ZN(new_n211));
  OAI21_X1  g025(.A(G131), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G237), .ZN(new_n213));
  INV_X1    g027(.A(G953), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G214), .ZN(new_n215));
  INV_X1    g029(.A(G143), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G131), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n209), .A2(G143), .A3(G214), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n212), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n200), .A2(new_n208), .A3(new_n221), .ZN(new_n222));
  OAI211_X1 g036(.A(G146), .B(new_n205), .C1(new_n206), .C2(new_n188), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT91), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n202), .A2(new_n201), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n190), .A2(new_n192), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n194), .B1(new_n227), .B2(G140), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT91), .A3(G146), .ZN(new_n229));
  AND2_X1   g043(.A1(KEYINPUT90), .A2(KEYINPUT18), .ZN(new_n230));
  OAI211_X1 g044(.A(G131), .B(new_n230), .C1(new_n210), .C2(new_n211), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(G131), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n217), .A2(new_n219), .A3(new_n232), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n226), .A2(new_n229), .A3(new_n231), .A4(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n222), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G113), .B(G122), .ZN(new_n236));
  INV_X1    g050(.A(G104), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n236), .B(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n235), .A2(KEYINPUT92), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n195), .A2(new_n199), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n201), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n200), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT17), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n212), .A2(new_n244), .A3(new_n220), .ZN(new_n245));
  OAI211_X1 g059(.A(KEYINPUT17), .B(G131), .C1(new_n210), .C2(new_n211), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n238), .B(new_n234), .C1(new_n243), .C2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n240), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT92), .B1(new_n235), .B2(new_n239), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n187), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT20), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT20), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n253), .B(new_n187), .C1(new_n249), .C2(new_n250), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G475), .ZN(new_n256));
  AOI211_X1 g070(.A(new_n201), .B(new_n198), .C1(new_n207), .C2(KEYINPUT16), .ZN(new_n257));
  AOI21_X1  g071(.A(G146), .B1(new_n195), .B2(new_n199), .ZN(new_n258));
  NOR3_X1   g072(.A1(new_n247), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n234), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n239), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n248), .ZN(new_n262));
  INV_X1    g076(.A(G902), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n256), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT93), .B1(new_n255), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT93), .ZN(new_n267));
  AOI211_X1 g081(.A(new_n267), .B(new_n264), .C1(new_n252), .C2(new_n254), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  XOR2_X1   g083(.A(G116), .B(G122), .Z(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G107), .ZN(new_n271));
  XNOR2_X1  g085(.A(G116), .B(G122), .ZN(new_n272));
  INV_X1    g086(.A(G107), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT94), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n271), .A2(KEYINPUT94), .A3(new_n274), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G128), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT13), .B1(new_n280), .B2(G143), .ZN(new_n281));
  INV_X1    g095(.A(G134), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(G128), .B(G143), .ZN(new_n284));
  OR2_X1    g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n284), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n279), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G116), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT14), .A3(G122), .ZN(new_n290));
  OAI211_X1 g104(.A(G107), .B(new_n290), .C1(new_n270), .C2(KEYINPUT14), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n284), .A2(G134), .ZN(new_n292));
  OR2_X1    g106(.A1(new_n284), .A2(G134), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n291), .A2(new_n274), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT9), .B(G234), .ZN(new_n295));
  INV_X1    g109(.A(G217), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n295), .A2(new_n296), .A3(G953), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n288), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n297), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n277), .A2(new_n278), .B1(new_n285), .B2(new_n286), .ZN(new_n300));
  INV_X1    g114(.A(new_n294), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n263), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT15), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(G478), .ZN(new_n306));
  INV_X1    g120(.A(G478), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n303), .B(new_n263), .C1(KEYINPUT15), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n201), .A2(G143), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n216), .A2(G146), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AND2_X1   g127(.A1(KEYINPUT0), .A2(G128), .ZN(new_n314));
  NOR2_X1   g128(.A1(KEYINPUT0), .A2(G128), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(new_n313), .B2(new_n314), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n227), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n319));
  INV_X1    g133(.A(new_n311), .ZN(new_n320));
  OAI21_X1  g134(.A(G128), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n311), .A2(new_n312), .A3(G128), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n321), .A2(new_n313), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n318), .B1(new_n323), .B2(new_n227), .ZN(new_n324));
  INV_X1    g138(.A(G224), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n324), .B(KEYINPUT7), .C1(new_n325), .C2(G953), .ZN(new_n326));
  XNOR2_X1  g140(.A(G110), .B(G122), .ZN(new_n327));
  XOR2_X1   g141(.A(new_n327), .B(KEYINPUT8), .Z(new_n328));
  INV_X1    g142(.A(G119), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G116), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n289), .A2(G119), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT2), .B(G113), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT5), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G113), .ZN(new_n338));
  INV_X1    g152(.A(new_n330), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n338), .B1(new_n339), .B2(new_n335), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n334), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(KEYINPUT3), .B1(new_n237), .B2(G107), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT3), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(new_n273), .A3(G104), .ZN(new_n344));
  INV_X1    g158(.A(G101), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n237), .A2(G107), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n342), .A2(new_n344), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n273), .A2(G104), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n237), .A2(G107), .ZN(new_n349));
  OAI21_X1  g163(.A(G101), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n328), .B1(new_n341), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n340), .A2(KEYINPUT88), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n353), .A2(new_n336), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n340), .A2(KEYINPUT88), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n334), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n352), .B1(new_n356), .B2(new_n351), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT7), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n325), .A2(G953), .ZN(new_n359));
  OAI221_X1 g173(.A(new_n318), .B1(new_n358), .B2(new_n359), .C1(new_n323), .C2(new_n227), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n326), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n351), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n341), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n334), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT66), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n332), .A2(new_n333), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n332), .A2(new_n333), .A3(KEYINPUT66), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n342), .A2(new_n344), .A3(new_n346), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT82), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(G101), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(KEYINPUT4), .A3(new_n347), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n370), .A2(new_n371), .A3(new_n374), .A4(G101), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n327), .B(new_n363), .C1(new_n369), .C2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(G902), .B1(new_n361), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n363), .B1(new_n369), .B2(new_n376), .ZN(new_n379));
  INV_X1    g193(.A(new_n327), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(KEYINPUT6), .A3(new_n377), .ZN(new_n382));
  XOR2_X1   g196(.A(new_n324), .B(new_n359), .Z(new_n383));
  INV_X1    g197(.A(KEYINPUT6), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n379), .A2(new_n384), .A3(new_n380), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n378), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT89), .ZN(new_n388));
  OAI21_X1  g202(.A(G210), .B1(G237), .B2(G902), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n387), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n378), .B(new_n386), .C1(KEYINPUT89), .C2(new_n389), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(G234), .A2(G237), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n394), .A2(G952), .A3(new_n214), .ZN(new_n395));
  XOR2_X1   g209(.A(KEYINPUT21), .B(G898), .Z(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(KEYINPUT95), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n394), .A2(G902), .A3(G953), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n395), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(G214), .B1(G237), .B2(G902), .ZN(new_n401));
  XOR2_X1   g215(.A(new_n401), .B(KEYINPUT87), .Z(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n269), .A2(new_n310), .A3(new_n393), .A4(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G469), .ZN(new_n407));
  XNOR2_X1  g221(.A(G110), .B(G140), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n408), .B(KEYINPUT80), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n214), .A2(G227), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT11), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n413), .B1(new_n282), .B2(G137), .ZN(new_n414));
  INV_X1    g228(.A(G137), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(KEYINPUT11), .A3(G134), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n282), .A2(G137), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(G131), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n414), .A2(new_n416), .A3(new_n218), .A4(new_n417), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT83), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n423), .B(KEYINPUT1), .C1(new_n216), .C2(G146), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G128), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n423), .B1(new_n311), .B2(KEYINPUT1), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n313), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n322), .A2(new_n319), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n351), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT84), .B1(new_n429), .B2(KEYINPUT10), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT84), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT10), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT1), .B1(new_n216), .B2(G146), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT83), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(G128), .A3(new_n424), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n435), .A2(new_n313), .B1(new_n319), .B2(new_n322), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n431), .B(new_n432), .C1(new_n436), .C2(new_n351), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n430), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT67), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n311), .A2(new_n312), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT65), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(KEYINPUT1), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT1), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(KEYINPUT65), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n311), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n440), .B1(new_n445), .B2(G128), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n443), .A2(KEYINPUT65), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n441), .A2(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n313), .A2(new_n449), .A3(new_n280), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n439), .B1(new_n446), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n280), .B1(new_n449), .B2(new_n311), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n428), .B(KEYINPUT67), .C1(new_n452), .C2(new_n440), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n351), .A2(new_n432), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n373), .A2(new_n317), .A3(new_n375), .ZN(new_n456));
  AND4_X1   g270(.A1(new_n422), .A2(new_n438), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n455), .A2(new_n456), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n422), .B1(new_n458), .B2(new_n438), .ZN(new_n459));
  OAI211_X1 g273(.A(KEYINPUT86), .B(new_n412), .C1(new_n457), .C2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n428), .B1(new_n452), .B2(new_n440), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(new_n362), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n421), .B1(new_n462), .B2(new_n429), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT12), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(KEYINPUT12), .B(new_n421), .C1(new_n462), .C2(new_n429), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n438), .A2(new_n422), .A3(new_n455), .A4(new_n456), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n468), .A3(new_n411), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n460), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n430), .A2(new_n437), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n455), .A2(new_n456), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n421), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n468), .ZN(new_n474));
  AOI21_X1  g288(.A(KEYINPUT86), .B1(new_n474), .B2(new_n412), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n407), .B(new_n263), .C1(new_n470), .C2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n407), .A2(new_n263), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n468), .A2(new_n411), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT85), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n468), .A2(new_n481), .A3(new_n411), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n473), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n467), .A2(new_n468), .ZN(new_n484));
  XOR2_X1   g298(.A(new_n411), .B(KEYINPUT81), .Z(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(G469), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n476), .A2(new_n478), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(G221), .B1(new_n295), .B2(G902), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n406), .A2(KEYINPUT96), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n209), .A2(G210), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(KEYINPUT27), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT26), .B(G101), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT64), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n497), .B1(new_n282), .B2(G137), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n415), .A2(KEYINPUT64), .A3(G134), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n417), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G131), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n501), .A2(new_n420), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n502), .A2(new_n461), .B1(new_n421), .B2(new_n317), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT69), .B1(new_n503), .B2(new_n369), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n451), .A2(new_n502), .A3(new_n453), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n317), .A2(new_n421), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n506), .A3(new_n369), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n313), .A2(new_n314), .ZN(new_n508));
  OR2_X1    g322(.A1(new_n314), .A2(new_n315), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n508), .B1(new_n313), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n501), .A2(new_n420), .ZN(new_n511));
  OAI22_X1  g325(.A1(new_n422), .A2(new_n510), .B1(new_n323), .B2(new_n511), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n367), .A2(new_n368), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT69), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n504), .A2(new_n507), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT28), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT28), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n507), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n496), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n507), .A2(new_n496), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT30), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n369), .B1(new_n512), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n523), .B1(new_n317), .B2(new_n421), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n505), .A2(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n524), .A2(KEYINPUT68), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(KEYINPUT68), .B1(new_n524), .B2(new_n526), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n522), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT31), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT68), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n505), .A2(new_n525), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n513), .B1(new_n503), .B2(KEYINPUT30), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n524), .A2(KEYINPUT68), .A3(new_n526), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(KEYINPUT31), .A3(new_n522), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n520), .B1(new_n531), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(G472), .A2(G902), .ZN(new_n540));
  XOR2_X1   g354(.A(new_n540), .B(KEYINPUT70), .Z(new_n541));
  OAI21_X1  g355(.A(KEYINPUT32), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n517), .A2(new_n519), .ZN(new_n543));
  INV_X1    g357(.A(new_n496), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT31), .B1(new_n537), .B2(new_n522), .ZN(new_n546));
  AOI211_X1 g360(.A(new_n530), .B(new_n521), .C1(new_n535), .C2(new_n536), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT32), .ZN(new_n549));
  INV_X1    g363(.A(new_n541), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n505), .A2(new_n506), .A3(new_n369), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n369), .B1(new_n505), .B2(new_n506), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT28), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n496), .A2(KEYINPUT29), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(new_n507), .B2(new_n518), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(KEYINPUT71), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n263), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT71), .B1(new_n554), .B2(new_n556), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT72), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n554), .A2(new_n556), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT71), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT72), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n563), .A2(new_n564), .A3(new_n263), .A4(new_n557), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n517), .A2(new_n519), .A3(new_n496), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT29), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n552), .B1(new_n535), .B2(new_n536), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n566), .B(new_n567), .C1(new_n496), .C2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n560), .A2(new_n565), .A3(new_n569), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n542), .A2(new_n551), .B1(new_n570), .B2(G472), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT25), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n329), .A2(G128), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT73), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n574), .B1(new_n280), .B2(G119), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n329), .A2(KEYINPUT73), .A3(G128), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n573), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT24), .B(G110), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(G110), .ZN(new_n581));
  OR2_X1    g395(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n582));
  NAND2_X1  g396(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n573), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n280), .A2(G119), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n329), .A2(G128), .ZN(new_n586));
  AND2_X1   g400(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n580), .B1(new_n581), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n242), .B2(new_n200), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(G110), .B1(new_n584), .B2(new_n588), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT76), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n575), .A2(new_n576), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n585), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n593), .A2(new_n594), .B1(new_n596), .B2(new_n578), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n589), .A2(new_n581), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT76), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n225), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n198), .B1(new_n207), .B2(KEYINPUT16), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n601), .B1(new_n602), .B2(G146), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n600), .A2(KEYINPUT77), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT77), .B1(new_n600), .B2(new_n603), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n592), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n214), .A2(G221), .A3(G234), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT78), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT22), .B(G137), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT77), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n593), .A2(new_n594), .ZN(new_n614));
  AOI211_X1 g428(.A(KEYINPUT76), .B(G110), .C1(new_n584), .C2(new_n588), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n577), .A2(new_n579), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n200), .A2(new_n225), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n613), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n600), .A2(new_n603), .A3(KEYINPUT77), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n621), .A2(new_n592), .A3(new_n610), .ZN(new_n622));
  AOI21_X1  g436(.A(G902), .B1(new_n612), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT79), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n572), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n610), .B1(new_n621), .B2(new_n592), .ZN(new_n626));
  AOI211_X1 g440(.A(new_n591), .B(new_n611), .C1(new_n619), .C2(new_n620), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n263), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n628), .A2(KEYINPUT79), .A3(KEYINPUT25), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n296), .B1(G234), .B2(new_n263), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n625), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n612), .A2(new_n622), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n630), .A2(G902), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n571), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT96), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n637), .B1(new_n405), .B2(new_n490), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n492), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT97), .B(G101), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G3));
  INV_X1    g455(.A(new_n635), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n491), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n539), .A2(G902), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT98), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n548), .A2(new_n263), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT98), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n646), .A2(G472), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n548), .A2(new_n550), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(KEYINPUT99), .B1(new_n643), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n490), .A2(new_n635), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT99), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n653), .A2(new_n654), .A3(new_n650), .A4(new_n649), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n254), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n235), .A2(new_n239), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT92), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n248), .A3(new_n240), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n253), .B1(new_n662), .B2(new_n187), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n265), .B1(new_n658), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n267), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n255), .A2(KEYINPUT93), .A3(new_n265), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n307), .A2(G902), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT33), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n298), .A2(new_n302), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n669), .B1(new_n298), .B2(new_n302), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n668), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT100), .B(G478), .Z(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n303), .B2(new_n263), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n667), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n401), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n387), .A2(new_n390), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n378), .A2(new_n386), .A3(new_n389), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n400), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n657), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT34), .B(G104), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G6));
  NAND3_X1  g501(.A1(new_n252), .A2(KEYINPUT101), .A3(new_n254), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n688), .B1(KEYINPUT101), .B2(new_n254), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n264), .A2(KEYINPUT102), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT102), .ZN(new_n691));
  AOI21_X1  g505(.A(G902), .B1(new_n261), .B2(new_n248), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n691), .B1(new_n692), .B2(new_n256), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n309), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n683), .A2(new_n689), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n657), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT103), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT35), .B(G107), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G9));
  NOR2_X1   g513(.A1(new_n610), .A2(KEYINPUT36), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT104), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n606), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n633), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n631), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n651), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n638), .A3(new_n492), .ZN(new_n707));
  XOR2_X1   g521(.A(KEYINPUT37), .B(G110), .Z(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G12));
  NAND2_X1  g523(.A1(new_n570), .A2(G472), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n549), .B1(new_n548), .B2(new_n550), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n539), .A2(KEYINPUT32), .A3(new_n541), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n682), .A3(new_n704), .ZN(new_n714));
  INV_X1    g528(.A(G900), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n398), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n395), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n689), .A2(new_n694), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n489), .A3(new_n488), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT105), .B1(new_n714), .B2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n721), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n704), .A2(new_n682), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n571), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT105), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n723), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n722), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G128), .ZN(G30));
  XNOR2_X1  g543(.A(new_n718), .B(KEYINPUT39), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n491), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT40), .ZN(new_n732));
  OR2_X1    g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  INV_X1    g548(.A(new_n568), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n496), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n552), .A2(new_n553), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n736), .B(new_n263), .C1(new_n496), .C2(new_n737), .ZN(new_n738));
  AOI22_X1  g552(.A1(new_n542), .A2(new_n551), .B1(G472), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n704), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT38), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n393), .B(new_n741), .ZN(new_n742));
  NOR4_X1   g556(.A1(new_n742), .A2(new_n269), .A3(new_n310), .A4(new_n679), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n733), .A2(new_n734), .A3(new_n740), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G143), .ZN(G45));
  NAND3_X1  g559(.A1(new_n667), .A2(new_n677), .A3(new_n718), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n490), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n725), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G146), .ZN(G48));
  INV_X1    g563(.A(new_n636), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n263), .B1(new_n470), .B2(new_n475), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT106), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI211_X1 g567(.A(KEYINPUT106), .B(new_n263), .C1(new_n470), .C2(new_n475), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(G469), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n476), .A2(new_n489), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n750), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n684), .ZN(new_n760));
  XNOR2_X1  g574(.A(KEYINPUT41), .B(G113), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(KEYINPUT107), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n760), .B(new_n762), .ZN(G15));
  NAND2_X1  g577(.A1(new_n759), .A2(new_n695), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G116), .ZN(G18));
  AOI21_X1  g579(.A(new_n407), .B1(new_n751), .B2(new_n752), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n756), .B1(new_n766), .B2(new_n754), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n667), .A2(new_n309), .A3(new_n399), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n725), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G119), .ZN(G21));
  AND2_X1   g584(.A1(new_n554), .A2(new_n519), .ZN(new_n771));
  OAI22_X1  g585(.A1(new_n546), .A2(new_n547), .B1(new_n496), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n550), .ZN(new_n773));
  INV_X1    g587(.A(G472), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n773), .B1(new_n644), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n635), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n776), .A2(new_n400), .A3(new_n767), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n680), .A2(new_n681), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n310), .A2(new_n679), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n778), .B(new_n779), .C1(new_n266), .C2(new_n268), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT108), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n667), .A2(KEYINPUT108), .A3(new_n778), .A4(new_n779), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n777), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G122), .ZN(G24));
  AND3_X1   g600(.A1(new_n755), .A2(new_n682), .A3(new_n757), .ZN(new_n787));
  INV_X1    g601(.A(new_n746), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n647), .A2(G472), .ZN(new_n790));
  AND4_X1   g604(.A1(new_n789), .A2(new_n790), .A3(new_n704), .A4(new_n773), .ZN(new_n791));
  AOI22_X1  g605(.A1(new_n647), .A2(G472), .B1(new_n550), .B2(new_n772), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n789), .B1(new_n792), .B2(new_n704), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n787), .B(new_n788), .C1(new_n791), .C2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G125), .ZN(G27));
  INV_X1    g609(.A(new_n489), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n391), .A2(new_n392), .A3(new_n401), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT110), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n486), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n484), .A2(KEYINPUT110), .A3(new_n485), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n483), .A2(new_n799), .A3(G469), .A4(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n801), .A2(new_n478), .ZN(new_n802));
  AOI211_X1 g616(.A(new_n796), .B(new_n797), .C1(new_n802), .C2(new_n476), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n636), .A2(new_n788), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT42), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n636), .A2(new_n803), .A3(KEYINPUT42), .A4(new_n788), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G131), .ZN(G33));
  NAND3_X1  g623(.A1(new_n636), .A2(new_n720), .A3(new_n803), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G134), .ZN(G36));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n483), .A2(new_n799), .A3(KEYINPUT45), .A4(new_n800), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n483), .A2(new_n486), .ZN(new_n814));
  OAI211_X1 g628(.A(G469), .B(new_n813), .C1(new_n814), .C2(KEYINPUT45), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n478), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT46), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n812), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n815), .A2(KEYINPUT111), .A3(KEYINPUT46), .A4(new_n478), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n476), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n816), .A2(new_n817), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n820), .B(new_n824), .C1(new_n823), .C2(new_n822), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n489), .A3(new_n730), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT113), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n269), .A2(KEYINPUT43), .A3(new_n677), .ZN(new_n828));
  INV_X1    g642(.A(new_n677), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n677), .A2(KEYINPUT114), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n665), .A2(new_n831), .A3(new_n666), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT43), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n833), .A2(KEYINPUT115), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT115), .B1(new_n833), .B2(new_n834), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n828), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n833), .A2(new_n834), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n833), .A2(KEYINPUT115), .A3(new_n834), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(KEYINPUT116), .A3(new_n828), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n651), .A2(new_n839), .A3(new_n845), .A4(new_n704), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n797), .B1(new_n846), .B2(KEYINPUT44), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n827), .B(new_n847), .C1(KEYINPUT44), .C2(new_n846), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(G137), .ZN(G39));
  NAND2_X1  g663(.A1(new_n825), .A2(new_n489), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT47), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n825), .A2(KEYINPUT47), .A3(new_n489), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n713), .A2(new_n642), .A3(new_n797), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n788), .A3(new_n855), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(G140), .ZN(G42));
  INV_X1    g671(.A(G952), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n214), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT52), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n726), .B1(new_n723), .B2(new_n725), .ZN(new_n861));
  NOR4_X1   g675(.A1(new_n721), .A2(new_n571), .A3(new_n724), .A4(KEYINPUT105), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n794), .A2(new_n748), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n782), .A2(new_n783), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n738), .A2(G472), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n868), .B1(new_n712), .B2(new_n711), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n802), .A2(new_n476), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n719), .A2(new_n796), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n869), .A2(new_n705), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n866), .B1(new_n867), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n870), .A2(new_n871), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n784), .A2(new_n874), .A3(new_n740), .A4(KEYINPUT118), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n860), .B1(new_n865), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT109), .B1(new_n775), .B2(new_n705), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n792), .A2(new_n789), .A3(new_n704), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n746), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n880), .A2(new_n787), .B1(new_n725), .B2(new_n747), .ZN(new_n881));
  AND4_X1   g695(.A1(new_n860), .A2(new_n876), .A3(new_n881), .A4(new_n728), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT119), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n725), .A2(new_n768), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n767), .A2(new_n884), .B1(new_n777), .B2(new_n784), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n393), .A2(new_n404), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n667), .A2(new_n310), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT117), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n887), .A2(new_n888), .B1(new_n667), .B2(new_n677), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT117), .B1(new_n667), .B2(new_n310), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n652), .A2(new_n891), .A3(new_n655), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n638), .B(new_n492), .C1(new_n706), .C2(new_n636), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n636), .B(new_n767), .C1(new_n684), .C2(new_n695), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n885), .A2(new_n892), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n810), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n896), .B1(new_n806), .B2(new_n807), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n310), .A2(new_n693), .A3(new_n690), .A4(new_n718), .ZN(new_n898));
  OR3_X1    g712(.A1(new_n797), .A2(new_n898), .A3(new_n689), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n899), .A2(new_n571), .A3(new_n705), .ZN(new_n900));
  AOI22_X1  g714(.A1(new_n880), .A2(new_n803), .B1(new_n900), .B2(new_n491), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n873), .A2(new_n875), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n794), .B(new_n748), .C1(new_n861), .C2(new_n862), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT52), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT119), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n876), .A2(new_n881), .A3(new_n728), .A4(new_n860), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n883), .A2(KEYINPUT53), .A3(new_n903), .A4(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT53), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n785), .A2(new_n894), .A3(new_n769), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n707), .A2(new_n639), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n914), .A2(new_n892), .A3(new_n897), .A4(new_n901), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n906), .A2(new_n908), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n911), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n910), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT54), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n903), .A2(KEYINPUT53), .A3(new_n908), .A4(new_n906), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n907), .B1(new_n906), .B2(new_n908), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n922), .A2(new_n923), .A3(new_n915), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n920), .B(new_n921), .C1(new_n924), .C2(KEYINPUT53), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n758), .A2(new_n797), .ZN(new_n926));
  AND4_X1   g740(.A1(new_n642), .A2(new_n926), .A3(new_n395), .A4(new_n739), .ZN(new_n927));
  INV_X1    g741(.A(new_n678), .ZN(new_n928));
  AOI211_X1 g742(.A(new_n858), .B(G953), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n787), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n837), .A2(new_n395), .A3(new_n776), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n717), .B1(new_n844), .B2(new_n828), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(new_n636), .A3(new_n926), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n933), .A2(KEYINPUT48), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n933), .A2(KEYINPUT48), .ZN(new_n935));
  OAI221_X1 g749(.A(new_n929), .B1(new_n930), .B2(new_n931), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n932), .B(new_n926), .C1(new_n791), .C2(new_n793), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n927), .A2(new_n269), .A3(new_n829), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(KEYINPUT51), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT50), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n942), .B1(new_n758), .B2(new_n401), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n755), .A2(new_n757), .A3(KEYINPUT121), .A4(new_n679), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n943), .A2(new_n742), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n941), .B1(new_n931), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n944), .A2(new_n742), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT121), .B1(new_n767), .B2(new_n679), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n932), .A2(KEYINPUT50), .A3(new_n949), .A4(new_n776), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n940), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n931), .A2(new_n797), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n755), .A2(new_n476), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n953), .A2(new_n489), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n952), .B1(new_n854), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n936), .B1(new_n951), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n919), .A2(new_n925), .A3(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT123), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n946), .A2(new_n950), .A3(KEYINPUT122), .ZN(new_n959));
  AOI21_X1  g773(.A(KEYINPUT122), .B1(new_n946), .B2(new_n950), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n939), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n853), .ZN(new_n962));
  AOI21_X1  g776(.A(KEYINPUT47), .B1(new_n825), .B2(new_n489), .ZN(new_n963));
  OAI21_X1  g777(.A(KEYINPUT120), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT120), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n852), .A2(new_n965), .A3(new_n853), .ZN(new_n966));
  INV_X1    g780(.A(new_n954), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n961), .B1(new_n968), .B2(new_n952), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n958), .B1(new_n969), .B2(KEYINPUT51), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT51), .ZN(new_n971));
  INV_X1    g785(.A(new_n952), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n954), .B1(new_n854), .B2(KEYINPUT120), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n972), .B1(new_n973), .B2(new_n966), .ZN(new_n974));
  OAI211_X1 g788(.A(KEYINPUT123), .B(new_n971), .C1(new_n974), .C2(new_n961), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n970), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n859), .B1(new_n957), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n742), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n642), .A2(new_n489), .A3(new_n402), .A4(new_n677), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n978), .A2(new_n979), .A3(new_n667), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n953), .A2(KEYINPUT49), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n953), .A2(KEYINPUT49), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n980), .A2(new_n739), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n977), .A2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT124), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n977), .A2(KEYINPUT124), .A3(new_n983), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(G75));
  NAND3_X1  g802(.A1(new_n883), .A2(new_n903), .A3(new_n909), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n911), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n921), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n991), .A2(G210), .A3(G902), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT56), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n382), .A2(new_n385), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(new_n383), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT55), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n992), .A2(new_n993), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n996), .B1(new_n992), .B2(new_n993), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n214), .A2(G952), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(G51));
  NAND2_X1  g814(.A1(new_n991), .A2(KEYINPUT54), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n925), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n477), .B(KEYINPUT57), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1004), .B1(new_n475), .B2(new_n470), .ZN(new_n1005));
  AND2_X1   g819(.A1(new_n990), .A2(new_n921), .ZN(new_n1006));
  OR3_X1    g820(.A1(new_n1006), .A2(new_n263), .A3(new_n815), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n999), .B1(new_n1005), .B2(new_n1007), .ZN(G54));
  NOR2_X1   g822(.A1(new_n1006), .A2(new_n263), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1009), .A2(KEYINPUT58), .A3(G475), .ZN(new_n1010));
  INV_X1    g824(.A(new_n662), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n999), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1009), .A2(KEYINPUT58), .A3(G475), .A4(new_n662), .ZN(new_n1014));
  AND3_X1   g828(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(G60));
  NOR2_X1   g829(.A1(new_n671), .A2(new_n672), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n919), .A2(new_n925), .ZN(new_n1018));
  XNOR2_X1  g832(.A(KEYINPUT125), .B(KEYINPUT59), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n307), .A2(new_n263), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1017), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  AND2_X1   g836(.A1(new_n1017), .A2(new_n1021), .ZN(new_n1023));
  AOI211_X1 g837(.A(new_n999), .B(new_n1022), .C1(new_n1002), .C2(new_n1023), .ZN(G63));
  NAND2_X1  g838(.A1(G217), .A2(G902), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1025), .B(KEYINPUT60), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1026), .B1(new_n990), .B2(new_n921), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n999), .B1(new_n1027), .B2(new_n702), .ZN(new_n1028));
  INV_X1    g842(.A(KEYINPUT61), .ZN(new_n1029));
  OAI221_X1 g843(.A(new_n1028), .B1(KEYINPUT126), .B2(new_n1029), .C1(new_n632), .C2(new_n1027), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1026), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n991), .A2(new_n702), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1032), .A2(KEYINPUT126), .A3(new_n1013), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1032), .A2(new_n1013), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n1027), .A2(new_n632), .ZN(new_n1035));
  OAI211_X1 g849(.A(new_n1033), .B(KEYINPUT61), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  AND2_X1   g850(.A1(new_n1030), .A2(new_n1036), .ZN(G66));
  OAI21_X1  g851(.A(G953), .B1(new_n397), .B2(new_n325), .ZN(new_n1038));
  INV_X1    g852(.A(new_n895), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1038), .B1(new_n1039), .B2(G953), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n994), .B1(G898), .B2(new_n214), .ZN(new_n1041));
  XOR2_X1   g855(.A(new_n1041), .B(KEYINPUT127), .Z(new_n1042));
  XNOR2_X1  g856(.A(new_n1040), .B(new_n1042), .ZN(G69));
  NAND2_X1  g857(.A1(new_n865), .A2(new_n897), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n750), .A2(new_n867), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n1044), .B1(new_n827), .B2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g860(.A1(new_n848), .A2(new_n1046), .A3(new_n214), .A4(new_n856), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n526), .B1(KEYINPUT30), .B2(new_n503), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n204), .B1(new_n207), .B2(new_n203), .ZN(new_n1049));
  XNOR2_X1  g863(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  OAI211_X1 g864(.A(new_n1047), .B(new_n1050), .C1(new_n715), .C2(new_n214), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n865), .A2(new_n744), .ZN(new_n1052));
  XOR2_X1   g866(.A(new_n1052), .B(KEYINPUT62), .Z(new_n1053));
  NOR2_X1   g867(.A1(new_n750), .A2(new_n797), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n889), .A2(new_n890), .ZN(new_n1055));
  NAND3_X1  g869(.A1(new_n1054), .A2(new_n1055), .A3(new_n731), .ZN(new_n1056));
  NAND4_X1  g870(.A1(new_n1053), .A2(new_n848), .A3(new_n856), .A4(new_n1056), .ZN(new_n1057));
  AND2_X1   g871(.A1(new_n1057), .A2(new_n214), .ZN(new_n1058));
  OAI21_X1  g872(.A(new_n1051), .B1(new_n1058), .B2(new_n1050), .ZN(new_n1059));
  AOI21_X1  g873(.A(new_n214), .B1(G227), .B2(G900), .ZN(new_n1060));
  XNOR2_X1  g874(.A(new_n1059), .B(new_n1060), .ZN(G72));
  OR2_X1    g875(.A1(new_n1057), .A2(new_n895), .ZN(new_n1062));
  NAND2_X1  g876(.A1(G472), .A2(G902), .ZN(new_n1063));
  XOR2_X1   g877(.A(new_n1063), .B(KEYINPUT63), .Z(new_n1064));
  AOI21_X1  g878(.A(new_n736), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g879(.A1(new_n848), .A2(new_n1046), .A3(new_n856), .A4(new_n1039), .ZN(new_n1066));
  AOI211_X1 g880(.A(new_n496), .B(new_n735), .C1(new_n1066), .C2(new_n1064), .ZN(new_n1067));
  OAI21_X1  g881(.A(new_n529), .B1(new_n568), .B2(new_n496), .ZN(new_n1068));
  AND3_X1   g882(.A1(new_n918), .A2(new_n1064), .A3(new_n1068), .ZN(new_n1069));
  NOR4_X1   g883(.A1(new_n1065), .A2(new_n999), .A3(new_n1067), .A4(new_n1069), .ZN(G57));
endmodule


