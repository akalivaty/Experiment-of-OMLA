//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT65), .Z(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT23), .ZN(new_n207));
  OR2_X1    g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209));
  AND3_X1   g008(.A1(new_n208), .A2(KEYINPUT24), .A3(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n205), .A2(KEYINPUT23), .ZN(new_n211));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(new_n209), .B2(KEYINPUT24), .ZN(new_n213));
  NOR3_X1   g012(.A1(new_n210), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n207), .A2(new_n214), .A3(KEYINPUT25), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n205), .A2(KEYINPUT23), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n215), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT27), .B(G183gat), .ZN(new_n220));
  INV_X1    g019(.A(G190gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(KEYINPUT28), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n220), .A2(KEYINPUT66), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT27), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT66), .B1(new_n224), .B2(G183gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(new_n221), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n222), .B1(new_n227), .B2(KEYINPUT28), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT26), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n206), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n212), .B1(new_n205), .B2(new_n229), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n228), .B(new_n209), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n219), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G226gat), .A2(G233gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(KEYINPUT72), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n233), .B1(KEYINPUT29), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G211gat), .A2(G218gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT22), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(KEYINPUT70), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G197gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G204gat), .ZN(new_n241));
  INV_X1    g040(.A(G204gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G197gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n239), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT70), .B1(new_n237), .B2(new_n238), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(G211gat), .B(G218gat), .Z(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT71), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(new_n244), .B2(new_n245), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n248), .A2(new_n249), .B1(new_n247), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n235), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n219), .A2(new_n232), .A3(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n252), .B1(new_n236), .B2(new_n254), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n204), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n257), .ZN(new_n259));
  INV_X1    g058(.A(new_n204), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n255), .A3(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(new_n261), .A3(KEYINPUT30), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT30), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n263), .B(new_n204), .C1(new_n256), .C2(new_n257), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G1gat), .B(G29gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT0), .ZN(new_n268));
  XNOR2_X1  g067(.A(G57gat), .B(G85gat), .ZN(new_n269));
  XOR2_X1   g068(.A(new_n268), .B(new_n269), .Z(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G225gat), .A2(G233gat), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n272), .B(KEYINPUT75), .Z(new_n273));
  XOR2_X1   g072(.A(G141gat), .B(G148gat), .Z(new_n274));
  INV_X1    g073(.A(G155gat), .ZN(new_n275));
  INV_X1    g074(.A(G162gat), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT2), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G155gat), .B(G162gat), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n274), .A2(new_n277), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n279), .B(KEYINPUT73), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n280), .B(KEYINPUT74), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  OR3_X1    g082(.A1(new_n282), .A2(KEYINPUT74), .A3(new_n281), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G127gat), .B(G134gat), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n286), .B1(KEYINPUT67), .B2(KEYINPUT1), .ZN(new_n287));
  XNOR2_X1  g086(.A(G113gat), .B(G120gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(KEYINPUT1), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n287), .B(new_n289), .Z(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n290), .B1(new_n283), .B2(new_n284), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n273), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT5), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT4), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT76), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n293), .A2(new_n296), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n293), .A2(KEYINPUT76), .A3(new_n296), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT3), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n290), .B1(new_n285), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT3), .B1(new_n283), .B2(new_n284), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n273), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n295), .B1(new_n303), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT5), .ZN(new_n311));
  INV_X1    g110(.A(new_n273), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n311), .B(new_n312), .C1(new_n305), .C2(new_n307), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT77), .ZN(new_n314));
  INV_X1    g113(.A(new_n297), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n314), .B1(new_n315), .B2(new_n300), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n301), .A2(KEYINPUT77), .A3(new_n297), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n313), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n271), .B1(new_n310), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT84), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g120(.A(KEYINPUT84), .B(new_n271), .C1(new_n310), .C2(new_n318), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n266), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n316), .A2(new_n317), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n306), .A2(new_n308), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n312), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT39), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n271), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n292), .A2(new_n293), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n327), .B1(new_n329), .B2(new_n312), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n316), .A2(new_n317), .B1(new_n308), .B2(new_n306), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n330), .B1(new_n331), .B2(new_n312), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT40), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n326), .A2(new_n327), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n336), .A2(KEYINPUT40), .A3(new_n332), .A4(new_n270), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT85), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT85), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n328), .A2(new_n339), .A3(KEYINPUT40), .A4(new_n332), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n323), .A2(new_n335), .A3(new_n338), .A4(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT37), .B1(new_n256), .B2(new_n257), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT37), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n259), .A2(new_n343), .A3(new_n255), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n204), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT38), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n258), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n347), .B1(new_n346), .B2(new_n345), .ZN(new_n348));
  XOR2_X1   g147(.A(KEYINPUT78), .B(KEYINPUT6), .Z(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n271), .B(new_n350), .C1(new_n310), .C2(new_n318), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n303), .A2(new_n309), .ZN(new_n352));
  INV_X1    g151(.A(new_n295), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n313), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n324), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n354), .A2(new_n356), .A3(new_n270), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n321), .A2(new_n357), .A3(new_n349), .A4(new_n322), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n348), .A2(new_n351), .A3(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G78gat), .B(G106gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(KEYINPUT80), .B(G50gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  XOR2_X1   g161(.A(KEYINPUT79), .B(KEYINPUT31), .Z(new_n363));
  XOR2_X1   g162(.A(new_n362), .B(new_n363), .Z(new_n364));
  INV_X1    g163(.A(G22gat), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n252), .B1(new_n307), .B2(KEYINPUT29), .ZN(new_n366));
  INV_X1    g165(.A(new_n285), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n304), .B1(new_n252), .B2(KEYINPUT29), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G228gat), .A2(G233gat), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n366), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT82), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n366), .A2(new_n369), .A3(new_n374), .A4(new_n371), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n366), .A2(KEYINPUT81), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n378), .B(new_n252), .C1(new_n307), .C2(KEYINPUT29), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n246), .A2(new_n247), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n380), .A2(new_n248), .A3(KEYINPUT29), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n367), .B1(KEYINPUT3), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n377), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n370), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n365), .B1(new_n376), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT83), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n364), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n376), .A2(new_n384), .A3(new_n365), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n387), .B1(new_n385), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n385), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n391), .A2(new_n388), .A3(new_n386), .A4(new_n364), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n341), .A2(new_n359), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n357), .A2(new_n319), .A3(new_n349), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n351), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n390), .A2(new_n392), .B1(new_n396), .B2(new_n265), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT36), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT69), .ZN(new_n399));
  OR2_X1    g198(.A1(new_n398), .A2(KEYINPUT69), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n290), .B1(new_n219), .B2(new_n232), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(G227gat), .A2(G233gat), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n219), .A2(new_n232), .A3(new_n290), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n406), .A2(KEYINPUT32), .ZN(new_n407));
  XNOR2_X1  g206(.A(G15gat), .B(G43gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(G71gat), .B(G99gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT33), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n410), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT34), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n413), .B1(new_n403), .B2(KEYINPUT68), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n402), .A2(new_n405), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n415), .B1(new_n416), .B2(new_n403), .ZN(new_n417));
  AOI211_X1 g216(.A(new_n404), .B(new_n414), .C1(new_n402), .C2(new_n405), .ZN(new_n418));
  NOR3_X1   g217(.A1(new_n412), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n412), .B1(new_n417), .B2(new_n418), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n407), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n421), .ZN(new_n423));
  INV_X1    g222(.A(new_n407), .ZN(new_n424));
  NOR3_X1   g223(.A1(new_n423), .A2(new_n419), .A3(new_n424), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n399), .B(new_n400), .C1(new_n422), .C2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n420), .A2(new_n407), .A3(new_n421), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n424), .B1(new_n423), .B2(new_n419), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n427), .A2(new_n428), .A3(KEYINPUT69), .A4(new_n398), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n397), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT35), .B1(new_n358), .B2(new_n351), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n422), .A2(new_n425), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n393), .A2(new_n432), .A3(new_n265), .A4(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n266), .B1(new_n395), .B2(new_n351), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n435), .A2(new_n390), .A3(new_n433), .A4(new_n392), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT35), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n394), .A2(new_n431), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(G15gat), .B(G22gat), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT16), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n439), .B1(new_n440), .B2(G1gat), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(KEYINPUT89), .A3(G8gat), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n439), .A2(G1gat), .ZN(new_n443));
  OR2_X1    g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(G8gat), .B1(new_n441), .B2(KEYINPUT90), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n445), .B1(KEYINPUT90), .B2(new_n441), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT89), .ZN(new_n447));
  INV_X1    g246(.A(G8gat), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n443), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n444), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(G50gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(G43gat), .ZN(new_n452));
  INV_X1    g251(.A(G43gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(G50gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT15), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT87), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT87), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n452), .A2(new_n454), .A3(new_n458), .A4(KEYINPUT15), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n455), .A2(new_n456), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT14), .ZN(new_n462));
  INV_X1    g261(.A(G29gat), .ZN(new_n463));
  INV_X1    g262(.A(G36gat), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n465), .A2(new_n466), .B1(G29gat), .B2(G36gat), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(KEYINPUT86), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n465), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n466), .A2(KEYINPUT86), .ZN(new_n471));
  OAI22_X1  g270(.A1(new_n470), .A2(new_n471), .B1(new_n463), .B2(new_n464), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n455), .A2(new_n456), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n460), .A2(new_n468), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n450), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(new_n473), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n457), .A2(new_n461), .A3(new_n459), .A4(new_n467), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT17), .ZN(new_n478));
  XOR2_X1   g277(.A(KEYINPUT88), .B(KEYINPUT17), .Z(new_n479));
  OAI211_X1 g278(.A(new_n450), .B(new_n478), .C1(new_n474), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(G229gat), .A2(G233gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n475), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT18), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n450), .B(new_n474), .ZN(new_n484));
  XOR2_X1   g283(.A(new_n481), .B(KEYINPUT13), .Z(new_n485));
  AOI22_X1  g284(.A1(new_n482), .A2(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(G113gat), .B(G141gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(G197gat), .ZN(new_n488));
  XOR2_X1   g287(.A(KEYINPUT11), .B(G169gat), .Z(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(KEYINPUT12), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n475), .A2(new_n480), .A3(KEYINPUT18), .A4(new_n481), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n486), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n491), .B1(new_n486), .B2(new_n492), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT91), .B1(new_n438), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n394), .A2(new_n431), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n434), .A2(new_n437), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT91), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n493), .A2(new_n494), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  XOR2_X1   g302(.A(G134gat), .B(G162gat), .Z(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  AND2_X1   g304(.A1(G232gat), .A2(G233gat), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n506), .A2(KEYINPUT41), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT96), .ZN(new_n509));
  NAND2_X1  g308(.A1(G85gat), .A2(G92gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT95), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT95), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n512), .A2(G85gat), .A3(G92gat), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n513), .A3(KEYINPUT7), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT7), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n510), .A2(KEYINPUT95), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(G99gat), .A2(G106gat), .ZN(new_n517));
  INV_X1    g316(.A(G85gat), .ZN(new_n518));
  INV_X1    g317(.A(G92gat), .ZN(new_n519));
  AOI22_X1  g318(.A1(KEYINPUT8), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n514), .A2(new_n516), .A3(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G99gat), .B(G106gat), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n514), .A2(new_n522), .A3(new_n516), .A4(new_n520), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n478), .B(new_n526), .C1(new_n474), .C2(new_n479), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n476), .A2(new_n477), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n517), .A2(KEYINPUT8), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n518), .A2(new_n519), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n516), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n522), .B1(new_n531), .B2(new_n514), .ZN(new_n532));
  AND4_X1   g331(.A1(new_n522), .A2(new_n514), .A3(new_n516), .A4(new_n520), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n528), .A2(new_n534), .B1(KEYINPUT41), .B2(new_n506), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n527), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G190gat), .B(G218gat), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n509), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n537), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n527), .A2(KEYINPUT96), .A3(new_n535), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n539), .B1(new_n527), .B2(new_n535), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n542), .A2(KEYINPUT97), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(KEYINPUT97), .ZN(new_n544));
  AND4_X1   g343(.A1(new_n508), .A2(new_n541), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT97), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n542), .B(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n508), .B1(new_n547), .B2(new_n541), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n505), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n507), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n547), .A2(new_n508), .A3(new_n541), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(new_n504), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G71gat), .A2(G78gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OR2_X1    g356(.A1(G57gat), .A2(G64gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(G57gat), .A2(G64gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI22_X1  g359(.A1(KEYINPUT92), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n561));
  OR2_X1    g360(.A1(G71gat), .A2(G78gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n560), .B(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n564), .A2(KEYINPUT21), .ZN(new_n565));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n565), .B(new_n566), .Z(new_n567));
  XNOR2_X1  g366(.A(G127gat), .B(G155gat), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n568), .B(KEYINPUT93), .Z(new_n569));
  XNOR2_X1  g368(.A(new_n567), .B(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT94), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n564), .A2(KEYINPUT21), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n571), .B1(new_n450), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n450), .A2(new_n571), .A3(new_n572), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n570), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n577));
  XNOR2_X1  g376(.A(G183gat), .B(G211gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n569), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n567), .B(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n575), .A2(new_n573), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n576), .A2(new_n579), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n579), .B1(new_n576), .B2(new_n583), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n554), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT98), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n554), .A2(KEYINPUT98), .A3(new_n586), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n534), .A2(KEYINPUT10), .A3(new_n564), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT100), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT99), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n525), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n564), .B(new_n595), .C1(new_n532), .C2(new_n533), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n560), .A2(new_n562), .A3(new_n561), .ZN(new_n597));
  AND2_X1   g396(.A1(G57gat), .A2(G64gat), .ZN(new_n598));
  NOR2_X1   g397(.A1(G57gat), .A2(G64gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n563), .A2(new_n557), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n525), .B(new_n524), .C1(new_n602), .C2(new_n594), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n596), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT10), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n593), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI211_X1 g405(.A(KEYINPUT100), .B(KEYINPUT10), .C1(new_n596), .C2(new_n603), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n592), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G230gat), .A2(G233gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n610), .B1(new_n609), .B2(new_n604), .ZN(new_n611));
  XNOR2_X1  g410(.A(G120gat), .B(G148gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT101), .ZN(new_n613));
  XNOR2_X1  g412(.A(G176gat), .B(G204gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n611), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n591), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n503), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n396), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g423(.A(KEYINPUT16), .B(G8gat), .Z(new_n625));
  NAND3_X1  g424(.A1(new_n621), .A2(new_n266), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n448), .B1(new_n621), .B2(new_n266), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT42), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n629), .B1(KEYINPUT42), .B2(new_n627), .ZN(G1325gat));
  INV_X1    g429(.A(new_n430), .ZN(new_n631));
  OAI21_X1  g430(.A(G15gat), .B1(new_n620), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(G15gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n433), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n632), .B1(new_n620), .B2(new_n634), .ZN(G1326gat));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n393), .ZN(new_n636));
  XOR2_X1   g435(.A(KEYINPUT43), .B(G22gat), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(G1327gat));
  INV_X1    g437(.A(KEYINPUT44), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n639), .B1(new_n438), .B2(new_n554), .ZN(new_n640));
  INV_X1    g439(.A(new_n554), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n499), .A2(KEYINPUT44), .A3(new_n641), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n586), .A2(new_n618), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n501), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT103), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(G29gat), .B1(new_n647), .B2(new_n396), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n644), .A2(new_n641), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n649), .B1(new_n496), .B2(new_n502), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n650), .A2(new_n463), .A3(new_n622), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(KEYINPUT102), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT45), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n650), .A2(new_n654), .A3(new_n463), .A4(new_n622), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n653), .B1(new_n652), .B2(new_n655), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n648), .B1(new_n656), .B2(new_n657), .ZN(G1328gat));
  NAND3_X1  g457(.A1(new_n650), .A2(new_n464), .A3(new_n266), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n659), .A2(KEYINPUT46), .ZN(new_n660));
  OAI21_X1  g459(.A(G36gat), .B1(new_n647), .B2(new_n265), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(KEYINPUT46), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(G1329gat));
  OAI21_X1  g462(.A(G43gat), .B1(new_n647), .B2(new_n631), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n650), .A2(new_n453), .A3(new_n433), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT47), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1330gat));
  INV_X1    g467(.A(KEYINPUT48), .ZN(new_n669));
  INV_X1    g468(.A(new_n393), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n640), .A2(new_n642), .A3(new_n670), .A4(new_n646), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n671), .A2(G50gat), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n393), .A2(G50gat), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n650), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n669), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n451), .B1(new_n671), .B2(new_n676), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n669), .B1(new_n650), .B2(new_n673), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n680), .B1(new_n679), .B2(new_n681), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n675), .B1(new_n682), .B2(new_n683), .ZN(G1331gat));
  INV_X1    g483(.A(new_n618), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n591), .A2(new_n501), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n499), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(new_n622), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g489(.A1(new_n687), .A2(new_n265), .ZN(new_n691));
  NOR2_X1   g490(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n692));
  AND2_X1   g491(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(new_n691), .B2(new_n692), .ZN(G1333gat));
  OAI21_X1  g494(.A(G71gat), .B1(new_n687), .B2(new_n631), .ZN(new_n696));
  INV_X1    g495(.A(G71gat), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n433), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n696), .B1(new_n687), .B2(new_n698), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g499(.A1(new_n688), .A2(new_n670), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g501(.A(new_n554), .B1(new_n497), .B2(new_n498), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n586), .A2(new_n501), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT51), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n703), .A2(KEYINPUT51), .A3(new_n704), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n685), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n709), .A2(new_n518), .A3(new_n622), .ZN(new_n710));
  INV_X1    g509(.A(new_n704), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n685), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n643), .A2(new_n622), .A3(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(G85gat), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n713), .A2(new_n714), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n710), .B1(new_n716), .B2(new_n717), .ZN(G1336gat));
  NOR2_X1   g517(.A1(new_n265), .A2(G92gat), .ZN(new_n719));
  NOR4_X1   g518(.A1(new_n438), .A2(new_n706), .A3(new_n554), .A4(new_n711), .ZN(new_n720));
  AOI21_X1  g519(.A(KEYINPUT51), .B1(new_n703), .B2(new_n704), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n618), .B(new_n719), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(KEYINPUT107), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT52), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n640), .A2(new_n642), .A3(new_n266), .A4(new_n712), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(G92gat), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n722), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n727), .B1(new_n722), .B2(new_n726), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n724), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n722), .A2(new_n726), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT108), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n733), .B1(new_n722), .B2(KEYINPUT107), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n722), .A2(new_n726), .A3(new_n727), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n732), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n730), .A2(new_n736), .ZN(G1337gat));
  INV_X1    g536(.A(G99gat), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n709), .A2(new_n738), .A3(new_n433), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n643), .A2(new_n430), .A3(new_n712), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n738), .B2(new_n740), .ZN(G1338gat));
  NOR2_X1   g540(.A1(new_n393), .A2(G106gat), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n709), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n640), .A2(new_n642), .A3(new_n670), .A4(new_n712), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n744), .A2(G106gat), .ZN(new_n745));
  OAI21_X1  g544(.A(KEYINPUT53), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n747));
  OR2_X1    g546(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(G106gat), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n744), .B2(new_n747), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT53), .B1(new_n709), .B2(new_n742), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n751), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n753), .B1(new_n751), .B2(new_n752), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n746), .B1(new_n754), .B2(new_n755), .ZN(G1339gat));
  NAND3_X1  g555(.A1(new_n393), .A2(new_n265), .A3(new_n433), .ZN(new_n757));
  INV_X1    g556(.A(new_n609), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n758), .B(new_n592), .C1(new_n606), .C2(new_n607), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n610), .A2(KEYINPUT54), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT54), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n608), .A2(new_n761), .A3(new_n609), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n762), .A2(new_n763), .A3(new_n615), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n762), .B2(new_n615), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n760), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g567(.A(KEYINPUT55), .B(new_n760), .C1(new_n764), .C2(new_n765), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n768), .A2(new_n501), .A3(new_n616), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n484), .A2(new_n485), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n481), .B1(new_n475), .B2(new_n480), .ZN(new_n772));
  OR2_X1    g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n493), .B1(new_n490), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n618), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n641), .B1(new_n770), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n774), .A2(new_n549), .A3(new_n553), .ZN(new_n777));
  INV_X1    g576(.A(new_n760), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n615), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT111), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n762), .A2(new_n763), .A3(new_n615), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(KEYINPUT55), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n769), .A2(new_n616), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n777), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(KEYINPUT112), .B1(new_n776), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n586), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n769), .A2(new_n616), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n641), .A2(new_n788), .A3(new_n774), .A4(new_n768), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n495), .B1(new_n766), .B2(new_n767), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n788), .A2(new_n791), .B1(new_n618), .B2(new_n774), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n789), .B(new_n790), .C1(new_n792), .C2(new_n641), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n786), .A2(new_n787), .A3(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n589), .A2(new_n495), .A3(new_n590), .A4(new_n685), .ZN(new_n795));
  AOI211_X1 g594(.A(new_n396), .B(new_n757), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(G113gat), .B1(new_n796), .B2(new_n501), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n670), .B1(new_n794), .B2(new_n795), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n622), .A2(new_n265), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n798), .A2(new_n433), .A3(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n501), .A2(G113gat), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n797), .B1(new_n801), .B2(new_n802), .ZN(G1340gat));
  AOI21_X1  g602(.A(G120gat), .B1(new_n796), .B2(new_n618), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n618), .A2(G120gat), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n804), .B1(new_n801), .B2(new_n805), .ZN(G1341gat));
  AND2_X1   g605(.A1(new_n796), .A2(new_n586), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(G127gat), .B1(new_n807), .B2(new_n808), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n586), .A2(G127gat), .ZN(new_n811));
  AOI22_X1  g610(.A1(new_n809), .A2(new_n810), .B1(new_n801), .B2(new_n811), .ZN(G1342gat));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813));
  INV_X1    g612(.A(G134gat), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n801), .B2(new_n641), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n796), .A2(new_n814), .A3(new_n641), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT56), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n813), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n815), .B(KEYINPUT114), .ZN(new_n821));
  INV_X1    g620(.A(new_n819), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(KEYINPUT115), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n820), .A2(new_n823), .ZN(G1343gat));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(KEYINPUT116), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n794), .A2(new_n795), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(new_n829), .A3(new_n670), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n800), .A2(new_n631), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n501), .B1(new_n782), .B2(KEYINPUT55), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n775), .B1(new_n832), .B2(new_n784), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n554), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n586), .B1(new_n834), .B2(new_n789), .ZN(new_n835));
  INV_X1    g634(.A(new_n795), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n670), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n831), .B1(new_n837), .B2(KEYINPUT57), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n830), .A2(new_n501), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n827), .B1(new_n839), .B2(G141gat), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n396), .B1(new_n794), .B2(new_n795), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n393), .A2(new_n430), .A3(new_n266), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n495), .A2(G141gat), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n841), .A2(KEYINPUT117), .A3(new_n842), .A4(new_n843), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n840), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n839), .A2(new_n850), .A3(G141gat), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n826), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n840), .A2(new_n844), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n825), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n851), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n856), .A2(new_n840), .A3(new_n848), .ZN(new_n857));
  OAI211_X1 g656(.A(KEYINPUT118), .B(new_n853), .C1(new_n857), .C2(new_n826), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n855), .A2(new_n858), .ZN(G1344gat));
  NAND2_X1  g658(.A1(new_n841), .A2(new_n842), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(G148gat), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n862), .A3(new_n618), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n393), .B1(new_n794), .B2(new_n795), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(new_n829), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n787), .B1(new_n776), .B2(new_n785), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n795), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n868), .A2(KEYINPUT119), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n670), .A2(new_n829), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n870), .B1(new_n868), .B2(KEYINPUT119), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n866), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n872), .A2(new_n631), .A3(new_n618), .A4(new_n800), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n864), .B1(new_n873), .B2(G148gat), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n830), .A2(new_n838), .ZN(new_n875));
  AOI211_X1 g674(.A(KEYINPUT59), .B(new_n862), .C1(new_n875), .C2(new_n618), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n863), .B1(new_n874), .B2(new_n876), .ZN(G1345gat));
  AND2_X1   g676(.A1(new_n875), .A2(new_n586), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n586), .A2(new_n275), .ZN(new_n879));
  OAI22_X1  g678(.A1(new_n878), .A2(new_n275), .B1(new_n860), .B2(new_n879), .ZN(G1346gat));
  AOI21_X1  g679(.A(G162gat), .B1(new_n861), .B2(new_n641), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n554), .A2(new_n276), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n875), .B2(new_n882), .ZN(G1347gat));
  NAND2_X1  g682(.A1(new_n396), .A2(new_n266), .ZN(new_n884));
  XOR2_X1   g683(.A(new_n884), .B(KEYINPUT120), .Z(new_n885));
  NOR3_X1   g684(.A1(new_n885), .A2(new_n425), .A3(new_n422), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n798), .ZN(new_n887));
  INV_X1    g686(.A(G169gat), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n887), .A2(new_n888), .A3(new_n495), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n622), .B1(new_n794), .B2(new_n795), .ZN(new_n890));
  AND4_X1   g689(.A1(new_n266), .A2(new_n890), .A3(new_n393), .A4(new_n433), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n501), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n889), .B1(new_n892), .B2(new_n888), .ZN(G1348gat));
  INV_X1    g692(.A(G176gat), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n891), .A2(new_n894), .A3(new_n618), .ZN(new_n895));
  OAI21_X1  g694(.A(G176gat), .B1(new_n887), .B2(new_n685), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(G1349gat));
  NAND3_X1  g696(.A1(new_n891), .A2(new_n220), .A3(new_n586), .ZN(new_n898));
  OAI21_X1  g697(.A(G183gat), .B1(new_n887), .B2(new_n787), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT122), .ZN(new_n901));
  NAND2_X1  g700(.A1(KEYINPUT121), .A2(KEYINPUT60), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n898), .A2(new_n899), .A3(new_n904), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n901), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n903), .B1(new_n901), .B2(new_n905), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(G1350gat));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n221), .A3(new_n641), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT123), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n221), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n911), .B1(new_n887), .B2(new_n554), .ZN(new_n912));
  NOR2_X1   g711(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n913), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n910), .A2(new_n914), .A3(new_n915), .ZN(G1351gat));
  NAND2_X1  g715(.A1(new_n869), .A2(new_n871), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n885), .A2(new_n430), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n917), .B(new_n918), .C1(new_n865), .C2(new_n829), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n919), .A2(new_n240), .A3(new_n495), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n393), .A2(new_n430), .A3(new_n265), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n890), .A2(new_n501), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n920), .B1(new_n240), .B2(new_n922), .ZN(G1352gat));
  OAI21_X1  g722(.A(G204gat), .B1(new_n919), .B2(new_n685), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n890), .A2(new_n242), .A3(new_n618), .A4(new_n921), .ZN(new_n925));
  AND2_X1   g724(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n926));
  NOR2_X1   g725(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n924), .B(new_n928), .C1(new_n926), .C2(new_n925), .ZN(G1353gat));
  INV_X1    g728(.A(G211gat), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n919), .A2(new_n787), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n931), .B2(KEYINPUT126), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n933), .B1(new_n919), .B2(new_n787), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT63), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n872), .A2(KEYINPUT126), .A3(new_n586), .A4(new_n918), .ZN(new_n936));
  AND4_X1   g735(.A1(KEYINPUT63), .A2(new_n936), .A3(G211gat), .A4(new_n934), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n890), .A2(new_n921), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n586), .A2(new_n930), .ZN(new_n939));
  OAI22_X1  g738(.A1(new_n935), .A2(new_n937), .B1(new_n938), .B2(new_n939), .ZN(G1354gat));
  INV_X1    g739(.A(G218gat), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n919), .A2(new_n941), .A3(new_n554), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n938), .B2(new_n554), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n943), .A2(KEYINPUT127), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(KEYINPUT127), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n942), .A2(new_n944), .A3(new_n945), .ZN(G1355gat));
endmodule


