//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n621, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT66), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT67), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT68), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n453), .A2(G567), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT69), .Z(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT70), .Z(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT71), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n469), .A2(KEYINPUT71), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n466), .A2(new_n471), .A3(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n462), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n462), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT72), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g052(.A(KEYINPUT72), .B1(new_n462), .B2(G2104), .ZN(new_n478));
  OAI21_X1  g053(.A(G101), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g054(.A(G137), .B(new_n462), .C1(new_n464), .C2(new_n465), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n474), .A2(new_n481), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT73), .Z(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  NOR2_X1   g059(.A1(new_n464), .A2(new_n465), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(new_n462), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G112), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(G2105), .ZN(new_n491));
  OR3_X1    g066(.A1(new_n485), .A2(KEYINPUT74), .A3(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT74), .B1(new_n485), .B2(G2105), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI211_X1 g069(.A(new_n488), .B(new_n491), .C1(new_n494), .C2(G136), .ZN(G162));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(G2105), .ZN(new_n498));
  AND2_X1   g073(.A1(G126), .A2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(new_n464), .B2(new_n465), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT75), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(KEYINPUT75), .B(new_n499), .C1(new_n464), .C2(new_n465), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n498), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G138), .ZN(new_n505));
  NOR3_X1   g080(.A1(new_n505), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n466), .A2(new_n471), .A3(new_n506), .ZN(new_n507));
  OAI211_X1 g082(.A(G138), .B(new_n462), .C1(new_n464), .C2(new_n465), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT4), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  OR2_X1    g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n520), .A2(G88), .B1(G50), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n523), .A2(new_n526), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n520), .A2(G89), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n517), .A2(new_n518), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G51), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT76), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n529), .B(new_n530), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n535), .A2(new_n536), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(G168));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n532), .A2(new_n515), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n540), .A2(new_n533), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n525), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n543), .A2(new_n545), .ZN(G171));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n547), .A2(new_n533), .B1(new_n541), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n525), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g129(.A(KEYINPUT77), .B(KEYINPUT8), .Z(new_n555));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  INV_X1    g134(.A(G78), .ZN(new_n560));
  OAI22_X1  g135(.A1(new_n516), .A2(new_n559), .B1(new_n560), .B2(new_n521), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT78), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT78), .ZN(new_n563));
  OAI221_X1 g138(.A(new_n563), .B1(new_n560), .B2(new_n521), .C1(new_n516), .C2(new_n559), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(G651), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n532), .A2(G53), .A3(G543), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(KEYINPUT9), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n522), .A2(new_n568), .A3(G53), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n567), .A2(new_n569), .B1(G91), .B2(new_n520), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n565), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  XNOR2_X1  g148(.A(G166), .B(KEYINPUT79), .ZN(G303));
  AOI22_X1  g149(.A1(new_n520), .A2(G87), .B1(G49), .B2(new_n522), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n576), .A2(KEYINPUT80), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(KEYINPUT80), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(G288));
  INV_X1    g154(.A(G48), .ZN(new_n580));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  OAI22_X1  g156(.A1(new_n580), .A2(new_n533), .B1(new_n541), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n513), .B2(new_n514), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT81), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n589), .B1(new_n585), .B2(new_n586), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n583), .A2(new_n591), .ZN(G305));
  AOI22_X1  g167(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n593), .A2(new_n525), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  INV_X1    g170(.A(G85), .ZN(new_n596));
  OAI221_X1 g171(.A(new_n594), .B1(new_n595), .B2(new_n533), .C1(new_n596), .C2(new_n541), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT82), .ZN(new_n599));
  XNOR2_X1  g174(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT84), .ZN(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n541), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT84), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n600), .B(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n605), .A2(G92), .A3(new_n520), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(G54), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT85), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n608), .B1(new_n533), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n609), .B2(new_n533), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  XNOR2_X1  g187(.A(KEYINPUT86), .B(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n516), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G651), .ZN(new_n615));
  AND3_X1   g190(.A1(new_n607), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n599), .B1(G868), .B2(new_n616), .ZN(G284));
  OAI21_X1  g192(.A(new_n599), .B1(G868), .B2(new_n616), .ZN(G321));
  MUX2_X1   g193(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g194(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n616), .B1(new_n621), .B2(G860), .ZN(G148));
  NAND2_X1  g197(.A1(new_n616), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g201(.A(new_n475), .B(new_n476), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n627), .A2(new_n466), .A3(new_n471), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  INV_X1    g204(.A(G2100), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT87), .B(KEYINPUT13), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(G111), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(G2105), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n636), .B1(new_n486), .B2(G123), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n492), .A2(new_n493), .ZN(new_n638));
  INV_X1    g213(.A(G135), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT88), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT89), .B(G2096), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n633), .A2(new_n643), .ZN(G156));
  INV_X1    g219(.A(KEYINPUT14), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(new_n648), .B2(new_n647), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n650), .B(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(G14), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n658), .B2(new_n656), .ZN(G401));
  INV_X1    g235(.A(KEYINPUT18), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n661), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(new_n630), .ZN(new_n668));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n664), .B2(KEYINPUT18), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(G2096), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT19), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n676), .A2(new_n677), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n675), .A2(new_n682), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n675), .A2(new_n678), .A3(new_n682), .ZN(new_n684));
  NOR3_X1   g259(.A1(new_n681), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(G229));
  NOR2_X1   g266(.A1(G16), .A2(G19), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(new_n552), .B2(G16), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT94), .Z(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(G1341), .Z(new_n695));
  NOR2_X1   g270(.A1(G4), .A2(G16), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n616), .B2(G16), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT93), .B(G1348), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n697), .B(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G27), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G164), .B2(new_n701), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n703), .A2(G2078), .ZN(new_n704));
  INV_X1    g279(.A(G1961), .ZN(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NOR2_X1   g281(.A1(G171), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G5), .B2(new_n706), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n704), .B1(new_n705), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G2078), .B2(new_n703), .ZN(new_n710));
  NOR3_X1   g285(.A1(new_n695), .A2(new_n700), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT96), .B(KEYINPUT28), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n701), .A2(G26), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n494), .A2(G140), .ZN(new_n715));
  NOR2_X1   g290(.A1(G104), .A2(G2105), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT95), .Z(new_n717));
  INV_X1    g292(.A(G116), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n468), .B1(new_n718), .B2(G2105), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n717), .A2(new_n719), .B1(new_n486), .B2(G128), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n714), .B1(new_n721), .B2(G29), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G2067), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n701), .A2(G33), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT25), .Z(new_n726));
  INV_X1    g301(.A(G139), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(new_n638), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n466), .A2(new_n471), .A3(G127), .ZN(new_n729));
  NAND2_X1  g304(.A1(G115), .A2(G2104), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n462), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n724), .B1(new_n732), .B2(new_n701), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G2072), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(G2072), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n723), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n701), .A2(G32), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n494), .A2(G141), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT97), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n627), .A2(G105), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT98), .ZN(new_n741));
  NAND3_X1  g316(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT26), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n486), .A2(G129), .ZN(new_n744));
  AND3_X1   g319(.A1(new_n741), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n739), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n737), .B1(new_n746), .B2(G29), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT27), .B(G1996), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n747), .A2(new_n749), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n736), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT102), .B(KEYINPUT23), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n706), .A2(G20), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G299), .B2(G16), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1956), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n701), .A2(G35), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G162), .B2(new_n701), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n759), .A2(KEYINPUT29), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(KEYINPUT29), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G2090), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n757), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(KEYINPUT103), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT103), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n766), .B(new_n757), .C1(new_n762), .C2(new_n763), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n711), .A2(new_n752), .A3(new_n765), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT31), .B(G11), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n770), .A2(G28), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n701), .B1(new_n770), .B2(G28), .ZN(new_n772));
  OAI221_X1 g347(.A(new_n769), .B1(new_n771), .B2(new_n772), .C1(new_n708), .C2(new_n705), .ZN(new_n773));
  INV_X1    g348(.A(G1966), .ZN(new_n774));
  NOR2_X1   g349(.A1(G168), .A2(new_n706), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n706), .B2(G21), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n773), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n641), .A2(G29), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT99), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n776), .A2(new_n774), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n777), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(KEYINPUT100), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT100), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n777), .A2(new_n780), .A3(new_n784), .A4(new_n781), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT24), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n786), .A2(G34), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(G34), .ZN(new_n788));
  AOI21_X1  g363(.A(G29), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n483), .B2(G29), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G2084), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n760), .A2(new_n763), .A3(new_n761), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT101), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n783), .A2(new_n785), .A3(new_n791), .A4(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n768), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n706), .A2(G23), .ZN(new_n796));
  INV_X1    g371(.A(G288), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n706), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT33), .B(G1976), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(G6), .A2(G16), .ZN(new_n801));
  INV_X1    g376(.A(new_n590), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(new_n587), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n582), .B1(new_n803), .B2(G651), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n801), .B1(new_n804), .B2(G16), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT32), .B(G1981), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n706), .A2(G22), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT92), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G166), .B2(new_n706), .ZN(new_n810));
  INV_X1    g385(.A(G1971), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n798), .A2(new_n799), .ZN(new_n813));
  AND4_X1   g388(.A1(new_n800), .A2(new_n807), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT34), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n706), .A2(G24), .ZN(new_n818));
  INV_X1    g393(.A(G290), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(new_n706), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G1986), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n486), .A2(G119), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT91), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n494), .A2(G131), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n462), .A2(G107), .ZN(new_n825));
  OAI21_X1  g400(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n823), .B(new_n824), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  MUX2_X1   g402(.A(G25), .B(new_n827), .S(G29), .Z(new_n828));
  XOR2_X1   g403(.A(KEYINPUT35), .B(G1991), .Z(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n828), .A2(new_n830), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n821), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n816), .A2(new_n817), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT36), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT36), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n816), .A2(new_n836), .A3(new_n817), .A4(new_n833), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n795), .A2(new_n838), .ZN(G311));
  INV_X1    g414(.A(KEYINPUT104), .ZN(new_n840));
  AND3_X1   g415(.A1(new_n795), .A2(new_n840), .A3(new_n838), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n840), .B1(new_n795), .B2(new_n838), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(new_n842), .ZN(G150));
  NAND2_X1  g418(.A1(new_n616), .A2(G559), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  INV_X1    g420(.A(G55), .ZN(new_n846));
  INV_X1    g421(.A(G93), .ZN(new_n847));
  OAI22_X1  g422(.A1(new_n846), .A2(new_n533), .B1(new_n541), .B2(new_n847), .ZN(new_n848));
  AOI22_X1  g423(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n849), .A2(new_n525), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n552), .A2(new_n851), .ZN(new_n852));
  OAI22_X1  g427(.A1(new_n549), .A2(new_n551), .B1(new_n848), .B2(new_n850), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n845), .B(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n856), .A2(KEYINPUT39), .ZN(new_n857));
  INV_X1    g432(.A(G860), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(KEYINPUT39), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n851), .A2(new_n858), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(G145));
  XNOR2_X1  g438(.A(new_n483), .B(new_n641), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(G162), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n827), .B(new_n629), .Z(new_n866));
  INV_X1    g441(.A(new_n732), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n746), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n739), .A2(new_n745), .A3(new_n732), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n827), .B(new_n629), .ZN(new_n871));
  INV_X1    g446(.A(new_n869), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n732), .B1(new_n739), .B2(new_n745), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT105), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n507), .A2(new_n509), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n876), .B1(new_n507), .B2(new_n509), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n504), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n721), .B(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n486), .A2(G130), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n462), .A2(G118), .ZN(new_n882));
  OAI21_X1  g457(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n883));
  INV_X1    g458(.A(G142), .ZN(new_n884));
  OAI221_X1 g459(.A(new_n881), .B1(new_n882), .B2(new_n883), .C1(new_n638), .C2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n880), .B(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n875), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n870), .A3(new_n874), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n865), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT107), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n865), .A3(new_n889), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT106), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n888), .A2(new_n865), .A3(KEYINPUT106), .A4(new_n889), .ZN(new_n895));
  AOI21_X1  g470(.A(G37), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n891), .A2(KEYINPUT40), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT40), .B1(new_n891), .B2(new_n896), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(G395));
  NAND2_X1  g474(.A1(G299), .A2(KEYINPUT108), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n565), .A2(new_n570), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n616), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT41), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n607), .A2(new_n611), .A3(new_n615), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n905), .A2(KEYINPUT108), .A3(G299), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n904), .B1(new_n903), .B2(new_n906), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT109), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n623), .B(new_n855), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT109), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n903), .A2(new_n906), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n911), .B1(new_n912), .B2(KEYINPUT41), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n909), .A2(new_n910), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n912), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT42), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n819), .A2(new_n797), .ZN(new_n919));
  NAND2_X1  g494(.A1(G290), .A2(G288), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT110), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n804), .B(G166), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT110), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n919), .A2(new_n925), .A3(new_n920), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n922), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n928), .A2(KEYINPUT111), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT42), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n914), .A2(new_n930), .A3(new_n916), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n918), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n929), .B1(new_n918), .B2(new_n931), .ZN(new_n933));
  OAI21_X1  g508(.A(G868), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(G868), .B2(new_n851), .ZN(G295));
  OAI21_X1  g510(.A(new_n934), .B1(G868), .B2(new_n851), .ZN(G331));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n852), .A2(new_n853), .A3(G301), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(G301), .B1(new_n852), .B2(new_n853), .ZN(new_n940));
  OAI21_X1  g515(.A(G286), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n940), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n942), .A2(G168), .A3(new_n938), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n944), .B1(new_n909), .B2(new_n913), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n912), .B1(new_n941), .B2(new_n943), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n945), .A2(new_n928), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G37), .ZN(new_n948));
  INV_X1    g523(.A(new_n944), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n912), .A2(KEYINPUT41), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n946), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n924), .A2(new_n927), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n948), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT112), .B1(new_n947), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n949), .A2(new_n952), .ZN(new_n957));
  INV_X1    g532(.A(new_n946), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(G37), .B1(new_n959), .B2(new_n928), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n911), .B1(new_n950), .B2(new_n951), .ZN(new_n962));
  INV_X1    g537(.A(new_n913), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n949), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(new_n954), .A3(new_n958), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n960), .A2(new_n961), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n956), .A2(new_n966), .A3(KEYINPUT43), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n928), .B1(new_n945), .B2(new_n946), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n968), .A2(new_n965), .A3(new_n969), .A4(new_n948), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n937), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n968), .A2(new_n965), .A3(new_n948), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n960), .A2(new_n969), .A3(new_n965), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n973), .A2(new_n937), .A3(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n971), .A2(new_n975), .ZN(G397));
  INV_X1    g551(.A(new_n746), .ZN(new_n977));
  INV_X1    g552(.A(G1384), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT45), .B1(new_n879), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G40), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n474), .A2(new_n980), .A3(new_n481), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(G1996), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n977), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT114), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n982), .B(KEYINPUT115), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n721), .A2(G2067), .ZN(new_n987));
  INV_X1    g562(.A(G2067), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n715), .A2(new_n988), .A3(new_n720), .ZN(new_n989));
  INV_X1    g564(.A(G1996), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n987), .B(new_n989), .C1(new_n977), .C2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n985), .B1(new_n986), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n827), .B(new_n829), .ZN(new_n993));
  INV_X1    g568(.A(new_n986), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OR3_X1    g570(.A1(new_n982), .A2(G1986), .A3(G290), .ZN(new_n996));
  NAND2_X1  g571(.A1(G290), .A2(G1986), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n996), .B1(new_n982), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT113), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1001), .A2(G1384), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n511), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n981), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n774), .B1(new_n979), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1006), .B1(new_n511), .B2(new_n978), .ZN(new_n1007));
  INV_X1    g582(.A(new_n481), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n472), .A2(new_n473), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1008), .B(G40), .C1(new_n1009), .C2(new_n462), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G2084), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n879), .A2(new_n1006), .A3(new_n978), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1005), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(G8), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT126), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT51), .ZN(new_n1018));
  INV_X1    g593(.A(G8), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1018), .B1(G168), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1017), .A2(KEYINPUT51), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1016), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1019), .B1(new_n1005), .B2(new_n1014), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1022), .B1(new_n1025), .B2(new_n1020), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT62), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1015), .A2(G8), .A3(G286), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n502), .A2(new_n503), .ZN(new_n1030));
  INV_X1    g605(.A(new_n498), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n510), .A2(KEYINPUT105), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n507), .A2(new_n509), .A3(new_n876), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1032), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1035), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1036));
  AOI21_X1  g611(.A(G1384), .B1(new_n504), .B2(new_n510), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n981), .B1(new_n1006), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n705), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n981), .A2(new_n1003), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(G2078), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1035), .A2(G1384), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1040), .B(new_n1042), .C1(new_n1043), .C2(KEYINPUT45), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1039), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G2078), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n879), .A2(new_n1002), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n511), .A2(new_n978), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n1001), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1047), .A2(new_n1049), .A3(KEYINPUT116), .A4(new_n981), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT45), .B1(new_n511), .B2(new_n978), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(new_n1010), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT116), .B1(new_n1053), .B2(new_n1047), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1046), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1045), .B1(new_n1055), .B2(new_n1041), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1056), .A2(G301), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1029), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(G305), .A2(G1981), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(G305), .A2(G1981), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT49), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OR2_X1    g637(.A1(G305), .A2(G1981), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT49), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(new_n1064), .A3(new_n1059), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n879), .A2(new_n981), .A3(new_n978), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(G8), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT118), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1067), .A2(new_n1070), .A3(G8), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1066), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n797), .A2(G1976), .ZN(new_n1074));
  INV_X1    g649(.A(G1976), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT52), .B1(G288), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1071), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1070), .B1(new_n1067), .B2(G8), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1074), .B(new_n1076), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1069), .A2(new_n1071), .B1(G1976), .B2(new_n797), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1073), .B(new_n1079), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1002), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1035), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n981), .B1(KEYINPUT45), .B2(new_n1037), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1083), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1087), .A2(new_n811), .A3(new_n1050), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1011), .A2(new_n763), .A3(new_n1013), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G8), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1089), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(G303), .A2(G8), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT55), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1082), .B1(new_n1094), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1099), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1087), .A2(new_n811), .A3(new_n1050), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n879), .A2(new_n978), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1010), .B1(new_n1103), .B2(KEYINPUT50), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT119), .B1(new_n1048), .B2(KEYINPUT50), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1037), .A2(new_n1106), .A3(new_n1006), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n1110));
  AOI21_X1  g685(.A(G2090), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1104), .A2(new_n1108), .A3(KEYINPUT120), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1102), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1101), .B1(new_n1113), .B2(new_n1019), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1058), .A2(new_n1100), .A3(KEYINPUT127), .A4(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT127), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1118), .A2(G8), .A3(new_n1099), .A4(new_n1091), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1073), .A2(new_n1079), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1081), .A2(new_n1080), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1114), .A2(new_n1119), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1029), .A2(new_n1057), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1116), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1024), .A2(new_n1028), .A3(new_n1026), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n1126), .A2(new_n1027), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1115), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1062), .A2(new_n1065), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n797), .A2(new_n1075), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1063), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n1072), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n1119), .B2(new_n1082), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT121), .B1(new_n1016), .B2(G286), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1025), .A2(new_n1135), .A3(G168), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1122), .B(new_n1137), .C1(new_n1094), .C2(new_n1099), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1133), .B1(new_n1138), .B2(KEYINPUT63), .ZN(new_n1139));
  AOI21_X1  g714(.A(KEYINPUT63), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n879), .A2(new_n981), .A3(new_n978), .A4(new_n988), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT123), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n699), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1141), .A2(KEYINPUT123), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT124), .B1(new_n1146), .B2(new_n905), .ZN(new_n1147));
  XNOR2_X1  g722(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(G2072), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1085), .A2(new_n1086), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(G1956), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1150), .B1(new_n1109), .B2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g727(.A(G299), .B(KEYINPUT57), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n698), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1043), .A2(new_n1157), .A3(new_n988), .A4(new_n981), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1156), .A2(new_n1142), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(new_n1160), .A3(new_n616), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1147), .A2(new_n1155), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(G1956), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1153), .B1(new_n1163), .B2(new_n1150), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT61), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n1166));
  NOR4_X1   g741(.A1(new_n1163), .A2(new_n1153), .A3(new_n1150), .A4(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1159), .A2(KEYINPUT60), .A3(new_n616), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1170));
  OR2_X1    g745(.A1(new_n616), .A2(KEYINPUT60), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n616), .A2(KEYINPUT60), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1170), .A2(new_n1142), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1047), .A2(new_n1049), .A3(new_n990), .A4(new_n981), .ZN(new_n1174));
  XOR2_X1   g749(.A(KEYINPUT58), .B(G1341), .Z(new_n1175));
  NAND2_X1  g750(.A1(new_n1067), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n552), .A2(KEYINPUT125), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT59), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1177), .A2(KEYINPUT59), .A3(new_n1178), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1169), .A2(new_n1173), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  OAI211_X1 g758(.A(new_n1162), .B(new_n1164), .C1(new_n1168), .C2(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g759(.A(G171), .B(KEYINPUT54), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1047), .A2(new_n981), .A3(new_n1042), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1185), .B1(new_n1186), .B2(new_n979), .ZN(new_n1187));
  AOI21_X1  g762(.A(G1961), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(G2078), .B1(new_n1087), .B2(new_n1050), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1189), .B1(KEYINPUT53), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1191), .B1(new_n1056), .B2(new_n1185), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1126), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1140), .B1(new_n1184), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1139), .B1(new_n1194), .B2(new_n1123), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1000), .B1(new_n1128), .B2(new_n1195), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n983), .B(KEYINPUT46), .Z(new_n1197));
  NAND2_X1  g772(.A1(new_n987), .A2(new_n989), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n986), .B1(new_n746), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1200), .B(KEYINPUT47), .ZN(new_n1201));
  XOR2_X1   g776(.A(new_n996), .B(KEYINPUT48), .Z(new_n1202));
  OAI21_X1  g777(.A(new_n1201), .B1(new_n995), .B2(new_n1202), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n827), .A2(new_n830), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n992), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n994), .B1(new_n1205), .B2(new_n989), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1203), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1196), .A2(new_n1207), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g783(.A(G227), .ZN(new_n1210));
  NAND2_X1  g784(.A1(G319), .A2(new_n1210), .ZN(new_n1211));
  OR2_X1    g785(.A1(new_n1211), .A2(G401), .ZN(new_n1212));
  OR2_X1    g786(.A1(new_n1212), .A2(G229), .ZN(new_n1213));
  INV_X1    g787(.A(new_n1213), .ZN(new_n1214));
  NAND2_X1  g788(.A1(new_n891), .A2(new_n896), .ZN(new_n1215));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n974), .ZN(new_n1216));
  AND3_X1   g790(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(G308));
  NAND3_X1  g791(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(G225));
endmodule


