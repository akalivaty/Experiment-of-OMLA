

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579;

  NOR2_X1 U319 ( .A1(n467), .A2(n415), .ZN(n417) );
  NOR2_X1 U320 ( .A1(n467), .A2(n563), .ZN(n468) );
  AND2_X1 U321 ( .A1(G230GAT), .A2(G233GAT), .ZN(n287) );
  OR2_X1 U322 ( .A1(n511), .A2(n513), .ZN(n414) );
  XNOR2_X1 U323 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n359) );
  NOR2_X1 U324 ( .A1(n521), .A2(n464), .ZN(n465) );
  XNOR2_X1 U325 ( .A(n308), .B(n287), .ZN(n309) );
  INV_X1 U326 ( .A(KEYINPUT33), .ZN(n316) );
  XNOR2_X1 U327 ( .A(n310), .B(n309), .ZN(n313) );
  XNOR2_X1 U328 ( .A(KEYINPUT107), .B(KEYINPUT37), .ZN(n445) );
  XNOR2_X1 U329 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U330 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U331 ( .A(n446), .B(n445), .ZN(n507) );
  XNOR2_X1 U332 ( .A(n374), .B(n373), .ZN(n522) );
  XNOR2_X1 U333 ( .A(n319), .B(n318), .ZN(n569) );
  NOR2_X1 U334 ( .A1(n513), .A2(n469), .ZN(n558) );
  XNOR2_X1 U335 ( .A(KEYINPUT38), .B(n448), .ZN(n493) );
  XNOR2_X1 U336 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n470) );
  INV_X1 U337 ( .A(G36GAT), .ZN(n449) );
  XNOR2_X1 U338 ( .A(n471), .B(n470), .ZN(G1351GAT) );
  XNOR2_X1 U339 ( .A(n450), .B(n449), .ZN(G1329GAT) );
  XNOR2_X1 U340 ( .A(KEYINPUT85), .B(KEYINPUT18), .ZN(n288) );
  XNOR2_X1 U341 ( .A(n288), .B(KEYINPUT17), .ZN(n289) );
  XOR2_X1 U342 ( .A(n289), .B(KEYINPUT19), .Z(n291) );
  XNOR2_X1 U343 ( .A(G183GAT), .B(G190GAT), .ZN(n290) );
  XNOR2_X1 U344 ( .A(n291), .B(n290), .ZN(n368) );
  XOR2_X1 U345 ( .A(KEYINPUT21), .B(G218GAT), .Z(n293) );
  XNOR2_X1 U346 ( .A(KEYINPUT89), .B(G211GAT), .ZN(n292) );
  XNOR2_X1 U347 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U348 ( .A(G197GAT), .B(n294), .Z(n378) );
  XNOR2_X1 U349 ( .A(n368), .B(n378), .ZN(n305) );
  XOR2_X1 U350 ( .A(G64GAT), .B(KEYINPUT74), .Z(n296) );
  XNOR2_X1 U351 ( .A(G204GAT), .B(G92GAT), .ZN(n295) );
  XNOR2_X1 U352 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U353 ( .A(G176GAT), .B(n297), .Z(n311) );
  XOR2_X1 U354 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n300) );
  XNOR2_X1 U355 ( .A(G169GAT), .B(G36GAT), .ZN(n298) );
  XNOR2_X1 U356 ( .A(n298), .B(G8GAT), .ZN(n326) );
  XNOR2_X1 U357 ( .A(n326), .B(KEYINPUT98), .ZN(n299) );
  XNOR2_X1 U358 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U359 ( .A(n311), .B(n301), .Z(n303) );
  NAND2_X1 U360 ( .A1(G226GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U361 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U362 ( .A(n305), .B(n304), .Z(n511) );
  XOR2_X1 U363 ( .A(G99GAT), .B(G85GAT), .Z(n434) );
  XOR2_X1 U364 ( .A(G57GAT), .B(KEYINPUT13), .Z(n338) );
  XOR2_X1 U365 ( .A(n434), .B(n338), .Z(n310) );
  XOR2_X1 U366 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n307) );
  XNOR2_X1 U367 ( .A(KEYINPUT32), .B(KEYINPUT72), .ZN(n306) );
  XNOR2_X1 U368 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U369 ( .A(G120GAT), .B(G71GAT), .Z(n355) );
  XNOR2_X1 U370 ( .A(n355), .B(n311), .ZN(n312) );
  XNOR2_X1 U371 ( .A(n313), .B(n312), .ZN(n319) );
  XOR2_X1 U372 ( .A(G78GAT), .B(G148GAT), .Z(n315) );
  XNOR2_X1 U373 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n314) );
  XNOR2_X1 U374 ( .A(n315), .B(n314), .ZN(n385) );
  XNOR2_X1 U375 ( .A(n385), .B(KEYINPUT31), .ZN(n317) );
  XOR2_X1 U376 ( .A(KEYINPUT29), .B(KEYINPUT65), .Z(n321) );
  XNOR2_X1 U377 ( .A(G197GAT), .B(G113GAT), .ZN(n320) );
  XNOR2_X1 U378 ( .A(n321), .B(n320), .ZN(n330) );
  XOR2_X1 U379 ( .A(G141GAT), .B(G22GAT), .Z(n386) );
  XNOR2_X1 U380 ( .A(G15GAT), .B(G1GAT), .ZN(n322) );
  XNOR2_X1 U381 ( .A(n322), .B(KEYINPUT68), .ZN(n342) );
  XOR2_X1 U382 ( .A(n386), .B(n342), .Z(n324) );
  NAND2_X1 U383 ( .A1(G229GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U384 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U385 ( .A(n325), .B(KEYINPUT30), .Z(n328) );
  XNOR2_X1 U386 ( .A(n326), .B(KEYINPUT66), .ZN(n327) );
  XNOR2_X1 U387 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n335) );
  XOR2_X1 U389 ( .A(G29GAT), .B(KEYINPUT67), .Z(n332) );
  XNOR2_X1 U390 ( .A(G50GAT), .B(G43GAT), .ZN(n331) );
  XNOR2_X1 U391 ( .A(n332), .B(n331), .ZN(n334) );
  XOR2_X1 U392 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n333) );
  XOR2_X1 U393 ( .A(n334), .B(n333), .Z(n427) );
  XOR2_X1 U394 ( .A(n335), .B(n427), .Z(n537) );
  INV_X1 U395 ( .A(n537), .ZN(n566) );
  XOR2_X1 U396 ( .A(KEYINPUT69), .B(n566), .Z(n550) );
  INV_X1 U397 ( .A(n550), .ZN(n459) );
  NOR2_X1 U398 ( .A1(n569), .A2(n459), .ZN(n476) );
  XOR2_X1 U399 ( .A(G155GAT), .B(G211GAT), .Z(n337) );
  XNOR2_X1 U400 ( .A(G183GAT), .B(G127GAT), .ZN(n336) );
  XNOR2_X1 U401 ( .A(n337), .B(n336), .ZN(n339) );
  XOR2_X1 U402 ( .A(n339), .B(n338), .Z(n341) );
  XNOR2_X1 U403 ( .A(G22GAT), .B(G78GAT), .ZN(n340) );
  XNOR2_X1 U404 ( .A(n341), .B(n340), .ZN(n346) );
  XOR2_X1 U405 ( .A(n342), .B(KEYINPUT12), .Z(n344) );
  NAND2_X1 U406 ( .A1(G231GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U407 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U408 ( .A(n346), .B(n345), .Z(n354) );
  XOR2_X1 U409 ( .A(KEYINPUT78), .B(G64GAT), .Z(n348) );
  XNOR2_X1 U410 ( .A(G8GAT), .B(G71GAT), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U412 ( .A(KEYINPUT77), .B(KEYINPUT15), .Z(n350) );
  XNOR2_X1 U413 ( .A(KEYINPUT76), .B(KEYINPUT14), .ZN(n349) );
  XNOR2_X1 U414 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U415 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U416 ( .A(n354), .B(n353), .Z(n573) );
  INV_X1 U417 ( .A(n573), .ZN(n544) );
  XOR2_X1 U418 ( .A(n355), .B(KEYINPUT84), .Z(n357) );
  NAND2_X1 U419 ( .A1(G227GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U420 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U421 ( .A(n358), .B(G99GAT), .Z(n364) );
  XNOR2_X1 U422 ( .A(n359), .B(KEYINPUT80), .ZN(n360) );
  XOR2_X1 U423 ( .A(n360), .B(KEYINPUT79), .Z(n362) );
  XNOR2_X1 U424 ( .A(G113GAT), .B(G134GAT), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n362), .B(n361), .ZN(n406) );
  XNOR2_X1 U426 ( .A(G43GAT), .B(n406), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n364), .B(n363), .ZN(n374) );
  XOR2_X1 U428 ( .A(KEYINPUT86), .B(KEYINPUT83), .Z(n366) );
  XNOR2_X1 U429 ( .A(KEYINPUT20), .B(KEYINPUT82), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U431 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U432 ( .A(G176GAT), .B(KEYINPUT81), .Z(n370) );
  XNOR2_X1 U433 ( .A(G169GAT), .B(G15GAT), .ZN(n369) );
  XNOR2_X1 U434 ( .A(n370), .B(n369), .ZN(n371) );
  INV_X1 U435 ( .A(n522), .ZN(n513) );
  XOR2_X1 U436 ( .A(KEYINPUT90), .B(G162GAT), .Z(n376) );
  XNOR2_X1 U437 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U439 ( .A(KEYINPUT3), .B(n377), .Z(n405) );
  XNOR2_X1 U440 ( .A(n378), .B(n405), .ZN(n393) );
  XOR2_X1 U441 ( .A(G204GAT), .B(KEYINPUT87), .Z(n380) );
  XNOR2_X1 U442 ( .A(KEYINPUT22), .B(KEYINPUT92), .ZN(n379) );
  XNOR2_X1 U443 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U444 ( .A(KEYINPUT91), .B(n381), .Z(n383) );
  NAND2_X1 U445 ( .A1(G228GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U446 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U447 ( .A(n384), .B(KEYINPUT23), .Z(n391) );
  XOR2_X1 U448 ( .A(n385), .B(KEYINPUT88), .Z(n388) );
  XNOR2_X1 U449 ( .A(G50GAT), .B(n386), .ZN(n387) );
  XNOR2_X1 U450 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n389), .B(KEYINPUT24), .ZN(n390) );
  XNOR2_X1 U452 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U453 ( .A(n393), .B(n392), .ZN(n467) );
  XNOR2_X1 U454 ( .A(n467), .B(KEYINPUT64), .ZN(n394) );
  XOR2_X1 U455 ( .A(n394), .B(KEYINPUT28), .Z(n516) );
  INV_X1 U456 ( .A(n516), .ZN(n525) );
  XOR2_X1 U457 ( .A(G57GAT), .B(G148GAT), .Z(n396) );
  XNOR2_X1 U458 ( .A(G141GAT), .B(G120GAT), .ZN(n395) );
  XNOR2_X1 U459 ( .A(n396), .B(n395), .ZN(n398) );
  XOR2_X1 U460 ( .A(G29GAT), .B(G85GAT), .Z(n397) );
  XNOR2_X1 U461 ( .A(n398), .B(n397), .ZN(n410) );
  XOR2_X1 U462 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n400) );
  XNOR2_X1 U463 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n399) );
  XNOR2_X1 U464 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U465 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n402) );
  XNOR2_X1 U466 ( .A(KEYINPUT93), .B(KEYINPUT6), .ZN(n401) );
  XNOR2_X1 U467 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U468 ( .A(n404), .B(n403), .Z(n408) );
  XNOR2_X1 U469 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U470 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U471 ( .A(n410), .B(n409), .ZN(n412) );
  NAND2_X1 U472 ( .A1(G225GAT), .A2(G233GAT), .ZN(n411) );
  XOR2_X1 U473 ( .A(n412), .B(n411), .Z(n423) );
  XOR2_X1 U474 ( .A(n511), .B(KEYINPUT27), .Z(n419) );
  NAND2_X1 U475 ( .A1(n423), .A2(n419), .ZN(n520) );
  NOR2_X1 U476 ( .A1(n525), .A2(n520), .ZN(n413) );
  NAND2_X1 U477 ( .A1(n513), .A2(n413), .ZN(n426) );
  XOR2_X1 U478 ( .A(KEYINPUT100), .B(n414), .Z(n415) );
  XOR2_X1 U479 ( .A(KEYINPUT25), .B(KEYINPUT101), .Z(n416) );
  XNOR2_X1 U480 ( .A(n417), .B(n416), .ZN(n422) );
  NAND2_X1 U481 ( .A1(n467), .A2(n513), .ZN(n418) );
  XOR2_X1 U482 ( .A(n418), .B(KEYINPUT26), .Z(n565) );
  AND2_X1 U483 ( .A1(n419), .A2(n565), .ZN(n420) );
  XNOR2_X1 U484 ( .A(KEYINPUT99), .B(n420), .ZN(n421) );
  NAND2_X1 U485 ( .A1(n422), .A2(n421), .ZN(n424) );
  INV_X1 U486 ( .A(n423), .ZN(n508) );
  NAND2_X1 U487 ( .A1(n424), .A2(n508), .ZN(n425) );
  NAND2_X1 U488 ( .A1(n426), .A2(n425), .ZN(n473) );
  NAND2_X1 U489 ( .A1(n544), .A2(n473), .ZN(n444) );
  INV_X1 U490 ( .A(n427), .ZN(n431) );
  XOR2_X1 U491 ( .A(G106GAT), .B(G134GAT), .Z(n429) );
  XNOR2_X1 U492 ( .A(G36GAT), .B(G190GAT), .ZN(n428) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U494 ( .A(n431), .B(n430), .Z(n442) );
  XOR2_X1 U495 ( .A(KEYINPUT75), .B(KEYINPUT11), .Z(n433) );
  XNOR2_X1 U496 ( .A(G162GAT), .B(KEYINPUT9), .ZN(n432) );
  XNOR2_X1 U497 ( .A(n433), .B(n432), .ZN(n438) );
  XOR2_X1 U498 ( .A(G92GAT), .B(KEYINPUT10), .Z(n436) );
  XNOR2_X1 U499 ( .A(G218GAT), .B(n434), .ZN(n435) );
  XNOR2_X1 U500 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U501 ( .A(n438), .B(n437), .Z(n440) );
  NAND2_X1 U502 ( .A1(G232GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U503 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U504 ( .A(n442), .B(n441), .Z(n548) );
  XOR2_X1 U505 ( .A(KEYINPUT36), .B(KEYINPUT106), .Z(n443) );
  XOR2_X1 U506 ( .A(n548), .B(n443), .Z(n576) );
  NOR2_X1 U507 ( .A1(n444), .A2(n576), .ZN(n446) );
  NAND2_X1 U508 ( .A1(n476), .A2(n507), .ZN(n447) );
  XNOR2_X1 U509 ( .A(n447), .B(KEYINPUT108), .ZN(n448) );
  NOR2_X1 U510 ( .A1(n511), .A2(n493), .ZN(n450) );
  INV_X1 U511 ( .A(n548), .ZN(n531) );
  XOR2_X1 U512 ( .A(KEYINPUT116), .B(KEYINPUT46), .Z(n452) );
  XNOR2_X1 U513 ( .A(KEYINPUT41), .B(n569), .ZN(n540) );
  INV_X1 U514 ( .A(n540), .ZN(n555) );
  NAND2_X1 U515 ( .A1(n555), .A2(n566), .ZN(n451) );
  XNOR2_X1 U516 ( .A(n452), .B(n451), .ZN(n453) );
  NOR2_X1 U517 ( .A1(n531), .A2(n453), .ZN(n454) );
  NAND2_X1 U518 ( .A1(n544), .A2(n454), .ZN(n455) );
  XNOR2_X1 U519 ( .A(KEYINPUT47), .B(n455), .ZN(n456) );
  XNOR2_X1 U520 ( .A(n456), .B(KEYINPUT117), .ZN(n462) );
  NOR2_X1 U521 ( .A1(n544), .A2(n576), .ZN(n457) );
  XOR2_X1 U522 ( .A(KEYINPUT45), .B(n457), .Z(n458) );
  NOR2_X1 U523 ( .A1(n569), .A2(n458), .ZN(n460) );
  NAND2_X1 U524 ( .A1(n460), .A2(n459), .ZN(n461) );
  NAND2_X1 U525 ( .A1(n462), .A2(n461), .ZN(n463) );
  XOR2_X1 U526 ( .A(KEYINPUT48), .B(n463), .Z(n521) );
  XNOR2_X1 U527 ( .A(KEYINPUT122), .B(n511), .ZN(n464) );
  XNOR2_X1 U528 ( .A(KEYINPUT54), .B(n465), .ZN(n466) );
  NAND2_X1 U529 ( .A1(n466), .A2(n508), .ZN(n563) );
  XNOR2_X1 U530 ( .A(n468), .B(KEYINPUT55), .ZN(n469) );
  NAND2_X1 U531 ( .A1(n558), .A2(n531), .ZN(n471) );
  NOR2_X1 U532 ( .A1(n531), .A2(n544), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n472), .B(KEYINPUT16), .ZN(n474) );
  NAND2_X1 U534 ( .A1(n474), .A2(n473), .ZN(n475) );
  XOR2_X1 U535 ( .A(KEYINPUT102), .B(n475), .Z(n495) );
  NAND2_X1 U536 ( .A1(n476), .A2(n495), .ZN(n485) );
  NOR2_X1 U537 ( .A1(n508), .A2(n485), .ZN(n478) );
  XNOR2_X1 U538 ( .A(KEYINPUT34), .B(KEYINPUT103), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U540 ( .A(G1GAT), .B(n479), .ZN(G1324GAT) );
  NOR2_X1 U541 ( .A1(n511), .A2(n485), .ZN(n480) );
  XOR2_X1 U542 ( .A(G8GAT), .B(n480), .Z(G1325GAT) );
  NOR2_X1 U543 ( .A1(n485), .A2(n513), .ZN(n484) );
  XOR2_X1 U544 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n482) );
  XNOR2_X1 U545 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n481) );
  XNOR2_X1 U546 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U547 ( .A(n484), .B(n483), .ZN(G1326GAT) );
  NOR2_X1 U548 ( .A1(n516), .A2(n485), .ZN(n486) );
  XOR2_X1 U549 ( .A(G22GAT), .B(n486), .Z(G1327GAT) );
  NOR2_X1 U550 ( .A1(n508), .A2(n493), .ZN(n488) );
  XNOR2_X1 U551 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n487) );
  XNOR2_X1 U552 ( .A(n488), .B(n487), .ZN(G1328GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT110), .B(KEYINPUT109), .Z(n490) );
  XNOR2_X1 U554 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n489) );
  XNOR2_X1 U555 ( .A(n490), .B(n489), .ZN(n492) );
  NOR2_X1 U556 ( .A1(n513), .A2(n493), .ZN(n491) );
  XOR2_X1 U557 ( .A(n492), .B(n491), .Z(G1330GAT) );
  NOR2_X1 U558 ( .A1(n516), .A2(n493), .ZN(n494) );
  XOR2_X1 U559 ( .A(G50GAT), .B(n494), .Z(G1331GAT) );
  NOR2_X1 U560 ( .A1(n566), .A2(n540), .ZN(n506) );
  NAND2_X1 U561 ( .A1(n506), .A2(n495), .ZN(n501) );
  NOR2_X1 U562 ( .A1(n508), .A2(n501), .ZN(n496) );
  XOR2_X1 U563 ( .A(G57GAT), .B(n496), .Z(n497) );
  XNOR2_X1 U564 ( .A(KEYINPUT42), .B(n497), .ZN(G1332GAT) );
  NOR2_X1 U565 ( .A1(n511), .A2(n501), .ZN(n498) );
  XOR2_X1 U566 ( .A(G64GAT), .B(n498), .Z(G1333GAT) );
  NOR2_X1 U567 ( .A1(n513), .A2(n501), .ZN(n500) );
  XNOR2_X1 U568 ( .A(G71GAT), .B(KEYINPUT111), .ZN(n499) );
  XNOR2_X1 U569 ( .A(n500), .B(n499), .ZN(G1334GAT) );
  NOR2_X1 U570 ( .A1(n501), .A2(n516), .ZN(n505) );
  XOR2_X1 U571 ( .A(KEYINPUT113), .B(KEYINPUT43), .Z(n503) );
  XNOR2_X1 U572 ( .A(G78GAT), .B(KEYINPUT112), .ZN(n502) );
  XNOR2_X1 U573 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U574 ( .A(n505), .B(n504), .ZN(G1335GAT) );
  NAND2_X1 U575 ( .A1(n507), .A2(n506), .ZN(n515) );
  NOR2_X1 U576 ( .A1(n508), .A2(n515), .ZN(n509) );
  XOR2_X1 U577 ( .A(G85GAT), .B(n509), .Z(n510) );
  XNOR2_X1 U578 ( .A(KEYINPUT114), .B(n510), .ZN(G1336GAT) );
  NOR2_X1 U579 ( .A1(n511), .A2(n515), .ZN(n512) );
  XOR2_X1 U580 ( .A(G92GAT), .B(n512), .Z(G1337GAT) );
  NOR2_X1 U581 ( .A1(n513), .A2(n515), .ZN(n514) );
  XOR2_X1 U582 ( .A(G99GAT), .B(n514), .Z(G1338GAT) );
  NOR2_X1 U583 ( .A1(n516), .A2(n515), .ZN(n518) );
  XNOR2_X1 U584 ( .A(KEYINPUT44), .B(KEYINPUT115), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n519), .ZN(G1339GAT) );
  NOR2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n536) );
  NAND2_X1 U588 ( .A1(n536), .A2(n522), .ZN(n523) );
  XNOR2_X1 U589 ( .A(KEYINPUT118), .B(n523), .ZN(n524) );
  NOR2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n532) );
  NAND2_X1 U591 ( .A1(n550), .A2(n532), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(n526), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT49), .Z(n528) );
  NAND2_X1 U594 ( .A1(n532), .A2(n555), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(G1341GAT) );
  NAND2_X1 U596 ( .A1(n573), .A2(n532), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n529), .B(KEYINPUT50), .ZN(n530) );
  XNOR2_X1 U598 ( .A(G127GAT), .B(n530), .ZN(G1342GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n534) );
  NAND2_X1 U600 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U601 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U602 ( .A(G134GAT), .B(n535), .Z(G1343GAT) );
  NAND2_X1 U603 ( .A1(n536), .A2(n565), .ZN(n547) );
  NOR2_X1 U604 ( .A1(n537), .A2(n547), .ZN(n538) );
  XOR2_X1 U605 ( .A(G141GAT), .B(n538), .Z(n539) );
  XNOR2_X1 U606 ( .A(KEYINPUT120), .B(n539), .ZN(G1344GAT) );
  NOR2_X1 U607 ( .A1(n540), .A2(n547), .ZN(n542) );
  XNOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(n543), .ZN(G1345GAT) );
  NOR2_X1 U611 ( .A1(n544), .A2(n547), .ZN(n546) );
  XNOR2_X1 U612 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G1346GAT) );
  NOR2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U615 ( .A(G162GAT), .B(n549), .Z(G1347GAT) );
  NAND2_X1 U616 ( .A1(n550), .A2(n558), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G169GAT), .B(n551), .ZN(G1348GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n553) );
  XNOR2_X1 U619 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U621 ( .A(KEYINPUT56), .B(n554), .Z(n557) );
  NAND2_X1 U622 ( .A1(n558), .A2(n555), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1349GAT) );
  XOR2_X1 U624 ( .A(G183GAT), .B(KEYINPUT125), .Z(n560) );
  NAND2_X1 U625 ( .A1(n558), .A2(n573), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1350GAT) );
  XNOR2_X1 U627 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(KEYINPUT59), .ZN(n562) );
  XOR2_X1 U629 ( .A(KEYINPUT60), .B(n562), .Z(n568) );
  INV_X1 U630 ( .A(n563), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n575) );
  INV_X1 U632 ( .A(n575), .ZN(n572) );
  NAND2_X1 U633 ( .A1(n572), .A2(n566), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .Z(n571) );
  NAND2_X1 U636 ( .A1(n572), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1353GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n578) );
  XNOR2_X1 U641 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

