//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0 0 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n562, new_n564, new_n565, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n631, new_n633,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1243, new_n1244, new_n1245;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT64), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  OAI211_X1 g035(.A(G137), .B(new_n458), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND4_X1  g039(.A1(new_n464), .A2(KEYINPUT67), .A3(G137), .A4(new_n458), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n458), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n468));
  XNOR2_X1  g043(.A(new_n467), .B(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  XNOR2_X1  g046(.A(new_n471), .B(KEYINPUT66), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OR2_X1    g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g051(.A(G2105), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  AND3_X1   g052(.A1(new_n466), .A2(new_n470), .A3(new_n477), .ZN(G160));
  AOI21_X1  g053(.A(new_n458), .B1(new_n474), .B2(new_n475), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n458), .A2(G112), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n464), .A2(new_n458), .ZN(new_n485));
  INV_X1    g060(.A(G136), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n485), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n488), .A2(KEYINPUT69), .A3(G136), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n483), .B1(new_n487), .B2(new_n489), .ZN(G162));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n459), .C2(new_n460), .ZN(new_n491));
  OR2_X1    g066(.A1(KEYINPUT70), .A2(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(KEYINPUT70), .A2(G114), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n458), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n458), .C1(new_n459), .C2(new_n460), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n464), .A2(new_n499), .A3(G138), .A4(new_n458), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n498), .B2(new_n500), .ZN(G164));
  AND2_X1   g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G62), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT74), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT74), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(new_n510), .A3(G62), .ZN(new_n511));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n506), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n517), .A2(KEYINPUT71), .ZN(new_n518));
  OAI21_X1  g093(.A(G651), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n507), .A2(new_n508), .B1(KEYINPUT6), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n517), .A2(KEYINPUT71), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n520), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n520), .A2(KEYINPUT6), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n527), .B1(new_n502), .B2(new_n503), .ZN(new_n528));
  OAI21_X1  g103(.A(KEYINPUT72), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT73), .B(G88), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n523), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G543), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n532), .B1(KEYINPUT6), .B2(new_n520), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n526), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G50), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n514), .A2(new_n531), .A3(new_n536), .ZN(G303));
  INV_X1    g112(.A(G303), .ZN(G166));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XOR2_X1   g114(.A(new_n539), .B(KEYINPUT7), .Z(new_n540));
  AND3_X1   g115(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n541));
  AOI211_X1 g116(.A(new_n540), .B(new_n541), .C1(G51), .C2(new_n535), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n523), .A2(new_n529), .A3(G89), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n504), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n535), .A2(G52), .B1(new_n548), .B2(G651), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n523), .A2(new_n529), .A3(G90), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  AOI22_X1  g127(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n520), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n523), .A2(new_n529), .A3(G81), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n535), .A2(G43), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n555), .A2(KEYINPUT75), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g132(.A(KEYINPUT75), .B1(new_n555), .B2(new_n556), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(G188));
  XNOR2_X1  g141(.A(KEYINPUT71), .B(KEYINPUT6), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n533), .B1(new_n567), .B2(new_n520), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT9), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n519), .A2(new_n571), .A3(G53), .A4(new_n533), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n523), .A2(new_n529), .A3(G91), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n507), .A2(new_n576), .A3(new_n508), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT76), .B1(new_n502), .B2(new_n503), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AND2_X1   g154(.A1(G78), .A2(G543), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n573), .A2(new_n574), .A3(new_n581), .ZN(G299));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n523), .A2(new_n529), .ZN(new_n584));
  INV_X1    g159(.A(G87), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n523), .A2(new_n529), .A3(KEYINPUT77), .A4(G87), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n509), .A2(G74), .ZN(new_n588));
  AOI22_X1  g163(.A1(G49), .A2(new_n535), .B1(new_n588), .B2(G651), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(G288));
  OAI21_X1  g165(.A(G61), .B1(new_n502), .B2(new_n503), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n520), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(G48), .B2(new_n535), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n523), .A2(new_n529), .A3(G86), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G305));
  AOI22_X1  g171(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(new_n520), .ZN(new_n598));
  OR2_X1    g173(.A1(KEYINPUT78), .A2(G85), .ZN(new_n599));
  NAND2_X1  g174(.A1(KEYINPUT78), .A2(G85), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n523), .A2(new_n529), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n535), .A2(G47), .ZN(new_n602));
  AND2_X1   g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(KEYINPUT79), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n603), .A2(KEYINPUT79), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n598), .B1(new_n605), .B2(new_n606), .ZN(G290));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NOR2_X1   g183(.A1(G301), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n523), .A2(new_n529), .A3(G92), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g187(.A1(new_n523), .A2(new_n529), .A3(KEYINPUT10), .A4(G92), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g189(.A1(new_n535), .A2(G54), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n577), .A2(new_n578), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G66), .ZN(new_n617));
  INV_X1    g192(.A(G79), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n532), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n615), .B1(new_n619), .B2(G651), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n614), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT80), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n614), .A2(new_n620), .A3(KEYINPUT80), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n609), .B1(new_n625), .B2(new_n608), .ZN(G284));
  AOI21_X1  g201(.A(new_n609), .B1(new_n625), .B2(new_n608), .ZN(G321));
  NAND2_X1  g202(.A1(G299), .A2(new_n608), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G168), .B2(new_n608), .ZN(G297));
  OAI21_X1  g204(.A(new_n628), .B1(G168), .B2(new_n608), .ZN(G280));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n625), .B1(new_n631), .B2(G860), .ZN(G148));
  NOR2_X1   g207(.A1(new_n560), .A2(G868), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n625), .A2(new_n631), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(G868), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT81), .Z(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n469), .A2(new_n464), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT13), .ZN(new_n640));
  AOI22_X1  g215(.A1(new_n639), .A2(new_n640), .B1(KEYINPUT82), .B2(G2100), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n640), .B2(new_n639), .ZN(new_n642));
  OR3_X1    g217(.A1(new_n642), .A2(KEYINPUT82), .A3(G2100), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n642), .B1(KEYINPUT82), .B2(G2100), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n479), .A2(G123), .ZN(new_n645));
  OR2_X1    g220(.A1(G99), .A2(G2105), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n646), .B(G2104), .C1(G111), .C2(new_n458), .ZN(new_n647));
  INV_X1    g222(.A(G135), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n645), .B(new_n647), .C1(new_n648), .C2(new_n485), .ZN(new_n649));
  INV_X1    g224(.A(G2096), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n643), .A2(new_n644), .A3(new_n651), .ZN(G156));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n654), .B(new_n655), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2435), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(KEYINPUT14), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(KEYINPUT83), .ZN(new_n664));
  INV_X1    g239(.A(G1341), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT83), .ZN(new_n666));
  NAND4_X1  g241(.A1(new_n661), .A2(new_n666), .A3(KEYINPUT14), .A4(new_n662), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n664), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n665), .B1(new_n664), .B2(new_n667), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n669), .A2(new_n670), .A3(G1348), .ZN(new_n671));
  INV_X1    g246(.A(G1348), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n663), .A2(KEYINPUT83), .ZN(new_n673));
  INV_X1    g248(.A(new_n667), .ZN(new_n674));
  OAI21_X1  g249(.A(G1341), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n672), .B1(new_n675), .B2(new_n668), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n657), .B1(new_n671), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g252(.A(G1348), .B1(new_n669), .B2(new_n670), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n675), .A2(new_n672), .A3(new_n668), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n678), .A2(new_n679), .A3(new_n656), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n677), .A2(G14), .A3(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT84), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g258(.A1(new_n677), .A2(KEYINPUT84), .A3(G14), .A4(new_n680), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(G401));
  INV_X1    g260(.A(KEYINPUT18), .ZN(new_n686));
  XOR2_X1   g261(.A(G2084), .B(G2090), .Z(new_n687));
  XNOR2_X1  g262(.A(G2067), .B(G2678), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(KEYINPUT17), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n687), .A2(new_n688), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n686), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G2072), .B(G2078), .Z(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(new_n689), .B2(KEYINPUT18), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(new_n650), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT85), .B(G2100), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(G227));
  XNOR2_X1  g274(.A(G1971), .B(G1976), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT19), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(G1956), .B(G2474), .Z(new_n703));
  XOR2_X1   g278(.A(G1961), .B(G1966), .Z(new_n704));
  AND2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n703), .A2(new_n704), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  MUX2_X1   g285(.A(new_n710), .B(new_n709), .S(new_n702), .Z(new_n711));
  NOR2_X1   g286(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(G1991), .B(G1996), .Z(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n712), .B(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(G1981), .B(G1986), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT87), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n715), .B(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(G229));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G25), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n488), .A2(G131), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n479), .A2(G119), .ZN(new_n725));
  OR2_X1    g300(.A1(G95), .A2(G2105), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n726), .B(G2104), .C1(G107), .C2(new_n458), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n723), .B1(new_n729), .B2(new_n722), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT35), .B(G1991), .Z(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n730), .B(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G16), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n734), .A2(G24), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G290), .B2(G16), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT88), .B(G1986), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n733), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n734), .A2(G22), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G166), .B2(new_n734), .ZN(new_n740));
  INV_X1    g315(.A(G1971), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(G6), .A2(G16), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G305), .B2(new_n734), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT32), .B(G1981), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n734), .A2(G23), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G288), .B2(G16), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT33), .B(G1976), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n746), .A2(new_n747), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n742), .B(new_n751), .C1(new_n749), .C2(new_n750), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT89), .B(KEYINPUT34), .ZN(new_n753));
  OAI221_X1 g328(.A(new_n738), .B1(new_n736), .B2(new_n737), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n753), .B2(new_n752), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT36), .Z(new_n756));
  NOR2_X1   g331(.A1(G4), .A2(G16), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n625), .B2(G16), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT90), .B(G1348), .Z(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT91), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n758), .B(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT95), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT25), .Z(new_n764));
  AOI22_X1  g339(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n765));
  INV_X1    g340(.A(G139), .ZN(new_n766));
  OAI22_X1  g341(.A1(new_n765), .A2(new_n458), .B1(new_n766), .B2(new_n485), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(new_n722), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n722), .B2(G33), .ZN(new_n771));
  INV_X1    g346(.A(G2072), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(G164), .A2(G29), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G27), .B2(G29), .ZN(new_n775));
  INV_X1    g350(.A(G2078), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n771), .A2(new_n772), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n775), .A2(new_n776), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n773), .A2(new_n777), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n734), .A2(G21), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G168), .B2(new_n734), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1966), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n722), .A2(G32), .ZN(new_n784));
  AOI22_X1  g359(.A1(G141), .A2(new_n488), .B1(new_n469), .B2(G105), .ZN(new_n785));
  NAND3_X1  g360(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT26), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G129), .B2(new_n479), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n784), .B1(new_n790), .B2(new_n722), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT27), .B(G1996), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT31), .B(G11), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT30), .B(G28), .Z(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(G29), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n649), .A2(new_n722), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n796), .B1(new_n798), .B2(KEYINPUT98), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n793), .B(new_n799), .C1(KEYINPUT98), .C2(new_n798), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT24), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n722), .B1(new_n801), .B2(G34), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(KEYINPUT96), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(KEYINPUT96), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n801), .B2(G34), .ZN(new_n805));
  AOI22_X1  g380(.A1(G160), .A2(G29), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT97), .B(G2084), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NOR4_X1   g383(.A1(new_n780), .A2(new_n783), .A3(new_n800), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n734), .A2(G19), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT92), .Z(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n560), .B2(new_n734), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT93), .B(G1341), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n722), .A2(G26), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT28), .Z(new_n816));
  NAND2_X1  g391(.A1(new_n479), .A2(G128), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT94), .ZN(new_n818));
  OAI21_X1  g393(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n819));
  INV_X1    g394(.A(G116), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(G2105), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n488), .B2(G140), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n816), .B1(new_n823), .B2(G29), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(G2067), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n722), .A2(G35), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G162), .B2(new_n722), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT29), .B(G2090), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(G5), .A2(G16), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT99), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(G301), .B2(new_n734), .ZN(new_n832));
  INV_X1    g407(.A(G1961), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT100), .B(KEYINPUT23), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n734), .A2(G20), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G299), .B2(G16), .ZN(new_n839));
  INV_X1    g414(.A(G1956), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n832), .A2(new_n833), .ZN(new_n842));
  NOR4_X1   g417(.A1(new_n825), .A2(new_n835), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  AND4_X1   g418(.A1(new_n761), .A2(new_n809), .A3(new_n814), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n756), .A2(new_n844), .ZN(G150));
  INV_X1    g420(.A(G150), .ZN(G311));
  NAND2_X1  g421(.A1(new_n625), .A2(G559), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT38), .ZN(new_n848));
  NAND2_X1  g423(.A1(G80), .A2(G543), .ZN(new_n849));
  INV_X1    g424(.A(G67), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n504), .B2(new_n850), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n535), .A2(G55), .B1(new_n851), .B2(G651), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n523), .A2(new_n529), .A3(G93), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n559), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n854), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n856), .B(new_n554), .C1(new_n557), .C2(new_n558), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n848), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n860));
  AOI21_X1  g435(.A(G860), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n860), .B2(new_n859), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n854), .A2(G860), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT37), .Z(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(G145));
  XNOR2_X1  g440(.A(G160), .B(new_n649), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G162), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n790), .A2(new_n818), .A3(new_n822), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n823), .A2(new_n789), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(new_n769), .ZN(new_n871));
  XNOR2_X1  g446(.A(G164), .B(KEYINPUT101), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n768), .A2(new_n868), .A3(new_n869), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n872), .B1(new_n871), .B2(new_n873), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT12), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n638), .B(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n488), .A2(G142), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n479), .A2(G130), .ZN(new_n881));
  OR2_X1    g456(.A1(G106), .A2(G2105), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n882), .B(G2104), .C1(G118), .C2(new_n458), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n884), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n639), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n729), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n885), .A2(new_n887), .A3(new_n729), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(KEYINPUT102), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT102), .ZN(new_n892));
  INV_X1    g467(.A(new_n890), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n892), .B1(new_n893), .B2(new_n888), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n867), .B1(new_n877), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n893), .A2(new_n888), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n875), .B2(new_n876), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT103), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n900), .B(new_n897), .C1(new_n875), .C2(new_n876), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n896), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n891), .B(new_n894), .C1(new_n875), .C2(new_n876), .ZN(new_n903));
  INV_X1    g478(.A(new_n876), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n895), .A2(new_n904), .A3(new_n874), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n867), .ZN(new_n907));
  INV_X1    g482(.A(G37), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n902), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g485(.A(new_n858), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n634), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n858), .A2(new_n631), .A3(new_n625), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n915));
  INV_X1    g490(.A(G299), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n621), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n614), .A2(new_n620), .A3(G299), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n915), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n614), .A2(G299), .A3(new_n620), .ZN(new_n922));
  AOI21_X1  g497(.A(G299), .B1(new_n614), .B2(new_n620), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n915), .B(new_n920), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n921), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n917), .A2(new_n927), .A3(new_n918), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n922), .B1(new_n923), .B2(KEYINPUT104), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n920), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n914), .B(KEYINPUT106), .C1(new_n926), .C2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n928), .A2(new_n929), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n912), .A2(new_n933), .A3(new_n913), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n914), .B1(new_n926), .B2(new_n930), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT106), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G288), .ZN(new_n940));
  NAND2_X1  g515(.A1(G290), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n606), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n604), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(G288), .A3(new_n598), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(G303), .B(G305), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n941), .A2(new_n944), .A3(new_n946), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT42), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT42), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n948), .A2(new_n952), .A3(new_n949), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n939), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n935), .A2(new_n954), .A3(new_n938), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n608), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n856), .A2(G868), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT107), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n957), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n954), .B1(new_n935), .B2(new_n938), .ZN(new_n962));
  OAI21_X1  g537(.A(G868), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n964));
  INV_X1    g539(.A(new_n959), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n960), .A2(new_n966), .ZN(G295));
  NAND2_X1  g542(.A1(new_n963), .A2(new_n965), .ZN(G331));
  NAND2_X1  g543(.A1(new_n555), .A2(new_n556), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT75), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n555), .A2(KEYINPUT75), .A3(new_n556), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n856), .B1(new_n973), .B2(new_n554), .ZN(new_n974));
  INV_X1    g549(.A(new_n857), .ZN(new_n975));
  OAI21_X1  g550(.A(G171), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n855), .A2(G301), .A3(new_n857), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(G168), .A3(new_n977), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n855), .A2(G301), .A3(new_n857), .ZN(new_n979));
  AOI21_X1  g554(.A(G301), .B1(new_n855), .B2(new_n857), .ZN(new_n980));
  OAI21_X1  g555(.A(G286), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n978), .B(new_n981), .C1(new_n926), .C2(new_n930), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n979), .A2(new_n980), .A3(G286), .ZN(new_n983));
  AOI21_X1  g558(.A(G168), .B1(new_n976), .B2(new_n977), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n933), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(new_n985), .A3(new_n950), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n986), .A2(new_n908), .ZN(new_n987));
  INV_X1    g562(.A(new_n950), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n932), .A2(new_n920), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n919), .A2(KEYINPUT41), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n981), .A2(new_n978), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n932), .B1(new_n981), .B2(new_n978), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n991), .B1(new_n992), .B2(KEYINPUT108), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT108), .ZN(new_n994));
  AOI211_X1 g569(.A(new_n994), .B(new_n932), .C1(new_n981), .C2(new_n978), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n988), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT43), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n987), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n986), .A2(new_n908), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n950), .B1(new_n982), .B2(new_n985), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT43), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n987), .A2(new_n996), .A3(KEYINPUT43), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n997), .B1(new_n999), .B2(new_n1000), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  MUX2_X1   g580(.A(new_n1002), .B(new_n1005), .S(KEYINPUT44), .Z(G397));
  NAND4_X1  g581(.A1(new_n466), .A2(new_n470), .A3(new_n477), .A4(G40), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n498), .A2(new_n500), .ZN(new_n1010));
  AND2_X1   g585(.A1(KEYINPUT70), .A2(G114), .ZN(new_n1011));
  NOR2_X1   g586(.A1(KEYINPUT70), .A2(G114), .ZN(new_n1012));
  OAI21_X1  g587(.A(G2105), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n495), .ZN(new_n1014));
  AOI22_X1  g589(.A1(G126), .A2(new_n479), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1010), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1384), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1008), .A2(new_n1009), .A3(new_n1018), .ZN(new_n1019));
  OR2_X1    g594(.A1(new_n1019), .A2(G1996), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1020), .B(KEYINPUT46), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1019), .B(KEYINPUT109), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n823), .B(G2067), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1022), .B1(new_n789), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1025), .B(KEYINPUT47), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1022), .A2(G1996), .A3(new_n789), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n1020), .A2(new_n789), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n729), .A2(new_n731), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n728), .A2(new_n732), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1022), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  NOR3_X1   g609(.A1(G290), .A2(G1986), .A3(new_n1019), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n1035), .B(KEYINPUT48), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n823), .A2(G2067), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1022), .ZN(new_n1039));
  OAI221_X1 g614(.A(new_n1026), .B1(new_n1034), .B2(new_n1036), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g615(.A(new_n1040), .B(KEYINPUT126), .Z(new_n1041));
  INV_X1    g616(.A(KEYINPUT63), .ZN(new_n1042));
  AOI21_X1  g617(.A(G1384), .B1(new_n1010), .B2(new_n1015), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT114), .B1(new_n1045), .B2(new_n1007), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1008), .B(new_n1047), .C1(new_n1044), .C2(new_n1043), .ZN(new_n1048));
  INV_X1    g623(.A(G2090), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1046), .A2(new_n1048), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1009), .B1(G164), .B2(G1384), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1043), .A2(KEYINPUT45), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(new_n1008), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n741), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(G8), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(KEYINPUT110), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(KEYINPUT110), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  AOI211_X1 g636(.A(new_n1059), .B(new_n1061), .C1(G303), .C2(G8), .ZN(new_n1062));
  NAND4_X1  g637(.A1(G303), .A2(KEYINPUT110), .A3(new_n1058), .A4(G8), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1057), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G8), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1068), .B1(new_n1008), .B2(new_n1043), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT111), .ZN(new_n1070));
  OAI21_X1  g645(.A(G1981), .B1(new_n593), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(G305), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n594), .A2(new_n595), .A3(new_n1071), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT49), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1069), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n594), .A2(new_n595), .A3(new_n1071), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1071), .B1(new_n594), .B2(new_n595), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1076), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT112), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT112), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1075), .A2(new_n1082), .A3(new_n1076), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1077), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G1976), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT52), .B1(G288), .B2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n586), .A2(G1976), .A3(new_n587), .A4(new_n589), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1086), .A2(new_n1069), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1089), .B1(new_n1069), .B2(new_n1087), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1084), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1007), .B1(new_n1018), .B2(KEYINPUT50), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1094), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1068), .B1(new_n1055), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n1065), .ZN(new_n1097));
  INV_X1    g672(.A(G1966), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1054), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G2084), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1094), .A2(new_n1100), .A3(new_n1050), .ZN(new_n1101));
  AOI211_X1 g676(.A(new_n1068), .B(G286), .C1(new_n1099), .C2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1067), .A2(new_n1093), .A3(new_n1097), .A4(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1055), .A2(new_n1095), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(G8), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT115), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1059), .B1(G303), .B2(G8), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n1060), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1106), .B1(new_n1108), .B2(new_n1063), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1096), .B1(new_n1065), .B2(new_n1106), .ZN(new_n1111));
  AND4_X1   g686(.A1(KEYINPUT63), .A2(new_n1110), .A3(new_n1102), .A4(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT113), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1084), .B2(new_n1092), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1077), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1087), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1008), .A2(new_n1043), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(G8), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1090), .B1(new_n1121), .B2(new_n1086), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1117), .A2(new_n1122), .A3(KEYINPUT113), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1114), .A2(new_n1123), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1042), .A2(new_n1103), .B1(new_n1112), .B2(new_n1124), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1084), .A2(G1976), .A3(G288), .ZN(new_n1126));
  NOR2_X1   g701(.A1(G305), .A2(G1981), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1069), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1114), .A2(new_n1123), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1128), .B1(new_n1129), .B2(new_n1097), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1125), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1097), .A2(new_n1117), .A3(new_n1122), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1065), .B1(new_n1056), .B2(G8), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT124), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1067), .A2(new_n1093), .A3(new_n1135), .A4(new_n1097), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1052), .A2(new_n1053), .A3(new_n776), .A4(new_n1008), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT53), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1094), .A2(new_n1050), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1140), .A2(KEYINPUT123), .B1(new_n833), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1138), .A2(new_n1143), .A3(new_n1139), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1138), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1007), .B1(KEYINPUT45), .B2(new_n1043), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1148), .A2(KEYINPUT122), .A3(new_n776), .A4(new_n1052), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1147), .A2(KEYINPUT53), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(G301), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1068), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1099), .A2(G168), .A3(new_n1101), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(G8), .ZN(new_n1154));
  AOI21_X1  g729(.A(G168), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1155));
  OAI221_X1 g730(.A(KEYINPUT51), .B1(KEYINPUT121), .B2(new_n1152), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(KEYINPUT51), .B1(new_n1152), .B2(KEYINPUT121), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1157), .A2(G8), .A3(new_n1153), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT62), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1156), .A2(new_n1161), .A3(new_n1158), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1137), .A2(new_n1151), .A3(new_n1160), .A4(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT57), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT116), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n573), .A2(new_n574), .A3(new_n581), .A4(new_n1165), .ZN(new_n1166));
  OR2_X1    g741(.A1(new_n1164), .A2(KEYINPUT116), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1166), .B(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1050), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1008), .B1(new_n1044), .B2(new_n1043), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1170), .B1(new_n1171), .B2(KEYINPUT114), .ZN(new_n1172));
  AOI21_X1  g747(.A(G1956), .B1(new_n1172), .B2(new_n1048), .ZN(new_n1173));
  XNOR2_X1  g748(.A(KEYINPUT56), .B(G2072), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1148), .A2(new_n1174), .A3(new_n1052), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(KEYINPUT117), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT117), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1148), .A2(new_n1177), .A3(new_n1174), .A4(new_n1052), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1169), .B1(new_n1173), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n625), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1119), .A2(G2067), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1182), .B1(new_n672), .B2(new_n1141), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1180), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1046), .A2(new_n1050), .A3(new_n1048), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(new_n840), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1186), .A2(new_n1168), .A3(new_n1178), .A4(new_n1176), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1180), .A2(KEYINPUT61), .A3(new_n1187), .ZN(new_n1189));
  AOI21_X1  g764(.A(KEYINPUT61), .B1(new_n1180), .B2(new_n1187), .ZN(new_n1190));
  NAND2_X1  g765(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n973), .A2(new_n554), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1192), .ZN(new_n1193));
  OR2_X1    g768(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1194));
  XOR2_X1   g769(.A(KEYINPUT58), .B(G1341), .Z(new_n1195));
  NAND2_X1  g770(.A1(new_n1119), .A2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1196), .B1(new_n1054), .B2(G1996), .ZN(new_n1197));
  AND3_X1   g772(.A1(new_n1193), .A2(new_n1194), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1194), .B1(new_n1193), .B2(new_n1197), .ZN(new_n1199));
  OR2_X1    g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NOR3_X1   g775(.A1(new_n1189), .A2(new_n1190), .A3(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT119), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n625), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n623), .A2(KEYINPUT119), .A3(new_n624), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1203), .A2(new_n1183), .A3(KEYINPUT60), .A4(new_n1204), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1171), .A2(new_n1170), .ZN(new_n1206));
  OAI22_X1  g781(.A1(new_n1206), .A2(G1348), .B1(G2067), .B2(new_n1119), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT60), .ZN(new_n1208));
  OAI211_X1 g783(.A(new_n1181), .B(KEYINPUT119), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1205), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT120), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND4_X1  g788(.A1(new_n1205), .A2(new_n1209), .A3(KEYINPUT120), .A4(new_n1210), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1188), .B1(new_n1201), .B2(new_n1215), .ZN(new_n1216));
  NAND4_X1  g791(.A1(new_n1142), .A2(G301), .A3(new_n1144), .A4(new_n1150), .ZN(new_n1217));
  AND2_X1   g792(.A1(new_n1217), .A2(KEYINPUT54), .ZN(new_n1218));
  OR2_X1    g793(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1142), .A2(new_n1144), .A3(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1220), .A2(G171), .ZN(new_n1221));
  AOI22_X1  g796(.A1(new_n1218), .A2(new_n1221), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT54), .ZN(new_n1223));
  NOR2_X1   g798(.A1(new_n1220), .A2(G171), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1223), .B1(new_n1151), .B2(new_n1224), .ZN(new_n1225));
  NAND4_X1  g800(.A1(new_n1222), .A2(new_n1225), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1226));
  OAI211_X1 g801(.A(new_n1131), .B(new_n1163), .C1(new_n1216), .C2(new_n1226), .ZN(new_n1227));
  INV_X1    g802(.A(new_n1019), .ZN(new_n1228));
  XNOR2_X1  g803(.A(G290), .B(G1986), .ZN(new_n1229));
  AOI21_X1  g804(.A(new_n1034), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  AND3_X1   g805(.A1(new_n1227), .A2(KEYINPUT125), .A3(new_n1230), .ZN(new_n1231));
  AOI21_X1  g806(.A(KEYINPUT125), .B1(new_n1227), .B2(new_n1230), .ZN(new_n1232));
  OAI21_X1  g807(.A(new_n1041), .B1(new_n1231), .B2(new_n1232), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g808(.A1(new_n720), .A2(G319), .A3(new_n698), .ZN(new_n1235));
  AOI21_X1  g809(.A(new_n1235), .B1(new_n683), .B2(new_n684), .ZN(new_n1236));
  NAND2_X1  g810(.A1(new_n909), .A2(new_n1236), .ZN(new_n1237));
  AOI211_X1 g811(.A(KEYINPUT127), .B(new_n1237), .C1(new_n998), .C2(new_n1001), .ZN(new_n1238));
  INV_X1    g812(.A(KEYINPUT127), .ZN(new_n1239));
  INV_X1    g813(.A(new_n1237), .ZN(new_n1240));
  AOI21_X1  g814(.A(new_n1239), .B1(new_n1002), .B2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g815(.A1(new_n1238), .A2(new_n1241), .ZN(G308));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n1240), .ZN(new_n1243));
  NAND2_X1  g817(.A1(new_n1243), .A2(KEYINPUT127), .ZN(new_n1244));
  NAND3_X1  g818(.A1(new_n1002), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1245));
  NAND2_X1  g819(.A1(new_n1244), .A2(new_n1245), .ZN(G225));
endmodule


