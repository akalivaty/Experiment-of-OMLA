//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n548, new_n549, new_n550, new_n551, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n568, new_n569, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n631, new_n633,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g041(.A(G137), .B1(new_n462), .B2(new_n463), .ZN(new_n467));
  NAND2_X1  g042(.A1(G101), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(G160));
  NOR2_X1   g045(.A1(new_n462), .A2(new_n463), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G136), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n471), .A2(new_n461), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G162));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n480));
  NAND2_X1  g055(.A1(G126), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n482), .B1(new_n462), .B2(new_n463), .ZN(new_n483));
  INV_X1    g058(.A(G102), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(new_n461), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n485), .A2(new_n487), .A3(G2104), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n483), .A2(new_n488), .A3(KEYINPUT66), .ZN(new_n489));
  AOI21_X1  g064(.A(KEYINPUT66), .B1(new_n483), .B2(new_n488), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(G138), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OR2_X1    g069(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .A3(G138), .A4(new_n461), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n480), .B1(new_n491), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT66), .ZN(new_n501));
  AND3_X1   g076(.A1(new_n485), .A2(new_n487), .A3(G2104), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n481), .B1(new_n495), .B2(new_n496), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n483), .A2(new_n488), .A3(KEYINPUT66), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n494), .A2(new_n498), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT67), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n500), .A2(new_n508), .ZN(G164));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G50), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G651), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  OAI211_X1 g093(.A(new_n514), .B(new_n516), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n511), .A2(new_n512), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  OR2_X1    g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G62), .ZN(new_n526));
  NAND2_X1  g101(.A1(G75), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n522), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT68), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n522), .A2(KEYINPUT68), .A3(new_n529), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(G166));
  NAND2_X1  g109(.A1(new_n511), .A2(KEYINPUT69), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n514), .A2(new_n516), .A3(G543), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT69), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n540), .A2(G51), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT7), .ZN(new_n544));
  INV_X1    g119(.A(G89), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n542), .B(new_n544), .C1(new_n545), .C2(new_n519), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n541), .A2(new_n546), .ZN(G168));
  AND3_X1   g122(.A1(new_n535), .A2(new_n538), .A3(G52), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G90), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n549), .A2(new_n513), .B1(new_n550), .B2(new_n519), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(G171));
  AND2_X1   g127(.A1(G68), .A2(G543), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n525), .B2(G56), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n554), .A2(new_n513), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT70), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n540), .A2(G43), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n554), .A2(new_n513), .ZN(new_n558));
  INV_X1    g133(.A(new_n519), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n558), .A2(KEYINPUT70), .B1(G81), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT71), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT71), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n557), .A2(new_n563), .A3(new_n560), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  NAND4_X1  g141(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(G188));
  INV_X1    g145(.A(KEYINPUT73), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n519), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n525), .A2(new_n510), .A3(KEYINPUT73), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n572), .A2(G91), .A3(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(KEYINPUT72), .ZN(new_n576));
  AND2_X1   g151(.A1(G53), .A2(G543), .ZN(new_n577));
  AND3_X1   g152(.A1(new_n510), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n576), .B1(new_n510), .B2(new_n577), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n525), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n523), .A2(KEYINPUT74), .A3(new_n524), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n584), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n574), .B(new_n580), .C1(new_n585), .C2(new_n513), .ZN(G299));
  INV_X1    g161(.A(G171), .ZN(G301));
  OR2_X1    g162(.A1(new_n541), .A2(new_n546), .ZN(G286));
  INV_X1    g163(.A(G166), .ZN(G303));
  NAND3_X1  g164(.A1(new_n572), .A2(G87), .A3(new_n573), .ZN(new_n590));
  INV_X1    g165(.A(G74), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n523), .A2(new_n591), .A3(new_n524), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n536), .A2(G49), .B1(new_n592), .B2(G651), .ZN(new_n593));
  AND3_X1   g168(.A1(new_n590), .A2(KEYINPUT75), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g169(.A(KEYINPUT75), .B1(new_n590), .B2(new_n593), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n594), .A2(new_n595), .ZN(G288));
  AND2_X1   g171(.A1(G48), .A2(G543), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n514), .A2(new_n516), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT77), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n510), .A2(KEYINPUT77), .A3(new_n597), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n525), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n602));
  OAI211_X1 g177(.A(new_n600), .B(new_n601), .C1(new_n602), .C2(new_n513), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n572), .A2(G86), .A3(new_n573), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT76), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n572), .A2(new_n573), .A3(KEYINPUT76), .A4(G86), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n603), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G305));
  NAND2_X1  g184(.A1(new_n559), .A2(G85), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n611));
  INV_X1    g186(.A(G47), .ZN(new_n612));
  OAI221_X1 g187(.A(new_n610), .B1(new_n513), .B2(new_n611), .C1(new_n539), .C2(new_n612), .ZN(G290));
  NAND2_X1  g188(.A1(G301), .A2(G868), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n584), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G54), .ZN(new_n616));
  OAI22_X1  g191(.A1(new_n615), .A2(new_n513), .B1(new_n539), .B2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n572), .A2(G92), .A3(new_n573), .ZN(new_n620));
  XOR2_X1   g195(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n614), .B1(new_n624), .B2(G868), .ZN(G284));
  OAI21_X1  g200(.A(new_n614), .B1(new_n624), .B2(G868), .ZN(G321));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(G299), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G168), .B2(new_n627), .ZN(G297));
  OAI21_X1  g204(.A(new_n628), .B1(G168), .B2(new_n627), .ZN(G280));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n624), .B1(new_n631), .B2(G860), .ZN(G148));
  NAND2_X1  g207(.A1(new_n565), .A2(new_n627), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n624), .A2(new_n631), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(new_n627), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT11), .Z(G282));
  INV_X1    g211(.A(new_n635), .ZN(G323));
  NAND2_X1  g212(.A1(new_n472), .A2(G2104), .ZN(new_n638));
  XOR2_X1   g213(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT13), .Z(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(G2100), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(G2100), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n472), .A2(G135), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n474), .A2(G123), .ZN(new_n645));
  NOR2_X1   g220(.A1(G99), .A2(G2105), .ZN(new_n646));
  OAI21_X1  g221(.A(G2104), .B1(new_n461), .B2(G111), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n644), .B(new_n645), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(G2096), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n642), .A2(new_n643), .A3(new_n650), .ZN(G156));
  XNOR2_X1  g226(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G1341), .B(G1348), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT82), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n656), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2427), .B(G2438), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2430), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT15), .B(G2435), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  AND3_X1   g239(.A1(new_n663), .A2(new_n664), .A3(KEYINPUT14), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n659), .A2(new_n665), .ZN(new_n667));
  AND3_X1   g242(.A1(new_n666), .A2(G14), .A3(new_n667), .ZN(G401));
  XNOR2_X1  g243(.A(G2072), .B(G2078), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT17), .Z(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(new_n671), .B2(new_n669), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT83), .Z(new_n678));
  NAND3_X1  g253(.A1(new_n674), .A2(new_n671), .A3(new_n669), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT18), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n675), .A2(new_n671), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n680), .B1(new_n670), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(new_n649), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G2100), .ZN(G227));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1956), .B(G2474), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1961), .B(G1966), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NOR3_X1   g266(.A1(new_n687), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n687), .A2(new_n690), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT20), .Z(new_n694));
  AOI211_X1 g269(.A(new_n692), .B(new_n694), .C1(new_n687), .C2(new_n691), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  INV_X1    g274(.A(G1981), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n698), .B(new_n701), .ZN(G229));
  NAND2_X1  g277(.A1(G168), .A2(G16), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT92), .Z(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G16), .B2(G21), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1966), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n472), .A2(G141), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n474), .A2(G129), .ZN(new_n708));
  NAND3_X1  g283(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT26), .Z(new_n710));
  NAND3_X1  g285(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n711));
  NAND4_X1  g286(.A1(new_n707), .A2(new_n708), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  MUX2_X1   g287(.A(G32), .B(new_n712), .S(G29), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT27), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G1996), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n565), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n716), .B2(G19), .ZN(new_n718));
  INV_X1    g293(.A(G1341), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT84), .B(G29), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n722), .A2(G35), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G162), .B2(new_n722), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT29), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n725), .A2(G2090), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT31), .B(G11), .Z(new_n727));
  NOR2_X1   g302(.A1(new_n648), .A2(new_n721), .ZN(new_n728));
  INV_X1    g303(.A(G28), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n729), .A2(KEYINPUT30), .ZN(new_n730));
  AOI21_X1  g305(.A(G29), .B1(new_n729), .B2(KEYINPUT30), .ZN(new_n731));
  AOI211_X1 g306(.A(new_n727), .B(new_n728), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT24), .B(G34), .ZN(new_n733));
  AOI22_X1  g308(.A1(G160), .A2(G29), .B1(new_n721), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G2084), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(G2084), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n732), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n716), .A2(G5), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G171), .B2(new_n716), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1961), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n472), .A2(G140), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n474), .A2(G128), .ZN(new_n742));
  OR2_X1    g317(.A1(G104), .A2(G2105), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n743), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n721), .A2(G26), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT28), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G2067), .ZN(new_n750));
  NOR4_X1   g325(.A1(new_n726), .A2(new_n737), .A3(new_n740), .A4(new_n750), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n706), .A2(new_n715), .A3(new_n720), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(G115), .A2(G2104), .ZN(new_n753));
  INV_X1    g328(.A(G127), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n471), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n461), .B1(new_n755), .B2(KEYINPUT90), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(KEYINPUT90), .B2(new_n755), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT25), .ZN(new_n758));
  NAND2_X1  g333(.A1(G103), .A2(G2104), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(G2105), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n461), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n472), .A2(G139), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  MUX2_X1   g338(.A(G33), .B(new_n763), .S(G29), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT91), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(G2072), .Z(new_n766));
  NOR2_X1   g341(.A1(new_n722), .A2(G27), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G164), .B2(new_n722), .ZN(new_n768));
  INV_X1    g343(.A(G2078), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n718), .B2(new_n719), .ZN(new_n771));
  NOR3_X1   g346(.A1(new_n752), .A2(new_n766), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n716), .A2(G4), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n624), .B2(new_n716), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT89), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1348), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n716), .A2(G20), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT23), .ZN(new_n778));
  INV_X1    g353(.A(G299), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(new_n716), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT93), .Z(new_n781));
  AOI22_X1  g356(.A1(new_n781), .A2(G1956), .B1(new_n725), .B2(G2090), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G1956), .B2(new_n781), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT94), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n772), .A2(new_n776), .A3(new_n784), .ZN(new_n785));
  MUX2_X1   g360(.A(G24), .B(G290), .S(G16), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(G1986), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n722), .A2(G25), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n472), .A2(G131), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n474), .A2(G119), .ZN(new_n790));
  OR2_X1    g365(.A1(G95), .A2(G2105), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n791), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n789), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n788), .B1(new_n794), .B2(new_n722), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT35), .B(G1991), .Z(new_n796));
  XOR2_X1   g371(.A(new_n795), .B(new_n796), .Z(new_n797));
  NOR2_X1   g372(.A1(new_n786), .A2(G1986), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n716), .A2(G22), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT87), .Z(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G166), .B2(new_n716), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1971), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n716), .A2(G23), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n590), .A2(new_n593), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(KEYINPUT86), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT86), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n590), .A2(new_n807), .A3(new_n593), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n804), .B1(new_n809), .B2(G16), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT33), .B(G1976), .Z(new_n812));
  AOI21_X1  g387(.A(new_n803), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n716), .A2(G6), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n608), .B2(new_n716), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT32), .B(G1981), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n811), .A2(new_n812), .ZN(new_n818));
  AND3_X1   g393(.A1(new_n813), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT85), .B(KEYINPUT34), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n787), .B(new_n799), .C1(new_n820), .C2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT88), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n820), .A2(new_n822), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n826), .A2(KEYINPUT36), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(KEYINPUT36), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n785), .B1(new_n827), .B2(new_n828), .ZN(G311));
  INV_X1    g404(.A(G311), .ZN(G150));
  NAND2_X1  g405(.A1(new_n562), .A2(new_n564), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n559), .A2(G93), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n833));
  INV_X1    g408(.A(G55), .ZN(new_n834));
  OAI221_X1 g409(.A(new_n832), .B1(new_n513), .B2(new_n833), .C1(new_n539), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n561), .B2(new_n835), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT38), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n624), .A2(G559), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n841), .A2(new_n842), .A3(G860), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n835), .A2(G860), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT37), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n843), .A2(new_n845), .ZN(G145));
  XNOR2_X1  g421(.A(new_n478), .B(G160), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT95), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n648), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n712), .B(new_n745), .ZN(new_n850));
  INV_X1    g425(.A(G2104), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(new_n486), .B2(G2105), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n497), .A2(new_n482), .B1(new_n852), .B2(new_n485), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n853), .A2(new_n494), .A3(new_n498), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n850), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT96), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n855), .A2(new_n856), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n763), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT97), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n763), .B2(new_n855), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n859), .A2(new_n860), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n474), .A2(G130), .ZN(new_n866));
  NOR2_X1   g441(.A1(G106), .A2(G2105), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(G142), .B2(new_n472), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n794), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n640), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n849), .B1(new_n865), .B2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(KEYINPUT98), .ZN(new_n874));
  OR3_X1    g449(.A1(new_n862), .A2(new_n863), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(G37), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n865), .A2(new_n874), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n875), .ZN(new_n878));
  AOI21_X1  g453(.A(KEYINPUT99), .B1(new_n878), .B2(new_n849), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n880));
  INV_X1    g455(.A(new_n849), .ZN(new_n881));
  AOI211_X1 g456(.A(new_n880), .B(new_n881), .C1(new_n877), .C2(new_n875), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n876), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g459(.A(new_n837), .B(new_n634), .Z(new_n885));
  NOR2_X1   g460(.A1(new_n624), .A2(G299), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n624), .A2(G299), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT100), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n885), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(KEYINPUT101), .Z(new_n892));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n893));
  INV_X1    g468(.A(new_n888), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n893), .B1(new_n894), .B2(new_n886), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n895), .A2(KEYINPUT102), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n890), .A2(KEYINPUT41), .A3(new_n887), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(KEYINPUT102), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n885), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n892), .A2(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(G290), .B(KEYINPUT103), .Z(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(new_n809), .ZN(new_n903));
  XNOR2_X1  g478(.A(G166), .B(G305), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n904), .A2(KEYINPUT104), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(KEYINPUT104), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n907), .B1(new_n906), .B2(new_n903), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT105), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n911), .B1(new_n910), .B2(new_n908), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n901), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n901), .A2(new_n912), .ZN(new_n915));
  OAI21_X1  g490(.A(G868), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n835), .A2(new_n627), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(G295));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n917), .ZN(G331));
  NAND2_X1  g494(.A1(G286), .A2(G171), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT107), .ZN(new_n921));
  NAND2_X1  g496(.A1(G168), .A2(G301), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT106), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  XOR2_X1   g499(.A(new_n924), .B(new_n837), .Z(new_n925));
  AOI21_X1  g500(.A(KEYINPUT41), .B1(new_n890), .B2(new_n887), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n894), .A2(new_n893), .A3(new_n886), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n925), .B(KEYINPUT108), .C1(new_n926), .C2(new_n927), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n890), .A2(new_n887), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n924), .B(new_n837), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT109), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n932), .A2(new_n933), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT109), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n930), .A2(new_n931), .A3(new_n935), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n909), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n934), .B1(new_n899), .B2(new_n925), .ZN(new_n942));
  INV_X1    g517(.A(new_n909), .ZN(new_n943));
  AOI21_X1  g518(.A(G37), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n940), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n899), .A2(new_n925), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n909), .B1(new_n946), .B2(new_n934), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n945), .B1(new_n948), .B2(new_n941), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n940), .A2(KEYINPUT43), .A3(new_n944), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT43), .B1(new_n944), .B2(new_n947), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT44), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n951), .A2(new_n954), .ZN(G397));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n956));
  INV_X1    g531(.A(G1384), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n854), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n956), .B1(new_n958), .B2(KEYINPUT110), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n959), .B1(KEYINPUT110), .B2(new_n958), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n464), .A2(new_n465), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(G2105), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n467), .A2(new_n468), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n461), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n962), .A2(new_n964), .A3(G40), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n960), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G1996), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT46), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT125), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n968), .A2(new_n969), .ZN(new_n972));
  INV_X1    g547(.A(G2067), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n745), .B(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n966), .B1(new_n712), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT126), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n971), .A2(new_n972), .A3(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT47), .ZN(new_n979));
  NOR2_X1   g554(.A1(G290), .A2(G1986), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n966), .A2(new_n980), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n981), .B(KEYINPUT48), .Z(new_n982));
  XNOR2_X1  g557(.A(new_n712), .B(G1996), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n966), .B1(new_n975), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT111), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n793), .B(new_n796), .Z(new_n986));
  AND2_X1   g561(.A1(new_n966), .A2(new_n986), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n982), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n794), .A2(new_n796), .ZN(new_n989));
  OAI22_X1  g564(.A1(new_n985), .A2(new_n989), .B1(G2067), .B2(new_n745), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n988), .B1(new_n966), .B2(new_n990), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n979), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n806), .A2(G1976), .A3(new_n808), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n854), .A2(new_n957), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n962), .A2(new_n964), .A3(G40), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n994), .B(G8), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(G160), .A2(new_n854), .A3(G40), .A4(new_n957), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n994), .B1(new_n999), .B2(G8), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n993), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT52), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n995), .A2(new_n996), .ZN(new_n1003));
  INV_X1    g578(.A(G8), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT112), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n997), .ZN(new_n1006));
  INV_X1    g581(.A(G1976), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT52), .B1(G288), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1008), .A3(new_n993), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1002), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n998), .A2(new_n1000), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT49), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n600), .A2(new_n601), .ZN(new_n1013));
  OAI21_X1  g588(.A(G61), .B1(new_n517), .B2(new_n518), .ZN(new_n1014));
  NAND2_X1  g589(.A1(G73), .A2(G543), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n513), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n559), .A2(G86), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n700), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1019), .B1(new_n608), .B2(new_n700), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1012), .B1(new_n1020), .B2(KEYINPUT113), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n1022));
  AOI211_X1 g597(.A(G1981), .B(new_n603), .C1(new_n606), .C2(new_n607), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1022), .B(KEYINPUT49), .C1(new_n1023), .C2(new_n1019), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1011), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1010), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n500), .A2(new_n1027), .A3(new_n957), .A4(new_n508), .ZN(new_n1028));
  INV_X1    g603(.A(G2090), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n996), .B1(new_n995), .B2(KEYINPUT50), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n965), .B1(new_n995), .B2(new_n956), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n500), .A2(new_n957), .A3(new_n508), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1032), .B1(new_n1033), .B2(new_n956), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1031), .B1(new_n1034), .B2(G1971), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(G8), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n532), .A2(new_n533), .A3(G8), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1037), .B(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1034), .A2(G1971), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n965), .B1(new_n995), .B2(KEYINPUT50), .ZN(new_n1043));
  AOI211_X1 g618(.A(G2090), .B(new_n1043), .C1(new_n1033), .C2(KEYINPUT50), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1039), .B(G8), .C1(new_n1042), .C2(new_n1044), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1026), .A2(new_n1041), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(G286), .A2(G8), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1043), .B1(new_n1033), .B2(KEYINPUT50), .ZN(new_n1048));
  INV_X1    g623(.A(G2084), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n957), .A4(new_n508), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n996), .B1(new_n995), .B2(new_n956), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G1966), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1048), .A2(new_n1049), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g629(.A(KEYINPUT51), .B(new_n1047), .C1(new_n1054), .C2(new_n1004), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1033), .A2(KEYINPUT50), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1043), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1049), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1056), .B(G8), .C1(new_n1061), .C2(G286), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT121), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1047), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1063), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  AOI211_X1 g640(.A(KEYINPUT121), .B(new_n1047), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1055), .B(new_n1062), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1034), .A2(new_n769), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1070));
  INV_X1    g645(.A(G1961), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1068), .A2(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT122), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n1052), .B2(G2078), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1050), .A2(KEYINPUT122), .A3(new_n769), .A4(new_n1051), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(KEYINPUT53), .A3(new_n1075), .ZN(new_n1076));
  XOR2_X1   g651(.A(G171), .B(KEYINPUT54), .Z(new_n1077));
  NAND3_X1  g652(.A1(new_n1072), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  AOI211_X1 g653(.A(G2078), .B(new_n1032), .C1(new_n1033), .C2(new_n956), .ZN(new_n1079));
  OAI22_X1  g654(.A1(new_n1079), .A2(KEYINPUT53), .B1(G1961), .B2(new_n1048), .ZN(new_n1080));
  NOR4_X1   g655(.A1(new_n960), .A2(new_n1069), .A3(G2078), .A4(new_n1032), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1078), .B1(new_n1082), .B2(new_n1077), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1046), .A2(new_n1067), .A3(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT56), .B(G2072), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1034), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1087));
  INV_X1    g662(.A(G1956), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n1092));
  INV_X1    g667(.A(new_n583), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT74), .B1(new_n523), .B2(new_n524), .ZN(new_n1094));
  OAI21_X1  g669(.A(G65), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(G78), .A2(G543), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n513), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n580), .A2(new_n574), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1092), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT57), .B1(G299), .B2(new_n1092), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1091), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1104));
  NAND3_X1  g679(.A1(G299), .A2(new_n1092), .A3(KEYINPUT57), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1104), .A2(new_n1105), .A3(KEYINPUT117), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1090), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1003), .A2(new_n973), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n1048), .B2(G1348), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n624), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1086), .A2(new_n1089), .A3(new_n1113), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1085), .ZN(new_n1117));
  AOI211_X1 g692(.A(new_n1117), .B(new_n1032), .C1(new_n1033), .C2(new_n956), .ZN(new_n1118));
  AOI21_X1  g693(.A(G1956), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1119));
  OAI22_X1  g694(.A1(new_n1118), .A2(new_n1119), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1114), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT61), .ZN(new_n1122));
  NAND2_X1  g697(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT58), .B(G1341), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1003), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1126), .B1(new_n1034), .B2(new_n967), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1124), .B1(new_n1127), .B2(new_n831), .ZN(new_n1128));
  AOI211_X1 g703(.A(G1996), .B(new_n1032), .C1(new_n1033), .C2(new_n956), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n565), .B(new_n1123), .C1(new_n1129), .C2(new_n1126), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1121), .A2(new_n1122), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1114), .A2(KEYINPUT119), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1086), .A2(new_n1089), .A3(new_n1133), .A4(new_n1113), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1132), .A2(new_n1108), .A3(KEYINPUT61), .A4(new_n1134), .ZN(new_n1135));
  OR2_X1    g710(.A1(new_n1048), .A2(G1348), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1136), .A2(KEYINPUT120), .A3(KEYINPUT60), .A4(new_n1109), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT60), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1138), .B1(new_n1110), .B2(new_n1139), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1137), .A2(new_n624), .A3(new_n1140), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1138), .B(new_n623), .C1(new_n1110), .C2(new_n1139), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1110), .A2(new_n1139), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1131), .B(new_n1135), .C1(new_n1141), .C2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1084), .B1(new_n1116), .B2(new_n1145), .ZN(new_n1146));
  AOI211_X1 g721(.A(new_n1004), .B(G286), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1026), .A2(new_n1041), .A3(new_n1045), .A4(new_n1147), .ZN(new_n1148));
  XOR2_X1   g723(.A(KEYINPUT114), .B(KEYINPUT63), .Z(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1010), .A2(new_n1025), .A3(new_n1151), .ZN(new_n1152));
  OAI221_X1 g727(.A(G8), .B1(new_n1042), .B2(new_n1044), .C1(KEYINPUT115), .C2(new_n1039), .ZN(new_n1153));
  OAI21_X1  g728(.A(G8), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT115), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1154), .A2(new_n1155), .A3(new_n1040), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1152), .A2(new_n1153), .A3(new_n1156), .A4(new_n1147), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1150), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1045), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n1026), .ZN(new_n1160));
  NOR2_X1   g735(.A1(G288), .A2(G1976), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1021), .A2(new_n1024), .A3(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1006), .B1(new_n1162), .B2(new_n1023), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1158), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT123), .B1(new_n1146), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT123), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1164), .B1(new_n1150), .B2(new_n1157), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1135), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1137), .A2(new_n624), .A3(new_n1140), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1173), .A2(new_n1143), .A3(new_n1142), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1115), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g750(.A(new_n1168), .B(new_n1169), .C1(new_n1175), .C2(new_n1084), .ZN(new_n1176));
  OR2_X1    g751(.A1(new_n1067), .A2(KEYINPUT62), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1067), .A2(KEYINPUT62), .ZN(new_n1178));
  AOI21_X1  g753(.A(G301), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1177), .A2(new_n1046), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1167), .A2(new_n1176), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n1182));
  XNOR2_X1  g757(.A(G290), .B(G1986), .ZN(new_n1183));
  AOI211_X1 g758(.A(new_n987), .B(new_n985), .C1(new_n966), .C2(new_n1183), .ZN(new_n1184));
  AND3_X1   g759(.A1(new_n1181), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1182), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n992), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(KEYINPUT127), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n1189));
  OAI211_X1 g764(.A(new_n1189), .B(new_n992), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1188), .A2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g766(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1193));
  AND3_X1   g767(.A1(new_n949), .A2(new_n883), .A3(new_n1193), .ZN(G308));
  NAND3_X1  g768(.A1(new_n949), .A2(new_n883), .A3(new_n1193), .ZN(G225));
endmodule


