//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  INV_X1    g003(.A(G8gat), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n205), .A2(KEYINPUT84), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n204), .B(new_n206), .C1(G1gat), .C2(new_n202), .ZN(new_n207));
  AND2_X1   g006(.A1(new_n205), .A2(KEYINPUT84), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(G57gat), .A2(G64gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G57gat), .A2(G64gat), .ZN(new_n211));
  AND2_X1   g010(.A1(G71gat), .A2(G78gat), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n210), .B(new_n211), .C1(new_n212), .C2(KEYINPUT9), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT86), .B1(G71gat), .B2(G78gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(G71gat), .A2(G78gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(new_n217), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT21), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n209), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(G183gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(G231gat), .A2(G233gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G127gat), .B(G155gat), .ZN(new_n227));
  XOR2_X1   g026(.A(new_n227), .B(KEYINPUT20), .Z(new_n228));
  XNOR2_X1  g027(.A(new_n226), .B(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n221), .A2(new_n222), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(G211gat), .ZN(new_n232));
  XOR2_X1   g031(.A(new_n230), .B(new_n232), .Z(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n229), .A2(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n226), .A2(new_n228), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n226), .A2(new_n228), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(new_n233), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(G43gat), .B(G50gat), .Z(new_n241));
  INV_X1    g040(.A(KEYINPUT15), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n242), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT14), .ZN(new_n245));
  INV_X1    g044(.A(G29gat), .ZN(new_n246));
  INV_X1    g045(.A(G36gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n248), .A2(new_n249), .B1(G29gat), .B2(G36gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n243), .A2(new_n244), .A3(new_n250), .ZN(new_n251));
  OR3_X1    g050(.A1(new_n250), .A2(new_n242), .A3(new_n241), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT17), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G99gat), .A2(G106gat), .ZN(new_n256));
  INV_X1    g055(.A(G85gat), .ZN(new_n257));
  INV_X1    g056(.A(G92gat), .ZN(new_n258));
  AOI22_X1  g057(.A1(KEYINPUT8), .A2(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT7), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(new_n257), .B2(new_n258), .ZN(new_n261));
  NAND3_X1  g060(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  XOR2_X1   g062(.A(G99gat), .B(G106gat), .Z(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(KEYINPUT88), .A3(new_n264), .ZN(new_n265));
  OR2_X1    g064(.A1(new_n263), .A2(new_n264), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT88), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n263), .A2(new_n264), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n251), .A2(KEYINPUT17), .A3(new_n252), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n255), .A2(new_n265), .A3(new_n269), .A4(new_n270), .ZN(new_n271));
  AND3_X1   g070(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n269), .A2(new_n265), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n272), .B1(new_n273), .B2(new_n253), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT89), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n271), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n275), .B1(new_n271), .B2(new_n274), .ZN(new_n278));
  OAI21_X1  g077(.A(G190gat), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n271), .A2(new_n274), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT89), .ZN(new_n281));
  INV_X1    g080(.A(G190gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(new_n276), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n279), .A2(G218gat), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(G218gat), .B1(new_n279), .B2(new_n283), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT90), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n279), .A2(new_n283), .ZN(new_n288));
  INV_X1    g087(.A(G218gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT90), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n291), .A3(new_n284), .ZN(new_n292));
  XNOR2_X1  g091(.A(G134gat), .B(G162gat), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n287), .A2(new_n292), .A3(new_n296), .ZN(new_n297));
  OAI211_X1 g096(.A(KEYINPUT90), .B(new_n295), .C1(new_n285), .C2(new_n286), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n240), .A2(new_n299), .ZN(new_n300));
  AND2_X1   g099(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n282), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT28), .ZN(new_n304));
  NOR2_X1   g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT26), .ZN(new_n307));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n305), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT28), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n311), .B(new_n282), .C1(new_n301), .C2(new_n302), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n304), .A2(new_n309), .A3(new_n310), .A4(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G169gat), .ZN(new_n314));
  INV_X1    g113(.A(G176gat), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n315), .A2(KEYINPUT64), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(KEYINPUT64), .ZN(new_n317));
  OAI211_X1 g116(.A(KEYINPUT23), .B(new_n314), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(G183gat), .A2(G190gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT23), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n306), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT25), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n318), .A2(new_n323), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n313), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G113gat), .B(G120gat), .ZN(new_n329));
  OAI21_X1  g128(.A(G127gat), .B1(new_n329), .B2(KEYINPUT1), .ZN(new_n330));
  INV_X1    g129(.A(G120gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(G113gat), .ZN(new_n332));
  INV_X1    g131(.A(G113gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G120gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT1), .ZN(new_n336));
  INV_X1    g135(.A(G127gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n330), .A2(new_n338), .A3(G134gat), .ZN(new_n339));
  INV_X1    g138(.A(G134gat), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n337), .B1(new_n335), .B2(new_n336), .ZN(new_n341));
  AOI211_X1 g140(.A(KEYINPUT1), .B(G127gat), .C1(new_n332), .C2(new_n334), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT65), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n322), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g144(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n321), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n305), .A2(KEYINPUT23), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n348), .A3(new_n325), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT25), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n328), .A2(new_n339), .A3(new_n343), .A4(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(new_n327), .A3(new_n313), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n343), .A2(new_n339), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G227gat), .A2(G233gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT67), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G15gat), .B(G43gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(G71gat), .ZN(new_n362));
  INV_X1    g161(.A(G99gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n356), .B1(new_n351), .B2(new_n354), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT66), .B(KEYINPUT33), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT32), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  AOI221_X4 g169(.A(new_n368), .B1(new_n366), .B2(new_n364), .C1(new_n355), .C2(new_n357), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n360), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT32), .ZN(new_n374));
  INV_X1    g173(.A(new_n366), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n374), .A2(new_n376), .A3(new_n364), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n367), .A2(new_n369), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(new_n359), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n372), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n358), .A2(KEYINPUT67), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n381), .A2(KEYINPUT34), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n372), .A2(new_n379), .A3(new_n382), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT36), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT36), .B1(new_n384), .B2(new_n385), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT3), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT29), .ZN(new_n392));
  INV_X1    g191(.A(G211gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT69), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT69), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(G211gat), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n396), .A3(G218gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT68), .B(KEYINPUT22), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AND2_X1   g198(.A1(G197gat), .A2(G204gat), .ZN(new_n400));
  NOR2_X1   g199(.A1(G197gat), .A2(G204gat), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G211gat), .B(G218gat), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n392), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n402), .B1(new_n397), .B2(new_n398), .ZN(new_n407));
  INV_X1    g206(.A(new_n405), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n391), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(G148gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(G141gat), .ZN(new_n412));
  INV_X1    g211(.A(G141gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(G148gat), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT2), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT73), .ZN(new_n416));
  INV_X1    g215(.A(G155gat), .ZN(new_n417));
  INV_X1    g216(.A(G162gat), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT73), .B1(G155gat), .B2(G162gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AND2_X1   g220(.A1(G155gat), .A2(G162gat), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n415), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT2), .ZN(new_n424));
  NOR2_X1   g223(.A1(G155gat), .A2(G162gat), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT74), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n427), .A2(G141gat), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n413), .A2(KEYINPUT74), .ZN(new_n429));
  OAI21_X1  g228(.A(G148gat), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n426), .B1(new_n430), .B2(new_n412), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n423), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n412), .A2(new_n414), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n424), .ZN(new_n435));
  INV_X1    g234(.A(new_n422), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n435), .A2(new_n436), .A3(new_n420), .A4(new_n419), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT74), .B(G141gat), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n412), .B1(new_n438), .B2(new_n411), .ZN(new_n439));
  INV_X1    g238(.A(new_n426), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n437), .A2(new_n441), .A3(new_n391), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n392), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT70), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n405), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n407), .B(new_n445), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n410), .A2(new_n433), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(G228gat), .A2(G233gat), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT79), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT29), .B1(new_n432), .B2(new_n391), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n404), .B(new_n445), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n404), .A2(new_n405), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT29), .B1(new_n407), .B2(new_n408), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT3), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI22_X1  g254(.A1(new_n451), .A2(new_n452), .B1(new_n455), .B2(new_n432), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT79), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(new_n448), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n391), .B1(new_n446), .B2(KEYINPUT29), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n459), .A2(new_n433), .B1(new_n446), .B2(new_n443), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n450), .A2(new_n458), .B1(new_n449), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(G22gat), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT81), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n460), .A2(new_n449), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n447), .A2(KEYINPUT79), .A3(new_n449), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n457), .B1(new_n456), .B2(new_n448), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n462), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT80), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT81), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n471), .A3(G22gat), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n461), .A2(KEYINPUT80), .A3(new_n462), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n463), .A2(new_n469), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(G78gat), .B(G106gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(KEYINPUT31), .ZN(new_n476));
  INV_X1    g275(.A(G50gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n476), .B(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n478), .B1(new_n461), .B2(new_n462), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n470), .A2(G22gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n343), .A2(new_n441), .A3(new_n437), .A4(new_n339), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT3), .B1(new_n423), .B2(new_n431), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n353), .A2(new_n487), .A3(new_n442), .ZN(new_n488));
  NAND2_X1  g287(.A1(G225gat), .A2(G233gat), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n432), .A2(KEYINPUT4), .A3(new_n339), .A4(new_n343), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n486), .A2(new_n488), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  XOR2_X1   g290(.A(KEYINPUT76), .B(KEYINPUT5), .Z(new_n492));
  AND2_X1   g291(.A1(new_n492), .A2(KEYINPUT75), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n491), .B(new_n493), .ZN(new_n494));
  XOR2_X1   g293(.A(G1gat), .B(G29gat), .Z(new_n495));
  XNOR2_X1  g294(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G57gat), .B(G85gat), .ZN(new_n498));
  XOR2_X1   g297(.A(new_n497), .B(new_n498), .Z(new_n499));
  NAND2_X1  g298(.A1(new_n433), .A2(new_n353), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n484), .ZN(new_n501));
  INV_X1    g300(.A(new_n489), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n502), .A3(new_n492), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n494), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT40), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n502), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n508), .B(KEYINPUT39), .C1(new_n502), .C2(new_n501), .ZN(new_n509));
  INV_X1    g308(.A(new_n499), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n509), .B(new_n510), .C1(KEYINPUT39), .C2(new_n508), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n505), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n511), .A2(new_n506), .ZN(new_n513));
  INV_X1    g312(.A(G226gat), .ZN(new_n514));
  INV_X1    g313(.A(G233gat), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n352), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT29), .B1(new_n328), .B2(new_n350), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n452), .B(new_n517), .C1(new_n518), .C2(new_n516), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT72), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n352), .A2(new_n392), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(new_n514), .B2(new_n515), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n523), .A2(KEYINPUT72), .A3(new_n452), .A4(new_n517), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT71), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n352), .A2(new_n526), .A3(new_n516), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n526), .B1(new_n352), .B2(new_n516), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n452), .B1(new_n530), .B2(new_n523), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n533));
  XOR2_X1   g332(.A(G8gat), .B(G36gat), .Z(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(G64gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(new_n258), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n532), .A2(new_n533), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n536), .B1(new_n525), .B2(new_n531), .ZN(new_n539));
  INV_X1    g338(.A(new_n529), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n527), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n518), .A2(new_n516), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n446), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n543), .A2(new_n524), .A3(new_n521), .A4(new_n537), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n539), .A2(KEYINPUT30), .A3(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n512), .A2(new_n513), .A3(new_n538), .A4(new_n545), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n494), .A2(KEYINPUT6), .A3(new_n499), .A4(new_n503), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n491), .A2(new_n493), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n491), .A2(new_n493), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n503), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n510), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT6), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(new_n552), .A3(new_n504), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n532), .A2(KEYINPUT37), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n543), .A2(new_n524), .A3(new_n521), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT37), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n537), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT38), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n547), .B(new_n553), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n452), .B1(new_n523), .B2(new_n517), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n561), .B(KEYINPUT82), .Z(new_n562));
  NOR2_X1   g361(.A1(new_n541), .A2(new_n542), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n556), .B1(new_n563), .B2(new_n452), .ZN(new_n564));
  AOI22_X1  g363(.A1(new_n562), .A2(new_n564), .B1(new_n556), .B2(new_n555), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n536), .A2(new_n559), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n544), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n483), .B(new_n546), .C1(new_n560), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n547), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n545), .A2(new_n538), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT78), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n474), .A2(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT78), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n569), .A2(new_n570), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n572), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n390), .A2(new_n568), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT35), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n569), .A2(new_n570), .A3(new_n578), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n372), .A2(new_n379), .A3(new_n382), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n382), .B1(new_n372), .B2(new_n379), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR3_X1   g381(.A1(new_n573), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n569), .A2(new_n570), .A3(new_n574), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n574), .B1(new_n569), .B2(new_n570), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n386), .B(new_n483), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n583), .B1(new_n586), .B2(KEYINPUT35), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT83), .B1(new_n577), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n584), .A2(new_n585), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n483), .A2(new_n386), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT35), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n583), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT83), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n390), .A2(new_n576), .A3(new_n568), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n588), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT11), .B(G169gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(G197gat), .ZN(new_n599));
  XOR2_X1   g398(.A(G113gat), .B(G141gat), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT12), .ZN(new_n602));
  INV_X1    g401(.A(new_n209), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(new_n253), .ZN(new_n604));
  NAND2_X1  g403(.A1(G229gat), .A2(G233gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n209), .A2(new_n255), .A3(new_n270), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT18), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT85), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n602), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n209), .B(new_n253), .Z(new_n612));
  XOR2_X1   g411(.A(new_n605), .B(KEYINPUT13), .Z(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n604), .A2(new_n606), .A3(KEYINPUT18), .A4(new_n605), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(new_n609), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n611), .B(new_n616), .ZN(new_n617));
  AOI22_X1  g416(.A1(new_n218), .A2(new_n219), .B1(new_n266), .B2(new_n268), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n618), .B1(new_n273), .B2(new_n221), .ZN(new_n619));
  OAI21_X1  g418(.A(KEYINPUT91), .B1(new_n619), .B2(KEYINPUT10), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT91), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n220), .B1(new_n265), .B2(new_n269), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n621), .B(new_n622), .C1(new_n623), .C2(new_n618), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n273), .A2(KEYINPUT10), .A3(new_n220), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(G230gat), .A2(G233gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT92), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n619), .A2(new_n629), .ZN(new_n632));
  XNOR2_X1  g431(.A(G120gat), .B(G148gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(new_n315), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n634), .B(G204gat), .Z(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n631), .A2(new_n632), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n626), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n638), .B1(new_n620), .B2(new_n624), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n632), .B1(new_n639), .B2(new_n629), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n635), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  AND4_X1   g442(.A1(new_n300), .A2(new_n597), .A3(new_n617), .A4(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n569), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT93), .B(G1gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(G1324gat));
  XOR2_X1   g447(.A(KEYINPUT16), .B(G8gat), .Z(new_n649));
  INV_X1    g448(.A(KEYINPUT42), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT95), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n649), .B(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n570), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n644), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n652), .B1(new_n655), .B2(new_n650), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n654), .B(KEYINPUT94), .Z(new_n657));
  NOR2_X1   g456(.A1(new_n650), .A2(G8gat), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(G1325gat));
  AOI21_X1  g458(.A(G15gat), .B1(new_n644), .B2(new_n386), .ZN(new_n660));
  INV_X1    g459(.A(new_n390), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n644), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n660), .B1(G15gat), .B2(new_n662), .ZN(G1326gat));
  NAND2_X1  g462(.A1(new_n644), .A2(new_n573), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT96), .B(KEYINPUT43), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G22gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n664), .B(new_n666), .ZN(G1327gat));
  NAND2_X1  g466(.A1(new_n297), .A2(new_n298), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n668), .B1(new_n588), .B2(new_n596), .ZN(new_n669));
  INV_X1    g468(.A(new_n617), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n239), .A2(new_n670), .A3(new_n642), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n672), .A2(new_n246), .A3(new_n645), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT45), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n675), .B(new_n299), .C1(new_n577), .C2(new_n587), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(new_n669), .B2(new_n675), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n671), .B(KEYINPUT97), .Z(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(G29gat), .B1(new_n679), .B2(new_n569), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n674), .A2(new_n680), .ZN(G1328gat));
  NAND4_X1  g480(.A1(new_n669), .A2(new_n247), .A3(new_n653), .A4(new_n671), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT98), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(KEYINPUT46), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT99), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT46), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n684), .A2(new_n690), .A3(new_n685), .ZN(new_n691));
  OAI21_X1  g490(.A(G36gat), .B1(new_n679), .B2(new_n570), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n686), .A2(KEYINPUT99), .A3(KEYINPUT46), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n689), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT100), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n689), .A2(new_n693), .A3(KEYINPUT100), .A4(new_n694), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(G1329gat));
  INV_X1    g498(.A(KEYINPUT47), .ZN(new_n700));
  INV_X1    g499(.A(G43gat), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n672), .A2(new_n701), .A3(new_n386), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(KEYINPUT101), .Z(new_n703));
  INV_X1    g502(.A(new_n679), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n701), .B1(new_n704), .B2(new_n661), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n700), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n700), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n707), .A2(KEYINPUT102), .A3(new_n702), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT102), .B1(new_n707), .B2(new_n702), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n706), .B1(new_n708), .B2(new_n709), .ZN(G1330gat));
  AOI21_X1  g509(.A(G50gat), .B1(new_n672), .B2(new_n573), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n679), .A2(new_n477), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n711), .B1(new_n712), .B2(new_n573), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n713), .B(KEYINPUT48), .Z(G1331gat));
  AOI21_X1  g513(.A(new_n643), .B1(new_n593), .B2(new_n595), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(new_n300), .A3(new_n670), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n569), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(G57gat), .Z(G1332gat));
  AOI211_X1 g517(.A(new_n570), .B(new_n716), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n719));
  NOR2_X1   g518(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1333gat));
  OAI21_X1  g520(.A(G71gat), .B1(new_n716), .B2(new_n390), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n386), .B(KEYINPUT103), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n723), .A2(G71gat), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n716), .B2(new_n724), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g525(.A1(new_n716), .A2(new_n483), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT104), .B(G78gat), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1335gat));
  NOR2_X1   g528(.A1(new_n239), .A2(new_n617), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n299), .B(new_n730), .C1(new_n577), .C2(new_n587), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n731), .A2(KEYINPUT51), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(KEYINPUT51), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n732), .A2(new_n642), .A3(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(G85gat), .B1(new_n735), .B2(new_n645), .ZN(new_n736));
  INV_X1    g535(.A(new_n676), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n577), .A2(new_n587), .A3(KEYINPUT83), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n594), .B1(new_n593), .B2(new_n595), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n299), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n737), .B1(new_n740), .B2(KEYINPUT44), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n730), .A2(new_n642), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT105), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n744));
  INV_X1    g543(.A(new_n742), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n677), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n257), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n736), .B1(new_n747), .B2(new_n645), .ZN(G1336gat));
  AOI21_X1  g547(.A(new_n570), .B1(new_n743), .B2(new_n746), .ZN(new_n749));
  OAI21_X1  g548(.A(KEYINPUT106), .B1(new_n749), .B2(new_n258), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n258), .A3(new_n653), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n677), .A2(new_n744), .A3(new_n745), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n744), .B1(new_n677), .B2(new_n745), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n653), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT106), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(new_n755), .A3(G92gat), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n750), .A2(new_n751), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT52), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n677), .A2(new_n745), .ZN(new_n759));
  OAI21_X1  g558(.A(G92gat), .B1(new_n759), .B2(new_n570), .ZN(new_n760));
  XOR2_X1   g559(.A(KEYINPUT107), .B(KEYINPUT52), .Z(new_n761));
  NAND3_X1  g560(.A1(new_n760), .A2(new_n751), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n758), .A2(new_n762), .ZN(G1337gat));
  NAND3_X1  g562(.A1(new_n735), .A2(new_n363), .A3(new_n386), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n390), .B1(new_n743), .B2(new_n746), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n765), .B2(new_n363), .ZN(G1338gat));
  OAI21_X1  g565(.A(G106gat), .B1(new_n759), .B2(new_n483), .ZN(new_n767));
  OR3_X1    g566(.A1(new_n734), .A2(G106gat), .A3(new_n483), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n573), .B1(new_n752), .B2(new_n753), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G106gat), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n772), .A2(new_n768), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n770), .B1(new_n773), .B2(new_n769), .ZN(G1339gat));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n639), .B2(new_n629), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n631), .A2(new_n778), .ZN(new_n779));
  XOR2_X1   g578(.A(KEYINPUT108), .B(KEYINPUT54), .Z(new_n780));
  NAND3_X1  g579(.A1(new_n627), .A2(new_n630), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n635), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n776), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n631), .A2(new_n778), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n784), .A2(KEYINPUT55), .A3(new_n635), .A4(new_n781), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n783), .A2(new_n617), .A3(new_n637), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n605), .B1(new_n604), .B2(new_n606), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n787), .A2(KEYINPUT109), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(KEYINPUT109), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n788), .B(new_n789), .C1(new_n612), .C2(new_n613), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n601), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT110), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n614), .A2(new_n609), .A3(new_n602), .A4(new_n615), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n790), .A2(new_n794), .A3(new_n601), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n792), .A2(new_n642), .A3(new_n793), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n786), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n786), .A2(KEYINPUT111), .A3(new_n796), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(new_n668), .A3(new_n800), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n792), .A2(new_n793), .A3(new_n795), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n783), .A2(new_n637), .A3(new_n785), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n299), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n239), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  NOR4_X1   g604(.A1(new_n240), .A2(new_n299), .A3(new_n617), .A4(new_n642), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT112), .B1(new_n807), .B2(new_n573), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n809), .B(new_n483), .C1(new_n805), .C2(new_n806), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n653), .A2(new_n569), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n812), .A2(new_n582), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n617), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n775), .B1(new_n816), .B2(G113gat), .ZN(new_n817));
  AOI211_X1 g616(.A(KEYINPUT113), .B(new_n333), .C1(new_n815), .C2(new_n617), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n807), .A2(new_n573), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n386), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(new_n814), .ZN(new_n821));
  XOR2_X1   g620(.A(new_n821), .B(KEYINPUT114), .Z(new_n822));
  NAND2_X1  g621(.A1(new_n617), .A2(new_n333), .ZN(new_n823));
  OAI22_X1  g622(.A1(new_n817), .A2(new_n818), .B1(new_n822), .B2(new_n823), .ZN(G1340gat));
  INV_X1    g623(.A(new_n815), .ZN(new_n825));
  OAI21_X1  g624(.A(G120gat), .B1(new_n825), .B2(new_n643), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n642), .A2(new_n331), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n826), .B1(new_n822), .B2(new_n827), .ZN(G1341gat));
  AOI21_X1  g627(.A(G127gat), .B1(new_n821), .B2(new_n239), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n825), .A2(new_n240), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(G127gat), .ZN(G1342gat));
  NAND3_X1  g630(.A1(new_n821), .A2(new_n340), .A3(new_n299), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n832), .B(KEYINPUT56), .Z(new_n833));
  OAI21_X1  g632(.A(G134gat), .B1(new_n825), .B2(new_n668), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(G1343gat));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(KEYINPUT58), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n836), .A2(KEYINPUT58), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n661), .A2(new_n814), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT115), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n797), .A2(new_n668), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n239), .B1(new_n804), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n573), .B1(new_n842), .B2(new_n806), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n845), .B(new_n846), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n786), .A2(KEYINPUT111), .A3(new_n796), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT111), .B1(new_n786), .B2(new_n796), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n848), .A2(new_n849), .A3(new_n299), .ZN(new_n850));
  INV_X1    g649(.A(new_n804), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n240), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n806), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n483), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(KEYINPUT57), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n617), .B(new_n840), .C1(new_n847), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n438), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n854), .A2(new_n839), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n413), .A3(new_n617), .ZN(new_n860));
  AOI211_X1 g659(.A(new_n837), .B(new_n838), .C1(new_n857), .C2(new_n860), .ZN(new_n861));
  AND4_X1   g660(.A1(new_n836), .A2(new_n857), .A3(KEYINPUT58), .A4(new_n860), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(G1344gat));
  OR2_X1    g662(.A1(new_n847), .A2(new_n855), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n864), .A2(new_n840), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n866), .A3(new_n642), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT118), .B1(new_n843), .B2(new_n844), .ZN(new_n868));
  OAI211_X1 g667(.A(KEYINPUT57), .B(new_n573), .C1(new_n805), .C2(new_n806), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n642), .A3(new_n840), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n866), .B1(new_n859), .B2(new_n642), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n867), .B(new_n875), .C1(G148gat), .C2(new_n876), .ZN(G1345gat));
  AOI21_X1  g676(.A(G155gat), .B1(new_n859), .B2(new_n239), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n239), .A2(G155gat), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT119), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n878), .B1(new_n865), .B2(new_n880), .ZN(G1346gat));
  NAND3_X1  g680(.A1(new_n865), .A2(G162gat), .A3(new_n299), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n418), .B1(new_n858), .B2(new_n668), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(G1347gat));
  NOR2_X1   g683(.A1(new_n645), .A2(new_n570), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n820), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n314), .A3(new_n617), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n723), .A2(new_n886), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n812), .A2(new_n670), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n888), .B1(new_n891), .B2(new_n314), .ZN(G1348gat));
  AOI21_X1  g691(.A(G176gat), .B1(new_n887), .B2(new_n642), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n812), .A2(new_n890), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n643), .A2(new_n316), .A3(new_n317), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(G1349gat));
  NAND2_X1  g695(.A1(new_n852), .A2(new_n853), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n809), .B1(new_n897), .B2(new_n483), .ZN(new_n898));
  INV_X1    g697(.A(new_n810), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n239), .B(new_n889), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n811), .A2(KEYINPUT120), .A3(new_n239), .A4(new_n889), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(G183gat), .A3(new_n903), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n887), .B(new_n239), .C1(new_n302), .C2(new_n301), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(KEYINPUT122), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT121), .ZN(new_n907));
  NAND2_X1  g706(.A1(KEYINPUT121), .A2(KEYINPUT60), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n904), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT60), .ZN(new_n910));
  AOI22_X1  g709(.A1(new_n907), .A2(new_n909), .B1(new_n910), .B2(new_n906), .ZN(G1350gat));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n299), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(G190gat), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n913), .A2(KEYINPUT123), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n887), .A2(new_n282), .A3(new_n299), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(KEYINPUT123), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n914), .A2(KEYINPUT123), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n912), .A2(G190gat), .A3(new_n917), .A4(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n915), .A2(new_n916), .A3(new_n919), .ZN(G1351gat));
  OAI21_X1  g719(.A(KEYINPUT124), .B1(new_n870), .B2(new_n872), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n661), .A2(new_n886), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n868), .A2(new_n869), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n923), .B(new_n924), .C1(new_n871), .C2(new_n869), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n921), .A2(new_n922), .A3(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(G197gat), .B1(new_n926), .B2(new_n670), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n854), .A2(new_n922), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n928), .A2(G197gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n927), .B1(new_n670), .B2(new_n929), .ZN(G1352gat));
  NAND4_X1  g729(.A1(new_n921), .A2(new_n642), .A3(new_n922), .A4(new_n925), .ZN(new_n931));
  XNOR2_X1  g730(.A(KEYINPUT125), .B(G204gat), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n928), .A2(new_n643), .A3(new_n932), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT62), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT126), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT126), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n933), .A2(new_n938), .A3(new_n935), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(G1353gat));
  NAND3_X1  g739(.A1(new_n873), .A2(new_n239), .A3(new_n922), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G211gat), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT63), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n942), .B(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n928), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n394), .A2(new_n396), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n945), .A2(new_n239), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n944), .A2(new_n947), .ZN(G1354gat));
  NAND4_X1  g747(.A1(new_n921), .A2(new_n299), .A3(new_n922), .A4(new_n925), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G218gat), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n945), .A2(new_n289), .A3(new_n299), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n950), .A2(KEYINPUT127), .A3(new_n951), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1355gat));
endmodule


