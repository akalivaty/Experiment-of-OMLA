//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983, new_n984;
  INV_X1    g000(.A(G36gat), .ZN(new_n202));
  AND2_X1   g001(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n206), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209));
  AND2_X1   g008(.A1(G43gat), .A2(G50gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(G43gat), .A2(G50gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NOR3_X1   g011(.A1(new_n208), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT88), .ZN(new_n215));
  INV_X1    g014(.A(G43gat), .ZN(new_n216));
  INV_X1    g015(.A(G50gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G43gat), .A2(G50gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(KEYINPUT87), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n209), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n218), .A2(KEYINPUT87), .A3(KEYINPUT15), .A4(new_n219), .ZN(new_n222));
  AOI221_X4 g021(.A(new_n215), .B1(new_n205), .B2(new_n207), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n222), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT88), .B1(new_n224), .B2(new_n208), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n214), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g025(.A1(G15gat), .A2(G22gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(G15gat), .A2(G22gat), .ZN(new_n228));
  INV_X1    g027(.A(G1gat), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n227), .A2(new_n228), .B1(KEYINPUT16), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT89), .ZN(new_n232));
  INV_X1    g031(.A(G8gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n227), .A2(new_n229), .A3(new_n228), .ZN(new_n235));
  NAND2_X1  g034(.A1(KEYINPUT89), .A2(G8gat), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n231), .A2(new_n234), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n235), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n232), .B(new_n233), .C1(new_n238), .C2(new_n230), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(KEYINPUT90), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT90), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n237), .A2(new_n239), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n226), .A2(KEYINPUT17), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT15), .B1(new_n212), .B2(KEYINPUT87), .ZN(new_n248));
  INV_X1    g047(.A(new_n222), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n208), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n215), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n224), .A2(KEYINPUT88), .A3(new_n208), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT17), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n254), .A3(new_n214), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n246), .B1(new_n247), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT91), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n242), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n246), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n254), .B1(new_n253), .B2(new_n214), .ZN(new_n260));
  AOI211_X1 g059(.A(KEYINPUT17), .B(new_n213), .C1(new_n251), .C2(new_n252), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n257), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G229gat), .A2(G233gat), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n264), .A2(KEYINPUT92), .A3(KEYINPUT18), .A4(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n242), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n267), .B1(new_n268), .B2(KEYINPUT91), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n269), .A2(KEYINPUT18), .A3(new_n265), .A4(new_n262), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT92), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G113gat), .B(G141gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(G197gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT11), .B(G169gat), .ZN(new_n276));
  XOR2_X1   g075(.A(new_n275), .B(new_n276), .Z(new_n277));
  XOR2_X1   g076(.A(new_n277), .B(KEYINPUT12), .Z(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(new_n265), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n213), .B1(new_n251), .B2(new_n252), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(new_n240), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n282), .B1(new_n242), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n265), .A3(new_n262), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT18), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AND3_X1   g087(.A1(new_n273), .A2(new_n279), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n279), .B1(new_n273), .B2(new_n288), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT36), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n293), .A2(KEYINPUT65), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(KEYINPUT65), .ZN(new_n295));
  NAND3_X1  g094(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n296), .B1(G183gat), .B2(G190gat), .ZN(new_n297));
  NOR3_X1   g096(.A1(new_n294), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT23), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT23), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n301), .B1(G169gat), .B2(G176gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n300), .B1(new_n302), .B2(new_n299), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT25), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n297), .A2(new_n293), .ZN(new_n305));
  NOR3_X1   g104(.A1(new_n305), .A2(new_n303), .A3(KEYINPUT25), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT27), .B(G183gat), .ZN(new_n308));
  INV_X1    g107(.A(G190gat), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT28), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT66), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n308), .B(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n309), .A2(KEYINPUT28), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n310), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n315), .B(KEYINPUT67), .ZN(new_n316));
  NOR3_X1   g115(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n317), .B1(G169gat), .B2(G176gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G183gat), .A2(G190gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n304), .B(new_n307), .C1(new_n314), .C2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G127gat), .B(G134gat), .ZN(new_n323));
  XOR2_X1   g122(.A(G113gat), .B(G120gat), .Z(new_n324));
  INV_X1    g123(.A(KEYINPUT1), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n327));
  AND2_X1   g126(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n323), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT68), .B(G120gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(G113gat), .ZN(new_n332));
  INV_X1    g131(.A(G113gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G120gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n330), .A2(new_n335), .A3(KEYINPUT70), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT70), .ZN(new_n337));
  INV_X1    g136(.A(new_n334), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n338), .B1(new_n331), .B2(G113gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n337), .B1(new_n339), .B2(new_n329), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n326), .B1(new_n336), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n322), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n336), .A2(new_n340), .ZN(new_n343));
  INV_X1    g142(.A(new_n326), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(KEYINPUT27), .B(G183gat), .Z(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(new_n311), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n308), .A2(KEYINPUT66), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n348), .A3(new_n313), .ZN(new_n349));
  INV_X1    g148(.A(new_n310), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n316), .A2(new_n318), .B1(G183gat), .B2(G190gat), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n306), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n345), .A2(new_n353), .A3(new_n304), .ZN(new_n354));
  NAND2_X1  g153(.A1(G227gat), .A2(G233gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(KEYINPUT64), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n342), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT32), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT33), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  XOR2_X1   g159(.A(G15gat), .B(G43gat), .Z(new_n361));
  XNOR2_X1  g160(.A(G71gat), .B(G99gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n358), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  OR2_X1    g163(.A1(new_n356), .A2(KEYINPUT34), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n365), .B1(new_n342), .B2(new_n354), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n345), .B1(new_n304), .B2(new_n353), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n322), .A2(new_n341), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n355), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n366), .B1(new_n369), .B2(KEYINPUT34), .ZN(new_n370));
  INV_X1    g169(.A(new_n363), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n357), .B(KEYINPUT32), .C1(new_n359), .C2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n364), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n370), .B1(new_n364), .B2(new_n372), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n292), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n364), .A2(new_n372), .ZN(new_n377));
  INV_X1    g176(.A(new_n370), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n379), .A2(KEYINPUT36), .A3(new_n373), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT30), .ZN(new_n382));
  INV_X1    g181(.A(G211gat), .ZN(new_n383));
  INV_X1    g182(.A(G218gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT72), .ZN(new_n386));
  NAND2_X1  g185(.A1(G211gat), .A2(G218gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT71), .ZN(new_n391));
  AND2_X1   g190(.A1(G197gat), .A2(G204gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(G197gat), .A2(G204gat), .ZN(new_n393));
  OAI22_X1  g192(.A1(new_n390), .A2(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n390), .A2(new_n391), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n389), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n392), .A2(new_n393), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT22), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n387), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT71), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n398), .A2(new_n388), .A3(new_n401), .A4(new_n395), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G226gat), .A2(G233gat), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT29), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n406), .B1(new_n322), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n405), .B1(new_n353), .B2(new_n304), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n404), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n322), .A2(new_n406), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT29), .B1(new_n353), .B2(new_n304), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n411), .B(new_n403), .C1(new_n412), .C2(new_n406), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G8gat), .B(G36gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(KEYINPUT73), .ZN(new_n416));
  XNOR2_X1  g215(.A(G64gat), .B(G92gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n382), .B1(new_n414), .B2(new_n419), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n410), .A2(KEYINPUT30), .A3(new_n413), .A4(new_n418), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n418), .B(KEYINPUT74), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n414), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT2), .ZN(new_n425));
  INV_X1    g224(.A(G148gat), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n426), .A2(G141gat), .ZN(new_n427));
  INV_X1    g226(.A(G141gat), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(G148gat), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n425), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT75), .ZN(new_n431));
  NAND2_X1  g230(.A1(G155gat), .A2(G162gat), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(G155gat), .A2(G162gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n430), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n428), .A2(G148gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n426), .A2(G141gat), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT2), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n434), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n432), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT75), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  OR3_X1    g241(.A1(new_n426), .A2(KEYINPUT76), .A3(G141gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n437), .A2(KEYINPUT76), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT77), .B(G148gat), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n443), .B(new_n444), .C1(new_n445), .C2(new_n428), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n432), .B1(new_n440), .B2(KEYINPUT2), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n436), .A2(new_n442), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n343), .A2(new_n448), .A3(new_n344), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT4), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT4), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n341), .A2(new_n451), .A3(new_n448), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(G225gat), .A2(G233gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n446), .A2(new_n447), .ZN(new_n455));
  NOR3_X1   g254(.A1(new_n439), .A2(new_n441), .A3(KEYINPUT75), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n431), .B1(new_n430), .B2(new_n435), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT78), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT3), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT3), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT78), .B1(new_n448), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n448), .A2(new_n461), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n460), .A2(new_n462), .A3(new_n345), .A4(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n453), .A2(new_n454), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n454), .ZN(new_n466));
  INV_X1    g265(.A(new_n449), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n341), .A2(new_n448), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT5), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n453), .A2(KEYINPUT5), .A3(new_n454), .A4(new_n464), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G1gat), .B(G29gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT0), .ZN(new_n475));
  XNOR2_X1  g274(.A(G57gat), .B(G85gat), .ZN(new_n476));
  XOR2_X1   g275(.A(new_n475), .B(new_n476), .Z(new_n477));
  NAND2_X1  g276(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n479));
  INV_X1    g278(.A(new_n477), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n471), .A2(new_n480), .A3(new_n472), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n471), .A2(KEYINPUT6), .A3(new_n480), .A4(new_n472), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n424), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n407), .B1(new_n458), .B2(KEYINPUT3), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n404), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT29), .B1(new_n397), .B2(new_n402), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n458), .B1(new_n487), .B2(KEYINPUT3), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT81), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n458), .B(KEYINPUT81), .C1(new_n487), .C2(KEYINPUT3), .ZN(new_n491));
  NAND2_X1  g290(.A1(G228gat), .A2(G233gat), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n486), .A2(new_n490), .A3(new_n491), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT82), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n492), .B1(new_n485), .B2(new_n404), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT82), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n496), .A2(new_n497), .A3(new_n491), .A4(new_n490), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n492), .B(KEYINPUT80), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n398), .A2(new_n395), .A3(new_n401), .ZN(new_n502));
  XNOR2_X1  g301(.A(G211gat), .B(G218gat), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT29), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(new_n503), .B2(new_n502), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n461), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n458), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n501), .B1(new_n507), .B2(new_n486), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n499), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G78gat), .B(G106gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(new_n217), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n512), .B(new_n513), .Z(new_n514));
  NAND2_X1  g313(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT83), .B(G22gat), .ZN(new_n516));
  INV_X1    g315(.A(new_n514), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n499), .A2(new_n509), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n516), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n517), .B1(new_n499), .B2(new_n509), .ZN(new_n521));
  AOI211_X1 g320(.A(new_n508), .B(new_n514), .C1(new_n495), .C2(new_n498), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n381), .B(KEYINPUT84), .C1(new_n484), .C2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n381), .B1(new_n484), .B2(new_n524), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT84), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT86), .ZN(new_n529));
  NOR2_X1   g328(.A1(KEYINPUT85), .A2(KEYINPUT40), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n454), .B1(new_n453), .B2(new_n464), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT39), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n345), .A2(new_n458), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(new_n454), .A3(new_n449), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT39), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n477), .B1(new_n531), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n530), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n536), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n453), .A2(new_n464), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n539), .B1(new_n540), .B2(new_n454), .ZN(new_n541));
  INV_X1    g340(.A(new_n530), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n531), .A2(new_n532), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n541), .A2(new_n477), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n538), .A2(new_n544), .A3(new_n481), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n545), .A2(new_n424), .B1(new_n519), .B2(new_n523), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n414), .A2(new_n419), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT37), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n410), .A2(new_n548), .A3(new_n413), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT38), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n422), .A2(new_n550), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n548), .B1(new_n410), .B2(new_n413), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n547), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n549), .A2(new_n419), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT38), .B1(new_n556), .B2(new_n553), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n482), .A2(new_n555), .A3(new_n483), .A4(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n529), .B1(new_n546), .B2(new_n558), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n424), .A2(new_n538), .A3(new_n544), .A4(new_n481), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n558), .A2(new_n529), .A3(new_n524), .A4(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n525), .B(new_n528), .C1(new_n559), .C2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT35), .ZN(new_n564));
  INV_X1    g363(.A(new_n484), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n374), .A2(new_n375), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n524), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n564), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n484), .A2(KEYINPUT35), .A3(new_n524), .A4(new_n566), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n291), .B1(new_n563), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G57gat), .B(G64gat), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G71gat), .B(G78gat), .Z(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT21), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(G127gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n576), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n241), .B1(new_n583), .B2(KEYINPUT21), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n582), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n586));
  INV_X1    g385(.A(G155gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G183gat), .B(G211gat), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n588), .B(new_n589), .Z(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n585), .A2(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n582), .A2(new_n584), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n582), .A2(new_n584), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n594), .A3(new_n590), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G232gat), .A2(G233gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT94), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT41), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G134gat), .B(G162gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(G85gat), .A2(G92gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT7), .ZN(new_n606));
  INV_X1    g405(.A(G99gat), .ZN(new_n607));
  INV_X1    g406(.A(G106gat), .ZN(new_n608));
  OAI21_X1  g407(.A(KEYINPUT8), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(KEYINPUT95), .B(G85gat), .Z(new_n610));
  OAI211_X1 g409(.A(new_n606), .B(new_n609), .C1(G92gat), .C2(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G99gat), .B(G106gat), .Z(new_n612));
  AND2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n615), .B1(new_n247), .B2(new_n255), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n598), .A2(new_n599), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n617), .B1(new_n226), .B2(new_n615), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n604), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n615), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n621), .B1(new_n260), .B2(new_n261), .ZN(new_n622));
  INV_X1    g421(.A(new_n604), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n622), .A2(new_n623), .A3(new_n618), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n603), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n622), .A2(new_n618), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT96), .B1(new_n627), .B2(new_n604), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n603), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n627), .A2(KEYINPUT96), .A3(new_n604), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT97), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n619), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n602), .B1(new_n633), .B2(new_n623), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT96), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n631), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT97), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n626), .B1(new_n632), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n641), .B(KEYINPUT98), .Z(new_n642));
  NAND2_X1  g441(.A1(new_n615), .A2(new_n583), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n576), .B1(new_n613), .B2(new_n614), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n615), .A2(KEYINPUT10), .A3(new_n583), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n642), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n643), .A2(new_n645), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n648), .B1(new_n649), .B2(new_n642), .ZN(new_n650));
  XNOR2_X1  g449(.A(G120gat), .B(G148gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(G176gat), .B(G204gat), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n651), .B(new_n652), .Z(new_n653));
  OR2_X1    g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n646), .A2(new_n647), .ZN(new_n655));
  INV_X1    g454(.A(new_n642), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n649), .A2(new_n642), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(new_n658), .A3(new_n653), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n596), .A2(new_n640), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n571), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n482), .ZN(new_n663));
  INV_X1    g462(.A(new_n483), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT99), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(new_n229), .ZN(G1324gat));
  INV_X1    g467(.A(new_n662), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT16), .B(G8gat), .Z(new_n670));
  NAND4_X1  g469(.A1(new_n669), .A2(KEYINPUT42), .A3(new_n424), .A4(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n424), .ZN(new_n672));
  OR3_X1    g471(.A1(new_n662), .A2(KEYINPUT101), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT101), .B1(new_n662), .B2(new_n672), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(G8gat), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n670), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n676), .B1(new_n673), .B2(new_n674), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT100), .B(KEYINPUT42), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n671), .B(new_n675), .C1(new_n677), .C2(new_n678), .ZN(G1325gat));
  INV_X1    g478(.A(G15gat), .ZN(new_n680));
  INV_X1    g479(.A(new_n566), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n680), .B1(new_n662), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(KEYINPUT102), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(KEYINPUT102), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n381), .A2(new_n680), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT103), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n683), .A2(new_n684), .B1(new_n669), .B2(new_n686), .ZN(G1326gat));
  OR3_X1    g486(.A1(new_n662), .A2(KEYINPUT104), .A3(new_n524), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT104), .B1(new_n662), .B2(new_n524), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT43), .B(G22gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  INV_X1    g491(.A(new_n660), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n596), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n630), .A2(KEYINPUT97), .A3(new_n631), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n637), .A2(new_n638), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n625), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n571), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n666), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(new_n206), .A3(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT45), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n563), .A2(new_n570), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n697), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n558), .A2(new_n524), .A3(new_n560), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT86), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n526), .B1(new_n709), .B2(new_n561), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n568), .A2(new_n569), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n640), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n705), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n707), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n694), .A2(new_n291), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n714), .A2(new_n700), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G29gat), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n717), .A3(new_n718), .ZN(G1328gat));
  NOR2_X1   g518(.A1(new_n672), .A2(G36gat), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n699), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT46), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n707), .A2(new_n713), .A3(new_n424), .A4(new_n715), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G36gat), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n699), .A2(new_n725), .A3(new_n720), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n722), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT105), .ZN(G1329gat));
  INV_X1    g527(.A(new_n381), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n707), .A2(new_n713), .A3(new_n729), .A4(new_n715), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G43gat), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT47), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n699), .A2(new_n216), .A3(new_n566), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n733), .B(new_n735), .ZN(G1330gat));
  INV_X1    g535(.A(new_n524), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n707), .A2(new_n713), .A3(new_n737), .A4(new_n715), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n217), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(new_n739), .B2(new_n738), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n699), .A2(new_n217), .A3(new_n737), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT48), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n738), .A2(G50gat), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n743), .B1(new_n746), .B2(new_n742), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1331gat));
  NAND2_X1  g547(.A1(new_n592), .A2(new_n595), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n291), .A2(new_n749), .A3(new_n697), .A4(new_n660), .ZN(new_n750));
  INV_X1    g549(.A(new_n526), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(new_n559), .B2(new_n562), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n750), .B1(new_n752), .B2(new_n570), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n700), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n424), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n757));
  XOR2_X1   g556(.A(KEYINPUT49), .B(G64gat), .Z(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n756), .B2(new_n758), .ZN(G1333gat));
  NAND2_X1  g558(.A1(new_n753), .A2(new_n566), .ZN(new_n760));
  AOI21_X1  g559(.A(G71gat), .B1(new_n760), .B2(KEYINPUT108), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(KEYINPUT108), .B2(new_n760), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n753), .A2(G71gat), .A3(new_n729), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g564(.A1(new_n753), .A2(new_n737), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g566(.A1(new_n273), .A2(new_n288), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n278), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n273), .A2(new_n279), .A3(new_n288), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n596), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT109), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n773), .A2(new_n693), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n714), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n700), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n610), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n712), .B2(new_n773), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n752), .A2(new_n570), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n771), .B(KEYINPUT109), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n780), .A2(KEYINPUT51), .A3(new_n640), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n780), .A2(new_n640), .A3(new_n781), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n784), .B1(new_n786), .B2(new_n778), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  OR3_X1    g589(.A1(new_n666), .A2(new_n610), .A3(new_n693), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n777), .B1(new_n790), .B2(new_n791), .ZN(G1336gat));
  NAND4_X1  g591(.A1(new_n707), .A2(new_n713), .A3(new_n424), .A4(new_n774), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n793), .A2(KEYINPUT111), .A3(G92gat), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT111), .B1(new_n793), .B2(G92gat), .ZN(new_n795));
  OR3_X1    g594(.A1(new_n693), .A2(new_n672), .A3(G92gat), .ZN(new_n796));
  XOR2_X1   g595(.A(new_n796), .B(KEYINPUT112), .Z(new_n797));
  AOI21_X1  g596(.A(new_n797), .B1(new_n779), .B2(new_n782), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n794), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n801));
  INV_X1    g600(.A(new_n797), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n801), .B1(new_n789), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT110), .B1(new_n779), .B2(new_n782), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n801), .B(new_n802), .C1(new_n804), .C2(new_n787), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(new_n793), .B2(G92gat), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI22_X1  g606(.A1(new_n799), .A2(new_n800), .B1(new_n803), .B2(new_n807), .ZN(G1337gat));
  AND2_X1   g607(.A1(new_n775), .A2(new_n729), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n566), .A2(new_n660), .A3(new_n607), .ZN(new_n810));
  OAI22_X1  g609(.A1(new_n809), .A2(new_n607), .B1(new_n790), .B2(new_n810), .ZN(G1338gat));
  NOR3_X1   g610(.A1(new_n524), .A2(new_n693), .A3(G106gat), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n789), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n714), .A2(new_n737), .A3(new_n774), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G106gat), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI22_X1  g616(.A1(new_n814), .A2(G106gat), .B1(new_n783), .B2(new_n812), .ZN(new_n818));
  OAI22_X1  g617(.A1(new_n813), .A2(new_n817), .B1(new_n818), .B2(new_n816), .ZN(G1339gat));
  NAND3_X1  g618(.A1(new_n242), .A2(new_n284), .A3(new_n282), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT114), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n242), .A2(new_n284), .A3(new_n822), .A4(new_n282), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n268), .A2(KEYINPUT91), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n262), .A3(new_n242), .ZN(new_n826));
  INV_X1    g625(.A(new_n265), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n824), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n277), .ZN(new_n829));
  OAI21_X1  g628(.A(KEYINPUT115), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n265), .B1(new_n269), .B2(new_n262), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n831), .B(new_n277), .C1(new_n832), .C2(new_n824), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n770), .A2(new_n834), .A3(new_n660), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n770), .A2(new_n834), .A3(KEYINPUT117), .A4(new_n660), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n646), .A2(new_n647), .A3(new_n642), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n657), .A2(KEYINPUT54), .A3(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n653), .B1(new_n648), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n840), .A2(KEYINPUT55), .A3(new_n842), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n845), .A2(new_n659), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(new_n289), .B2(new_n290), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n837), .A2(new_n838), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n697), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n640), .A2(new_n770), .A3(new_n847), .A4(new_n834), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT116), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n770), .A2(new_n834), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n845), .A2(new_n659), .A3(new_n846), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n695), .A2(new_n696), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n854), .B1(new_n855), .B2(new_n626), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n853), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n852), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n749), .B1(new_n850), .B2(new_n859), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n661), .A2(new_n291), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n862), .A2(new_n567), .A3(new_n666), .ZN(new_n863));
  INV_X1    g662(.A(new_n291), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n864), .A3(new_n672), .ZN(new_n865));
  AND2_X1   g664(.A1(KEYINPUT118), .A2(G113gat), .ZN(new_n866));
  NOR2_X1   g665(.A1(KEYINPUT118), .A2(G113gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n868), .B1(new_n865), .B2(new_n866), .ZN(G1340gat));
  NAND2_X1  g668(.A1(new_n863), .A2(new_n672), .ZN(new_n870));
  OAI21_X1  g669(.A(G120gat), .B1(new_n870), .B2(new_n693), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n660), .A2(new_n331), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT119), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n871), .B1(new_n870), .B2(new_n873), .ZN(G1341gat));
  NAND3_X1  g673(.A1(new_n863), .A2(new_n672), .A3(new_n749), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(G127gat), .ZN(G1342gat));
  NOR3_X1   g675(.A1(new_n697), .A2(G134gat), .A3(new_n424), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n863), .A2(new_n877), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n878), .A2(KEYINPUT56), .ZN(new_n879));
  OAI21_X1  g678(.A(G134gat), .B1(new_n870), .B2(new_n697), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(KEYINPUT56), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(G1343gat));
  AOI21_X1  g681(.A(new_n854), .B1(new_n769), .B2(new_n770), .ZN(new_n883));
  INV_X1    g682(.A(new_n835), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n697), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n859), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n861), .B1(new_n886), .B2(new_n596), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT57), .B1(new_n887), .B2(new_n524), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n889), .B(new_n737), .C1(new_n860), .C2(new_n861), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n666), .A2(new_n424), .A3(new_n729), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n888), .A2(new_n890), .A3(new_n864), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(G141gat), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n862), .A2(new_n666), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n729), .A2(new_n524), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n864), .A2(new_n428), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT120), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n894), .A2(new_n672), .A3(new_n895), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT58), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT58), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n893), .A2(new_n901), .A3(new_n898), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(G1344gat));
  OR2_X1    g702(.A1(new_n860), .A2(new_n861), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n904), .A2(new_n672), .A3(new_n700), .A4(new_n895), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT59), .B1(new_n905), .B2(new_n693), .ZN(new_n906));
  INV_X1    g705(.A(new_n445), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n737), .B1(new_n860), .B2(new_n861), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n661), .A2(KEYINPUT121), .A3(new_n291), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT121), .B1(new_n661), .B2(new_n291), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n856), .A2(KEYINPUT122), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n914), .B1(new_n697), .B2(new_n854), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n913), .A2(new_n853), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n885), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n596), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n912), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n524), .A2(KEYINPUT57), .ZN(new_n920));
  AOI22_X1  g719(.A1(new_n909), .A2(KEYINPUT57), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n660), .A3(new_n891), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(new_n924));
  OR3_X1    g723(.A1(new_n924), .A2(KEYINPUT59), .A3(new_n693), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n908), .A2(new_n923), .A3(new_n925), .ZN(G1345gat));
  OAI21_X1  g725(.A(G155gat), .B1(new_n924), .B2(new_n596), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n749), .A2(new_n587), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n905), .B2(new_n928), .ZN(G1346gat));
  OAI21_X1  g728(.A(G162gat), .B1(new_n924), .B2(new_n697), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n697), .A2(G162gat), .A3(new_n424), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n894), .A2(new_n895), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(G1347gat));
  NAND2_X1  g732(.A1(new_n666), .A2(new_n424), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n934), .A2(new_n567), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n862), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n864), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n660), .ZN(new_n939));
  XOR2_X1   g738(.A(KEYINPUT123), .B(G176gat), .Z(new_n940));
  XNOR2_X1  g739(.A(new_n939), .B(new_n940), .ZN(G1349gat));
  INV_X1    g740(.A(G183gat), .ZN(new_n942));
  INV_X1    g741(.A(new_n935), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n904), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n942), .B1(new_n944), .B2(new_n596), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT60), .ZN(new_n946));
  INV_X1    g745(.A(new_n312), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n936), .A2(new_n947), .A3(new_n749), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n946), .B1(new_n945), .B2(new_n948), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n949), .A2(new_n950), .ZN(G1350gat));
  OAI22_X1  g750(.A1(new_n944), .A2(new_n697), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n952));
  NAND2_X1  g751(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n952), .B(new_n953), .ZN(G1351gat));
  NAND3_X1  g753(.A1(new_n666), .A2(new_n424), .A3(new_n381), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n904), .A2(KEYINPUT124), .A3(new_n737), .A4(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n958), .B1(new_n909), .B2(new_n955), .ZN(new_n959));
  INV_X1    g758(.A(G197gat), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n957), .A2(new_n959), .A3(new_n960), .A4(new_n864), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n921), .A2(new_n864), .A3(new_n956), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n962), .B2(new_n960), .ZN(G1352gat));
  NAND2_X1  g762(.A1(new_n909), .A2(KEYINPUT57), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n919), .A2(new_n920), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n964), .A2(new_n660), .A3(new_n965), .A4(new_n956), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n921), .A2(KEYINPUT126), .A3(new_n660), .A4(new_n956), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n968), .A2(G204gat), .A3(new_n969), .ZN(new_n970));
  AOI211_X1 g769(.A(G204gat), .B(new_n693), .C1(KEYINPUT125), .C2(KEYINPUT62), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n904), .A2(new_n737), .A3(new_n956), .A4(new_n971), .ZN(new_n972));
  NOR2_X1   g771(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n973));
  XNOR2_X1  g772(.A(new_n972), .B(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n970), .A2(new_n974), .ZN(G1353gat));
  NAND4_X1  g774(.A1(new_n957), .A2(new_n959), .A3(new_n383), .A4(new_n749), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n964), .A2(new_n749), .A3(new_n965), .A4(new_n956), .ZN(new_n977));
  AND3_X1   g776(.A1(new_n977), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n978));
  AOI21_X1  g777(.A(KEYINPUT63), .B1(new_n977), .B2(G211gat), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(G1354gat));
  AND2_X1   g779(.A1(new_n921), .A2(new_n956), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n640), .A2(G218gat), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(KEYINPUT127), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n957), .A2(new_n640), .A3(new_n959), .ZN(new_n984));
  AOI22_X1  g783(.A1(new_n981), .A2(new_n983), .B1(new_n984), .B2(new_n384), .ZN(G1355gat));
endmodule


