//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1033, new_n1034, new_n1035,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091,
    new_n1092, new_n1093, new_n1094, new_n1095, new_n1096, new_n1097,
    new_n1098, new_n1099, new_n1100, new_n1101, new_n1102;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G469), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G137), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT11), .A3(G134), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(G137), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G131), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n196), .A2(new_n198), .A3(new_n202), .A4(new_n199), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  OR2_X1    g018(.A1(KEYINPUT84), .A2(KEYINPUT12), .ZN(new_n205));
  INV_X1    g019(.A(G101), .ZN(new_n206));
  INV_X1    g020(.A(G107), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G104), .ZN(new_n208));
  INV_X1    g022(.A(G104), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G107), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n206), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT82), .ZN(new_n212));
  OR2_X1    g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT3), .B1(new_n209), .B2(G107), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(new_n207), .A3(G104), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n214), .A2(new_n216), .A3(new_n206), .A4(new_n210), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n211), .A2(new_n212), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n213), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT65), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G146), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n221), .A2(new_n223), .A3(G143), .ZN(new_n224));
  INV_X1    g038(.A(G143), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT64), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G143), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(new_n228), .A3(G146), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT1), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n224), .A2(new_n229), .A3(new_n230), .A4(G128), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n224), .A2(new_n229), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n226), .A2(new_n228), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n230), .B1(new_n234), .B2(new_n220), .ZN(new_n235));
  INV_X1    g049(.A(G128), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n233), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT83), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n232), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT64), .B(G143), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT1), .B1(new_n240), .B2(G146), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n241), .A2(G128), .B1(new_n224), .B2(new_n229), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT83), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n219), .B1(new_n239), .B2(new_n243), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n213), .A2(new_n217), .A3(new_n218), .ZN(new_n245));
  AOI21_X1  g059(.A(G146), .B1(new_n226), .B2(new_n228), .ZN(new_n246));
  AOI21_X1  g060(.A(G143), .B1(new_n221), .B2(new_n223), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n236), .B1(new_n224), .B2(KEYINPUT1), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n231), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n204), .B(new_n205), .C1(new_n244), .C2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n204), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n231), .B1(new_n242), .B2(KEYINPUT83), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n237), .A2(new_n238), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n245), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n250), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n219), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n253), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  XOR2_X1   g073(.A(KEYINPUT84), .B(KEYINPUT12), .Z(new_n260));
  OAI21_X1  g074(.A(new_n252), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT85), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n214), .A2(new_n216), .A3(new_n210), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G101), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(KEYINPUT4), .A3(new_n217), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT80), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AND2_X1   g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  NOR2_X1   g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  OR2_X1    g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n234), .A2(new_n220), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n222), .A2(G146), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n220), .A2(KEYINPUT65), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n225), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n270), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n224), .A2(new_n229), .A3(new_n268), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n264), .A2(KEYINPUT80), .A3(KEYINPUT4), .A4(new_n217), .ZN(new_n278));
  OR2_X1    g092(.A1(new_n264), .A2(KEYINPUT4), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n267), .A2(new_n277), .A3(new_n278), .A4(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT81), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n264), .A2(KEYINPUT4), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(new_n266), .B2(new_n265), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n284), .A2(KEYINPUT81), .A3(new_n277), .A4(new_n278), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT10), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n287), .B(new_n245), .C1(new_n254), .C2(new_n255), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT10), .B1(new_n257), .B2(new_n219), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n286), .A2(new_n290), .A3(new_n253), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n261), .A2(new_n262), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(G110), .B(G140), .ZN(new_n293));
  INV_X1    g107(.A(G953), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n294), .A2(G227), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n293), .B(new_n295), .ZN(new_n296));
  XOR2_X1   g110(.A(new_n296), .B(KEYINPUT79), .Z(new_n297));
  NAND2_X1  g111(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n262), .B1(new_n261), .B2(new_n291), .ZN(new_n299));
  INV_X1    g113(.A(new_n296), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n291), .A2(KEYINPUT86), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n286), .A2(new_n290), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n204), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT86), .B1(new_n291), .B2(new_n300), .ZN(new_n305));
  OAI22_X1  g119(.A1(new_n298), .A2(new_n299), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n193), .B1(new_n306), .B2(new_n190), .ZN(new_n307));
  XOR2_X1   g121(.A(KEYINPUT87), .B(G469), .Z(new_n308));
  NAND3_X1  g122(.A1(new_n261), .A2(new_n291), .A3(new_n300), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n300), .B1(new_n303), .B2(new_n291), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n190), .B(new_n308), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n192), .B1(new_n307), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT88), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT88), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n316), .B(new_n192), .C1(new_n307), .C2(new_n313), .ZN(new_n317));
  INV_X1    g131(.A(G217), .ZN(new_n318));
  NOR3_X1   g132(.A1(new_n188), .A2(new_n318), .A3(G953), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n240), .A2(G128), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n236), .A2(G143), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n195), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n321), .A2(new_n195), .A3(new_n322), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G116), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT95), .B1(new_n327), .B2(G122), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT95), .ZN(new_n329));
  INV_X1    g143(.A(G122), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(G116), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n327), .A2(G122), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n207), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(KEYINPUT14), .ZN(new_n335));
  OR3_X1    g149(.A1(new_n330), .A2(KEYINPUT14), .A3(G116), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n332), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G107), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(KEYINPUT96), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT96), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n340), .B1(new_n337), .B2(G107), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n326), .B(new_n334), .C1(new_n339), .C2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT97), .ZN(new_n343));
  INV_X1    g157(.A(new_n334), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n207), .B1(new_n332), .B2(new_n333), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n321), .A2(new_n322), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT13), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(G134), .B1(new_n321), .B2(KEYINPUT13), .ZN(new_n349));
  OAI221_X1 g163(.A(new_n325), .B1(new_n344), .B2(new_n345), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n342), .A2(new_n343), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n343), .B1(new_n342), .B2(new_n350), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n320), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n325), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n334), .B1(new_n354), .B2(new_n323), .ZN(new_n355));
  INV_X1    g169(.A(new_n339), .ZN(new_n356));
  INV_X1    g170(.A(new_n341), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n348), .A2(new_n349), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n325), .B1(new_n344), .B2(new_n345), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT97), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n342), .A2(new_n350), .A3(new_n343), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n363), .A3(new_n319), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n353), .A2(new_n364), .A3(new_n190), .ZN(new_n365));
  INV_X1    g179(.A(G478), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(KEYINPUT15), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n367), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n353), .A2(new_n364), .A3(new_n190), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(G234), .A2(G237), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(G952), .A3(new_n294), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT21), .B(G898), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n372), .A2(G902), .A3(G953), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  XOR2_X1   g191(.A(new_n377), .B(KEYINPUT98), .Z(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n371), .A2(new_n379), .ZN(new_n380));
  AND2_X1   g194(.A1(KEYINPUT69), .A2(G237), .ZN(new_n381));
  NOR2_X1   g195(.A1(KEYINPUT69), .A2(G237), .ZN(new_n382));
  OAI211_X1 g196(.A(G214), .B(new_n294), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n240), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT69), .B(G237), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n385), .A2(G143), .A3(G214), .A4(new_n294), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n202), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT17), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT92), .B1(new_n387), .B2(G131), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT92), .ZN(new_n392));
  AOI211_X1 g206(.A(new_n392), .B(new_n202), .C1(new_n384), .C2(new_n386), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n389), .B(new_n390), .C1(new_n391), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n387), .A2(G131), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n392), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n387), .A2(KEYINPUT92), .A3(G131), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(KEYINPUT17), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G125), .ZN(new_n399));
  NOR3_X1   g213(.A1(new_n399), .A2(KEYINPUT16), .A3(G140), .ZN(new_n400));
  XNOR2_X1  g214(.A(G125), .B(G140), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n400), .B1(new_n401), .B2(KEYINPUT16), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT74), .B1(new_n402), .B2(G146), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(G146), .B2(new_n402), .ZN(new_n404));
  INV_X1    g218(.A(new_n402), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(KEYINPUT74), .A3(new_n220), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n394), .A2(new_n398), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT65), .B(G146), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n401), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n410), .B1(new_n220), .B2(new_n401), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT18), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(new_n202), .ZN(new_n413));
  OAI221_X1 g227(.A(new_n411), .B1(new_n387), .B2(new_n413), .C1(new_n395), .C2(new_n412), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(G113), .B(G122), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(new_n209), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n408), .A2(new_n417), .A3(new_n414), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n190), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G475), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT94), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n408), .A2(new_n417), .A3(new_n414), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n389), .B1(new_n391), .B2(new_n393), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n402), .A2(G146), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT93), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n401), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(KEYINPUT19), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n409), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n426), .A2(new_n427), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n417), .B1(new_n433), .B2(new_n414), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n424), .B1(new_n425), .B2(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(G475), .A2(G902), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n433), .A2(new_n414), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n418), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n420), .A3(KEYINPUT94), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n435), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n440), .A2(KEYINPUT20), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n436), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(new_n438), .B2(new_n420), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n380), .B(new_n423), .C1(new_n441), .C2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT2), .B(G113), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT67), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G113), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT2), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT2), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G113), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n450), .A2(new_n452), .A3(new_n447), .ZN(new_n453));
  XNOR2_X1  g267(.A(G116), .B(G119), .ZN(new_n454));
  OAI22_X1  g268(.A1(new_n448), .A2(new_n453), .B1(KEYINPUT66), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n454), .A2(KEYINPUT66), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n450), .A2(new_n452), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT67), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n446), .A2(new_n447), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n456), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n267), .A2(new_n461), .A3(new_n278), .A4(new_n279), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n457), .A2(new_n454), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT5), .ZN(new_n464));
  INV_X1    g278(.A(G119), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n464), .A2(new_n465), .A3(G116), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT89), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n449), .B1(new_n454), .B2(KEYINPUT5), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n245), .A2(new_n463), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n462), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT6), .ZN(new_n472));
  XNOR2_X1  g286(.A(G110), .B(G122), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n471), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n462), .A2(new_n470), .A3(new_n473), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT6), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n473), .B1(new_n462), .B2(new_n470), .ZN(new_n478));
  OAI211_X1 g292(.A(KEYINPUT90), .B(new_n475), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n478), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT90), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT6), .A4(new_n476), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n230), .B1(new_n409), .B2(G143), .ZN(new_n484));
  OAI22_X1  g298(.A1(new_n484), .A2(new_n236), .B1(new_n246), .B2(new_n247), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(new_n399), .A3(new_n231), .ZN(new_n486));
  OAI21_X1  g300(.A(G125), .B1(new_n275), .B2(new_n276), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G224), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n489), .A2(G953), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(KEYINPUT91), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n488), .B(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n483), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(G210), .B1(G237), .B2(G902), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n469), .A2(new_n463), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n219), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n470), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n473), .B(KEYINPUT8), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT7), .B1(new_n489), .B2(G953), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n488), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n488), .A2(new_n500), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n499), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n476), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n190), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n493), .A2(new_n494), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n494), .ZN(new_n508));
  INV_X1    g322(.A(new_n492), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n509), .B1(new_n479), .B2(new_n482), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n508), .B1(new_n510), .B2(new_n505), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(G214), .B1(G237), .B2(G902), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n445), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n315), .A2(new_n317), .A3(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(G472), .A2(G902), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n455), .A2(new_n460), .ZN(new_n518));
  INV_X1    g332(.A(new_n199), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n195), .A2(G137), .ZN(new_n520));
  OAI21_X1  g334(.A(G131), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n203), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n250), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT68), .B1(new_n277), .B2(new_n204), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n268), .A2(new_n269), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n526), .B1(new_n246), .B2(new_n247), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n224), .A2(new_n229), .A3(new_n268), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n204), .A2(KEYINPUT68), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n518), .B(new_n524), .C1(new_n525), .C2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n385), .A2(G210), .A3(new_n294), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n532), .B(KEYINPUT27), .ZN(new_n533));
  XNOR2_X1  g347(.A(KEYINPUT26), .B(G101), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n533), .B(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT30), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n204), .A2(new_n527), .A3(new_n528), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n524), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n524), .B1(new_n525), .B2(new_n530), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n538), .B1(new_n539), .B2(KEYINPUT30), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n531), .B(new_n535), .C1(new_n540), .C2(new_n518), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT70), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n524), .A2(new_n536), .A3(new_n537), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n522), .B1(new_n485), .B2(new_n231), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT68), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n537), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n544), .B1(new_n546), .B2(new_n529), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n543), .B1(new_n547), .B2(new_n536), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n461), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT70), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n549), .A2(new_n550), .A3(new_n531), .A4(new_n535), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n542), .A2(KEYINPUT31), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n535), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n524), .A2(new_n518), .A3(new_n537), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT28), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n518), .B1(new_n524), .B2(new_n537), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n555), .B1(new_n531), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT71), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n556), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n557), .B1(new_n547), .B2(new_n518), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n562), .A2(KEYINPUT71), .A3(new_n555), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n553), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  AOI211_X1 g378(.A(new_n461), .B(new_n544), .C1(new_n546), .C2(new_n529), .ZN(new_n565));
  AOI211_X1 g379(.A(new_n553), .B(new_n565), .C1(new_n548), .C2(new_n461), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT31), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n517), .B1(new_n552), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT32), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT71), .B1(new_n562), .B2(new_n555), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n560), .B(KEYINPUT28), .C1(new_n565), .C2(new_n557), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n574), .A3(new_n556), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n553), .A2(new_n575), .B1(new_n566), .B2(new_n567), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n542), .A2(KEYINPUT31), .A3(new_n551), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n578), .A2(KEYINPUT32), .A3(new_n517), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n549), .A2(new_n531), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n553), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT29), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n581), .B(new_n582), .C1(new_n575), .C2(new_n553), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n546), .A2(new_n529), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n518), .B1(new_n584), .B2(new_n524), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT28), .B1(new_n565), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n556), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n553), .A2(new_n582), .ZN(new_n589));
  AOI21_X1  g403(.A(G902), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n583), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G472), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n572), .A2(new_n579), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT25), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT23), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(new_n465), .B2(G128), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT72), .B1(new_n465), .B2(G128), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT73), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n598), .A2(KEYINPUT73), .A3(new_n599), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(new_n603), .A3(G110), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT24), .B(G110), .Z(new_n605));
  XNOR2_X1  g419(.A(G119), .B(G128), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n604), .A2(new_n406), .A3(new_n404), .A4(new_n607), .ZN(new_n608));
  OAI22_X1  g422(.A1(new_n600), .A2(G110), .B1(new_n606), .B2(new_n605), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(new_n427), .A3(new_n410), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT22), .B(G137), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n294), .A2(G221), .A3(G234), .ZN(new_n613));
  XOR2_X1   g427(.A(new_n612), .B(new_n613), .Z(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n608), .A2(new_n610), .A3(new_n614), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n594), .B1(new_n618), .B2(G902), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n616), .A2(KEYINPUT25), .A3(new_n190), .A4(new_n617), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n318), .B1(G234), .B2(new_n190), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(G902), .ZN(new_n624));
  XOR2_X1   g438(.A(new_n624), .B(KEYINPUT75), .Z(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n616), .A2(new_n617), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(new_n627), .B(KEYINPUT76), .Z(new_n628));
  INV_X1    g442(.A(KEYINPUT77), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n623), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n622), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n631), .B1(new_n619), .B2(new_n620), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n627), .B(KEYINPUT76), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT77), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n593), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT78), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n593), .A2(KEYINPUT78), .A3(new_n636), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n516), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(new_n206), .ZN(G3));
  INV_X1    g456(.A(new_n317), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n261), .A2(new_n291), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT85), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(new_n292), .A3(new_n297), .ZN(new_n646));
  INV_X1    g460(.A(new_n305), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(new_n303), .A3(new_n301), .ZN(new_n648));
  AOI21_X1  g462(.A(G902), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n312), .B1(new_n649), .B2(new_n193), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n316), .B1(new_n650), .B2(new_n192), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n643), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n512), .A2(new_n513), .A3(new_n378), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n444), .B1(new_n440), .B2(KEYINPUT20), .ZN(new_n654));
  INV_X1    g468(.A(new_n423), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n366), .A2(G902), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT100), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n353), .A2(new_n364), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT33), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n353), .A2(new_n364), .A3(new_n658), .A4(KEYINPUT33), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n657), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n365), .A2(new_n366), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  OAI22_X1  g479(.A1(new_n654), .A2(new_n655), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n653), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(KEYINPUT99), .A2(G472), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n578), .B2(new_n190), .ZN(new_n669));
  INV_X1    g483(.A(new_n668), .ZN(new_n670));
  AOI211_X1 g484(.A(G902), .B(new_n670), .C1(new_n576), .C2(new_n577), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n635), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n652), .A2(new_n667), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G104), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT101), .B(KEYINPUT34), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G6));
  INV_X1    g490(.A(new_n513), .ZN(new_n677));
  AOI211_X1 g491(.A(new_n677), .B(new_n379), .C1(new_n507), .C2(new_n511), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n440), .A2(KEYINPUT20), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n440), .A2(KEYINPUT102), .A3(KEYINPUT20), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n425), .A2(new_n424), .A3(new_n434), .ZN(new_n683));
  AOI21_X1  g497(.A(KEYINPUT94), .B1(new_n438), .B2(new_n420), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n683), .A2(new_n684), .A3(new_n443), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n681), .A2(new_n682), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n371), .A2(new_n423), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n678), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n652), .A2(new_n672), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n207), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT103), .B(KEYINPUT35), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G9));
  NOR2_X1   g508(.A1(new_n615), .A2(KEYINPUT36), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n611), .B(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n632), .B1(new_n626), .B2(new_n696), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n669), .A2(new_n671), .A3(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n315), .A2(new_n698), .A3(new_n317), .A4(new_n515), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT37), .B(G110), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G12));
  XNOR2_X1  g515(.A(new_n373), .B(KEYINPUT104), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n702), .B1(G900), .B2(new_n376), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n704));
  OR2_X1    g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n703), .A2(new_n704), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n685), .B1(new_n679), .B2(new_n680), .ZN(new_n709));
  AOI211_X1 g523(.A(new_n688), .B(new_n708), .C1(new_n709), .C2(new_n682), .ZN(new_n710));
  INV_X1    g524(.A(new_n514), .ZN(new_n711));
  INV_X1    g525(.A(new_n697), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n710), .A2(new_n593), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n315), .A2(new_n317), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(new_n236), .ZN(G30));
  XNOR2_X1  g530(.A(new_n707), .B(KEYINPUT39), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n315), .A2(new_n317), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT40), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n513), .B(new_n371), .C1(new_n654), .C2(new_n655), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n507), .A2(KEYINPUT38), .A3(new_n511), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT38), .B1(new_n507), .B2(new_n511), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n553), .B1(new_n565), .B2(new_n585), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n542), .A2(new_n551), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n190), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(G472), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n572), .A2(new_n579), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n723), .A2(new_n728), .A3(new_n697), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT40), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n315), .A2(new_n732), .A3(new_n317), .A4(new_n717), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n723), .A2(new_n728), .A3(KEYINPUT106), .A4(new_n697), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n719), .A2(new_n731), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n234), .ZN(G45));
  NOR2_X1   g550(.A1(new_n666), .A2(new_n708), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n593), .A2(new_n711), .A3(new_n737), .A4(new_n712), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n714), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n220), .ZN(G48));
  NAND2_X1  g554(.A1(new_n303), .A2(new_n291), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n296), .ZN(new_n742));
  AOI21_X1  g556(.A(G902), .B1(new_n742), .B2(new_n309), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n192), .B(new_n312), .C1(new_n743), .C2(new_n193), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n593), .A2(new_n667), .A3(new_n636), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT41), .B(G113), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G15));
  NAND4_X1  g562(.A1(new_n690), .A2(new_n593), .A3(new_n636), .A4(new_n745), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G116), .ZN(G18));
  INV_X1    g564(.A(new_n445), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n514), .A2(new_n744), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n593), .A2(new_n751), .A3(new_n712), .A4(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G119), .ZN(G21));
  INV_X1    g568(.A(new_n512), .ZN(new_n755));
  NOR4_X1   g569(.A1(new_n720), .A2(new_n744), .A3(new_n755), .A4(new_n379), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n190), .B1(new_n552), .B2(new_n569), .ZN(new_n757));
  AOI22_X1  g571(.A1(new_n566), .A2(new_n567), .B1(new_n587), .B2(new_n553), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n577), .A2(new_n758), .ZN(new_n759));
  AOI22_X1  g573(.A1(new_n757), .A2(G472), .B1(new_n517), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n632), .A2(new_n633), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT107), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n759), .A2(new_n517), .ZN(new_n763));
  AOI21_X1  g577(.A(G902), .B1(new_n576), .B2(new_n577), .ZN(new_n764));
  INV_X1    g578(.A(G472), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n763), .B(new_n761), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT107), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n756), .B1(new_n762), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G122), .ZN(G24));
  NAND2_X1  g584(.A1(new_n757), .A2(G472), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n771), .A2(new_n712), .A3(new_n763), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n737), .A3(new_n752), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G125), .ZN(G27));
  NAND3_X1  g588(.A1(new_n593), .A2(new_n761), .A3(new_n737), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n507), .A2(new_n511), .A3(new_n513), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n650), .A2(new_n192), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT42), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT32), .B1(new_n578), .B2(new_n517), .ZN(new_n780));
  INV_X1    g594(.A(new_n517), .ZN(new_n781));
  AOI211_X1 g595(.A(new_n571), .B(new_n781), .C1(new_n576), .C2(new_n577), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n635), .B1(new_n783), .B2(new_n592), .ZN(new_n784));
  INV_X1    g598(.A(new_n778), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n661), .A2(new_n662), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n656), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n664), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n788), .B(new_n707), .C1(new_n654), .C2(new_n655), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(KEYINPUT42), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n784), .A2(new_n785), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n779), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(new_n202), .ZN(G33));
  NAND3_X1  g607(.A1(new_n687), .A2(new_n689), .A3(new_n707), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT108), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n708), .B1(new_n709), .B2(new_n682), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT108), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n797), .A3(new_n689), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n784), .A2(new_n785), .A3(new_n795), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G134), .ZN(G36));
  NOR2_X1   g614(.A1(new_n654), .A2(new_n655), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT110), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n788), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT43), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n801), .B(new_n788), .C1(new_n802), .C2(KEYINPUT43), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT111), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n757), .A2(new_n670), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n764), .A2(new_n668), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n809), .B1(new_n812), .B2(new_n712), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n809), .B(new_n712), .C1(new_n669), .C2(new_n671), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n808), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT44), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n717), .A2(new_n192), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT45), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n306), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n646), .A2(new_n648), .A3(KEYINPUT45), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(G469), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n193), .A2(new_n190), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n823), .A2(KEYINPUT46), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT109), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n193), .B1(new_n306), .B2(new_n820), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n824), .B1(new_n829), .B2(new_n822), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(KEYINPUT109), .A3(KEYINPUT46), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n823), .A2(new_n825), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT46), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n313), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n819), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n808), .B(KEYINPUT44), .C1(new_n813), .C2(new_n815), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n818), .A2(new_n777), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(G137), .ZN(G39));
  OAI21_X1  g653(.A(new_n312), .B1(new_n830), .B2(KEYINPUT46), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n828), .B2(new_n831), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT47), .B1(new_n841), .B2(new_n191), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n826), .A2(new_n827), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT109), .B1(new_n830), .B2(KEYINPUT46), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n835), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT47), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n845), .A2(new_n846), .A3(new_n192), .ZN(new_n847));
  NOR4_X1   g661(.A1(new_n593), .A2(new_n789), .A3(new_n636), .A4(new_n776), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n842), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(G140), .ZN(G42));
  INV_X1    g664(.A(new_n804), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n851), .A2(new_n761), .A3(new_n192), .A4(new_n513), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT112), .ZN(new_n853));
  INV_X1    g667(.A(new_n728), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n721), .A2(new_n722), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n743), .A2(new_n193), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n313), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT49), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n697), .B1(new_n783), .B2(new_n592), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n776), .A2(new_n655), .A3(new_n371), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n796), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n860), .A2(new_n315), .A3(new_n862), .A4(new_n317), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n306), .A2(new_n190), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(G469), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n191), .B1(new_n865), .B2(new_n312), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n772), .A2(new_n866), .A3(new_n737), .A4(new_n777), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n799), .A2(new_n863), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n792), .B1(new_n868), .B2(KEYINPUT113), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n769), .A2(new_n746), .A3(new_n749), .A4(new_n753), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n423), .B(new_n371), .C1(new_n441), .C2(new_n444), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n653), .B1(new_n871), .B2(new_n666), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n672), .A2(new_n315), .A3(new_n872), .A4(new_n317), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n699), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n870), .A2(new_n641), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT113), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n799), .A2(new_n863), .A3(new_n876), .A4(new_n867), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n869), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT114), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT52), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n773), .B1(new_n713), .B2(new_n714), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n707), .B(KEYINPUT116), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n720), .A2(new_n755), .A3(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n883), .A2(new_n728), .A3(new_n866), .A4(new_n697), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n884), .B1(new_n738), .B2(new_n714), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n880), .B1(new_n881), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT115), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n881), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n739), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n773), .B(KEYINPUT115), .C1(new_n713), .C2(new_n714), .ZN(new_n890));
  NOR4_X1   g704(.A1(new_n314), .A2(new_n755), .A3(new_n720), .A4(new_n882), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n712), .B1(new_n783), .B2(new_n727), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n880), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n888), .A2(new_n889), .A3(new_n890), .A4(new_n893), .ZN(new_n894));
  AOI22_X1  g708(.A1(new_n878), .A2(new_n879), .B1(new_n886), .B2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n869), .A2(new_n875), .A3(KEYINPUT114), .A4(new_n877), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT53), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n873), .A2(new_n699), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n315), .A2(new_n317), .A3(new_n515), .ZN(new_n899));
  INV_X1    g713(.A(new_n640), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT78), .B1(new_n593), .B2(new_n636), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n593), .A2(new_n636), .A3(new_n745), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n766), .A2(new_n767), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n771), .A2(KEYINPUT107), .A3(new_n761), .A4(new_n763), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI22_X1  g720(.A1(new_n903), .A2(new_n690), .B1(new_n906), .B2(new_n756), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n746), .A2(new_n753), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n898), .A2(new_n902), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  AND4_X1   g723(.A1(new_n876), .A2(new_n799), .A3(new_n863), .A4(new_n867), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AND4_X1   g725(.A1(new_n712), .A2(new_n737), .A3(new_n752), .A4(new_n760), .ZN(new_n912));
  AND4_X1   g726(.A1(new_n593), .A2(new_n710), .A3(new_n711), .A4(new_n712), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n912), .B1(new_n913), .B2(new_n652), .ZN(new_n914));
  AND4_X1   g728(.A1(new_n593), .A2(new_n711), .A3(new_n737), .A4(new_n712), .ZN(new_n915));
  AOI22_X1  g729(.A1(new_n915), .A2(new_n652), .B1(new_n891), .B2(new_n892), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n914), .A2(new_n916), .A3(KEYINPUT52), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n886), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n911), .A2(KEYINPUT53), .A3(new_n918), .A4(new_n869), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT117), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND4_X1   g735(.A1(new_n746), .A2(new_n769), .A3(new_n749), .A4(new_n753), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n922), .A2(new_n877), .A3(new_n902), .A4(new_n898), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n795), .A2(new_n798), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n593), .A2(new_n866), .A3(new_n636), .A4(new_n777), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n867), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n593), .A2(new_n712), .A3(new_n796), .A4(new_n861), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n927), .A2(new_n714), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT113), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n792), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n923), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n932), .A2(KEYINPUT117), .A3(KEYINPUT53), .A4(new_n918), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n921), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT54), .B1(new_n897), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n894), .A2(new_n886), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n932), .A2(KEYINPUT53), .A3(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT53), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n917), .A2(new_n886), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n938), .B1(new_n878), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT54), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n937), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n935), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n702), .B1(new_n806), .B2(new_n807), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n744), .A2(new_n776), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n944), .A2(new_n772), .A3(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n635), .A2(new_n373), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n854), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n801), .A2(new_n664), .A3(new_n787), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n944), .A2(new_n906), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n951), .A2(new_n677), .A3(new_n855), .A4(new_n745), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT50), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n952), .A2(new_n953), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n950), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI22_X1  g770(.A1(new_n842), .A2(new_n847), .B1(new_n191), .B2(new_n857), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n951), .A2(new_n777), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT51), .ZN(new_n961));
  OAI21_X1  g775(.A(KEYINPUT118), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT118), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n956), .A2(new_n963), .A3(KEYINPUT51), .A4(new_n959), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n960), .A2(new_n961), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n593), .A2(new_n761), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n944), .A2(new_n966), .A3(new_n945), .ZN(new_n967));
  AND2_X1   g781(.A1(KEYINPUT119), .A2(KEYINPUT48), .ZN(new_n968));
  NOR2_X1   g782(.A1(KEYINPUT119), .A2(KEYINPUT48), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n967), .A2(new_n968), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n951), .A2(new_n752), .ZN(new_n972));
  OAI211_X1 g786(.A(G952), .B(new_n294), .C1(new_n948), .C2(new_n666), .ZN(new_n973));
  NOR4_X1   g787(.A1(new_n970), .A2(new_n971), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n962), .A2(new_n964), .A3(new_n965), .A4(new_n974), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n943), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(G952), .A2(G953), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n859), .B1(new_n976), .B2(new_n977), .ZN(G75));
  XNOR2_X1  g792(.A(new_n483), .B(new_n492), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT55), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n190), .B1(new_n937), .B2(new_n940), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n981), .A2(G210), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n980), .B1(new_n982), .B2(KEYINPUT56), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n294), .A2(G952), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n982), .A2(KEYINPUT56), .A3(new_n980), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n986), .A2(new_n987), .ZN(G51));
  AOI21_X1  g802(.A(KEYINPUT53), .B1(new_n932), .B2(new_n918), .ZN(new_n989));
  INV_X1    g803(.A(new_n936), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n869), .A2(new_n875), .A3(KEYINPUT53), .A4(new_n877), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(KEYINPUT54), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n993), .A2(KEYINPUT120), .A3(new_n942), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n937), .A2(new_n940), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT120), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n995), .A2(new_n996), .A3(KEYINPUT54), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n824), .B(KEYINPUT57), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n994), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n742), .A2(new_n309), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n981), .A2(new_n822), .A3(new_n829), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n984), .B1(new_n1001), .B2(new_n1002), .ZN(G54));
  NOR2_X1   g817(.A1(new_n683), .A2(new_n684), .ZN(new_n1004));
  AND2_X1   g818(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n981), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1004), .B1(new_n981), .B2(new_n1005), .ZN(new_n1007));
  NOR3_X1   g821(.A1(new_n1006), .A2(new_n1007), .A3(new_n984), .ZN(G60));
  XOR2_X1   g822(.A(new_n786), .B(KEYINPUT121), .Z(new_n1009));
  NAND2_X1  g823(.A1(G478), .A2(G902), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1010), .B(KEYINPUT59), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1009), .B1(new_n943), .B2(new_n1011), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n994), .A2(new_n997), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(new_n985), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1012), .A2(new_n1015), .ZN(G63));
  INV_X1    g830(.A(KEYINPUT61), .ZN(new_n1017));
  OR2_X1    g831(.A1(new_n1017), .A2(KEYINPUT122), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(KEYINPUT122), .ZN(new_n1019));
  NAND2_X1  g833(.A1(G217), .A2(G902), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT60), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1021), .B1(new_n937), .B2(new_n940), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(new_n696), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(new_n618), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n985), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  OAI211_X1 g840(.A(new_n1018), .B(new_n1019), .C1(new_n1024), .C2(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1021), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n995), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n984), .B1(new_n1029), .B2(new_n618), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n1030), .A2(KEYINPUT122), .A3(new_n1017), .A4(new_n1023), .ZN(new_n1031));
  AND2_X1   g845(.A1(new_n1027), .A2(new_n1031), .ZN(G66));
  OAI21_X1  g846(.A(G953), .B1(new_n374), .B2(new_n489), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1033), .B1(new_n875), .B2(G953), .ZN(new_n1034));
  OAI211_X1 g848(.A(new_n479), .B(new_n482), .C1(G898), .C2(new_n294), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1034), .B(new_n1035), .ZN(G69));
  INV_X1    g850(.A(KEYINPUT124), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n739), .B1(new_n881), .B2(new_n887), .ZN(new_n1038));
  AND3_X1   g852(.A1(new_n779), .A2(new_n799), .A3(new_n791), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n838), .A2(new_n890), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  INV_X1    g854(.A(new_n1040), .ZN(new_n1041));
  INV_X1    g855(.A(KEYINPUT123), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n720), .A2(new_n755), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n593), .A2(new_n761), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g858(.A(new_n1044), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n1042), .B1(new_n836), .B2(new_n1045), .ZN(new_n1046));
  NOR4_X1   g860(.A1(new_n841), .A2(KEYINPUT123), .A3(new_n819), .A4(new_n1044), .ZN(new_n1047));
  NOR2_X1   g861(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g862(.A(new_n1048), .ZN(new_n1049));
  NAND4_X1  g863(.A1(new_n1041), .A2(new_n294), .A3(new_n1049), .A4(new_n849), .ZN(new_n1050));
  XNOR2_X1  g864(.A(new_n548), .B(new_n431), .ZN(new_n1051));
  NAND2_X1  g865(.A1(G900), .A2(G953), .ZN(new_n1052));
  AND3_X1   g866(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n639), .A2(new_n640), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n776), .B1(new_n871), .B2(new_n666), .ZN(new_n1055));
  NAND4_X1  g869(.A1(new_n1054), .A2(new_n652), .A3(new_n717), .A4(new_n1055), .ZN(new_n1056));
  AND3_X1   g870(.A1(new_n849), .A2(new_n838), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g871(.A(KEYINPUT62), .ZN(new_n1058));
  NAND4_X1  g872(.A1(new_n1038), .A2(new_n1058), .A3(new_n735), .A4(new_n890), .ZN(new_n1059));
  NAND4_X1  g873(.A1(new_n888), .A2(new_n735), .A3(new_n889), .A4(new_n890), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n1060), .A2(KEYINPUT62), .ZN(new_n1061));
  NAND3_X1  g875(.A1(new_n1057), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g876(.A(new_n1051), .B1(new_n1062), .B2(new_n294), .ZN(new_n1063));
  OAI21_X1  g877(.A(new_n1037), .B1(new_n1053), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g878(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1065));
  AND2_X1   g879(.A1(new_n1062), .A2(new_n294), .ZN(new_n1066));
  OAI211_X1 g880(.A(new_n1065), .B(KEYINPUT124), .C1(new_n1066), .C2(new_n1051), .ZN(new_n1067));
  AOI21_X1  g881(.A(new_n294), .B1(G227), .B2(G900), .ZN(new_n1068));
  NAND3_X1  g882(.A1(new_n1064), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g883(.A(new_n1068), .ZN(new_n1070));
  OAI211_X1 g884(.A(new_n1037), .B(new_n1070), .C1(new_n1053), .C2(new_n1063), .ZN(new_n1071));
  AND2_X1   g885(.A1(new_n1069), .A2(new_n1071), .ZN(G72));
  NAND4_X1  g886(.A1(new_n1057), .A2(new_n875), .A3(new_n1059), .A4(new_n1061), .ZN(new_n1073));
  NAND2_X1  g887(.A1(G472), .A2(G902), .ZN(new_n1074));
  XOR2_X1   g888(.A(new_n1074), .B(KEYINPUT63), .Z(new_n1075));
  NAND2_X1  g889(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g890(.A(KEYINPUT125), .ZN(new_n1077));
  NAND2_X1  g891(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g892(.A1(new_n1073), .A2(KEYINPUT125), .A3(new_n1075), .ZN(new_n1079));
  AOI21_X1  g893(.A(new_n553), .B1(new_n549), .B2(new_n531), .ZN(new_n1080));
  NAND3_X1  g894(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  AND3_X1   g895(.A1(new_n842), .A2(new_n847), .A3(new_n848), .ZN(new_n1082));
  NOR4_X1   g896(.A1(new_n1040), .A2(new_n1048), .A3(new_n1082), .A4(new_n909), .ZN(new_n1083));
  INV_X1    g897(.A(new_n1075), .ZN(new_n1084));
  OAI21_X1  g898(.A(KEYINPUT126), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g899(.A1(new_n1041), .A2(new_n849), .A3(new_n1049), .A4(new_n875), .ZN(new_n1086));
  INV_X1    g900(.A(KEYINPUT126), .ZN(new_n1087));
  NAND3_X1  g901(.A1(new_n1086), .A2(new_n1087), .A3(new_n1075), .ZN(new_n1088));
  NOR2_X1   g902(.A1(new_n580), .A2(new_n535), .ZN(new_n1089));
  NAND3_X1  g903(.A1(new_n1085), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  AND2_X1   g904(.A1(new_n542), .A2(new_n551), .ZN(new_n1091));
  AOI21_X1  g905(.A(new_n1084), .B1(new_n1091), .B2(new_n581), .ZN(new_n1092));
  OAI21_X1  g906(.A(new_n1092), .B1(new_n897), .B2(new_n934), .ZN(new_n1093));
  NAND4_X1  g907(.A1(new_n1081), .A2(new_n1090), .A3(new_n1093), .A4(new_n985), .ZN(new_n1094));
  INV_X1    g908(.A(KEYINPUT127), .ZN(new_n1095));
  NAND2_X1  g909(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g910(.A(new_n879), .B1(new_n923), .B2(new_n931), .ZN(new_n1097));
  NAND3_X1  g911(.A1(new_n1097), .A2(new_n896), .A3(new_n936), .ZN(new_n1098));
  NAND2_X1  g912(.A1(new_n1098), .A2(new_n938), .ZN(new_n1099));
  NAND3_X1  g913(.A1(new_n1099), .A2(new_n921), .A3(new_n933), .ZN(new_n1100));
  AOI21_X1  g914(.A(new_n984), .B1(new_n1100), .B2(new_n1092), .ZN(new_n1101));
  NAND4_X1  g915(.A1(new_n1101), .A2(KEYINPUT127), .A3(new_n1081), .A4(new_n1090), .ZN(new_n1102));
  NAND2_X1  g916(.A1(new_n1096), .A2(new_n1102), .ZN(G57));
endmodule


