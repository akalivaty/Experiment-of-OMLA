//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n792, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n989, new_n990, new_n991;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203));
  INV_X1    g002(.A(G85gat), .ZN(new_n204));
  INV_X1    g003(.A(G92gat), .ZN(new_n205));
  AOI22_X1  g004(.A1(KEYINPUT8), .A2(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT7), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(new_n204), .B2(new_n205), .ZN(new_n208));
  NAND3_X1  g007(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(G99gat), .B(G106gat), .Z(new_n211));
  XOR2_X1   g010(.A(new_n210), .B(new_n211), .Z(new_n212));
  INV_X1    g011(.A(G71gat), .ZN(new_n213));
  INV_X1    g012(.A(G78gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(G71gat), .A2(G78gat), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n215), .B1(KEYINPUT9), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G57gat), .B(G64gat), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n216), .B(KEYINPUT95), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT9), .ZN(new_n221));
  OAI221_X1 g020(.A(new_n220), .B1(new_n221), .B2(new_n218), .C1(new_n213), .C2(new_n214), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n212), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n219), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n210), .B(new_n211), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n202), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(KEYINPUT102), .ZN(new_n228));
  XNOR2_X1  g027(.A(G120gat), .B(G148gat), .ZN(new_n229));
  INV_X1    g028(.A(G176gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G204gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n228), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n223), .A2(KEYINPUT101), .A3(KEYINPUT10), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT101), .B1(new_n224), .B2(new_n225), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT10), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n235), .A2(new_n238), .A3(new_n202), .A4(new_n226), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n227), .A2(KEYINPUT102), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n234), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n239), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n233), .B1(new_n242), .B2(new_n227), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G155gat), .A2(G162gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT2), .ZN(new_n246));
  INV_X1    g045(.A(G141gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n247), .A2(G148gat), .ZN(new_n248));
  INV_X1    g047(.A(G148gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(G141gat), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n246), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  AND2_X1   g050(.A1(G155gat), .A2(G162gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(G155gat), .A2(G162gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT75), .ZN(new_n254));
  NOR3_X1   g053(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G155gat), .ZN(new_n256));
  INV_X1    g055(.A(G162gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT75), .B1(new_n258), .B2(new_n245), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n251), .B1(new_n255), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT76), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n254), .B1(new_n252), .B2(new_n253), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n258), .A2(KEYINPUT75), .A3(new_n245), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT76), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n265), .A3(new_n251), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n258), .A2(new_n245), .ZN(new_n267));
  XNOR2_X1  g066(.A(G141gat), .B(G148gat), .ZN(new_n268));
  OR2_X1    g067(.A1(KEYINPUT77), .A2(G155gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(KEYINPUT77), .A2(G155gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(G162gat), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n268), .B1(new_n271), .B2(KEYINPUT2), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n261), .A2(new_n266), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n274));
  XOR2_X1   g073(.A(G127gat), .B(G134gat), .Z(new_n275));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT1), .ZN(new_n277));
  INV_X1    g076(.A(G113gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n278), .A2(G120gat), .ZN(new_n279));
  INV_X1    g078(.A(G120gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n280), .A2(G113gat), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n276), .B(new_n277), .C1(new_n279), .C2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n275), .B1(new_n282), .B2(KEYINPUT68), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(KEYINPUT68), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n280), .A2(G113gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n278), .A2(G120gat), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT1), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT68), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n284), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n283), .B1(new_n290), .B2(new_n275), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n273), .A2(new_n274), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT79), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n272), .A2(new_n267), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n264), .A2(new_n265), .A3(new_n251), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n265), .B1(new_n264), .B2(new_n251), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n288), .B1(new_n287), .B2(new_n276), .ZN(new_n298));
  AOI211_X1 g097(.A(KEYINPUT68), .B(KEYINPUT1), .C1(new_n285), .C2(new_n286), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n275), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n283), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT4), .B1(new_n297), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT79), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n273), .A2(new_n291), .A3(new_n304), .A4(new_n274), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n293), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT5), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n297), .A2(KEYINPUT3), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT3), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n309), .B(new_n294), .C1(new_n295), .C2(new_n296), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n310), .A3(new_n302), .ZN(new_n311));
  NAND2_X1  g110(.A1(G225gat), .A2(G233gat), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n306), .A2(new_n307), .A3(new_n311), .A4(new_n312), .ZN(new_n313));
  OAI211_X1 g112(.A(KEYINPUT4), .B(new_n312), .C1(new_n297), .C2(new_n302), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(new_n292), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(new_n311), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT78), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n273), .A2(new_n291), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n297), .A2(new_n302), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n312), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n307), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n316), .A2(new_n317), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n317), .B1(new_n316), .B2(new_n322), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n313), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT0), .B(G57gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(G85gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(G1gat), .B(G29gat), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n327), .B(new_n328), .Z(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n329), .B(new_n313), .C1(new_n323), .C2(new_n324), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT6), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT80), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT80), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n331), .A2(new_n332), .A3(new_n336), .A4(new_n333), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n325), .A2(KEYINPUT6), .A3(new_n330), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n340));
  NAND2_X1  g139(.A1(G226gat), .A2(G233gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n341), .B(KEYINPUT72), .Z(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT73), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT67), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT28), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT27), .B(G183gat), .ZN(new_n348));
  INV_X1    g147(.A(G190gat), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AND2_X1   g149(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n349), .B(new_n347), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n346), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  OR3_X1    g154(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n357));
  INV_X1    g156(.A(G169gat), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n356), .B(new_n357), .C1(new_n358), .C2(new_n230), .ZN(new_n359));
  NAND2_X1  g158(.A1(G183gat), .A2(G190gat), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT65), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT24), .ZN(new_n365));
  INV_X1    g164(.A(G183gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n349), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT66), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n366), .A2(new_n349), .A3(KEYINPUT66), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT24), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n360), .A2(new_n363), .A3(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n365), .A2(new_n369), .A3(new_n370), .A4(new_n372), .ZN(new_n373));
  OR3_X1    g172(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n374), .A2(new_n375), .B1(G169gat), .B2(G176gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n373), .A2(KEYINPUT25), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT25), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n367), .A2(KEYINPUT24), .A3(new_n360), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n371), .A2(G183gat), .A3(G190gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n375), .ZN(new_n382));
  NOR3_X1   g181(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n383));
  OAI22_X1  g182(.A1(new_n382), .A2(new_n383), .B1(new_n358), .B2(new_n230), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n378), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n377), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n362), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT29), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n343), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g188(.A1(G211gat), .A2(G218gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(G211gat), .A2(G218gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(G197gat), .A2(G204gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(G197gat), .A2(G204gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n392), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G211gat), .B(G218gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(G197gat), .B(G204gat), .ZN(new_n399));
  INV_X1    g198(.A(new_n396), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n342), .B1(new_n362), .B2(new_n386), .ZN(new_n403));
  NOR3_X1   g202(.A1(new_n389), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n402), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n361), .A2(new_n355), .B1(new_n377), .B2(new_n385), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n342), .B1(new_n406), .B2(KEYINPUT29), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n387), .A2(new_n343), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n340), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT29), .B1(new_n362), .B2(new_n386), .ZN(new_n411));
  OAI221_X1 g210(.A(new_n405), .B1(new_n406), .B2(new_n342), .C1(new_n411), .C2(new_n343), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n387), .A2(new_n388), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n413), .A2(new_n342), .B1(new_n387), .B2(new_n343), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n412), .B(KEYINPUT74), .C1(new_n414), .C2(new_n405), .ZN(new_n415));
  XOR2_X1   g214(.A(G8gat), .B(G36gat), .Z(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(G64gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(new_n205), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n410), .A2(new_n415), .A3(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n412), .B1(new_n414), .B2(new_n405), .ZN(new_n420));
  INV_X1    g219(.A(new_n418), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(KEYINPUT30), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n421), .B1(new_n404), .B2(new_n409), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT30), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n419), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n339), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT86), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT85), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(G50gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(G78gat), .ZN(new_n432));
  XOR2_X1   g231(.A(new_n432), .B(G106gat), .Z(new_n433));
  INV_X1    g232(.A(G228gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n402), .A2(new_n388), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n309), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n297), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT82), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n434), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT3), .B1(new_n402), .B2(new_n388), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n261), .A2(new_n266), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n440), .B1(new_n441), .B2(new_n294), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n402), .B1(new_n310), .B2(new_n388), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n439), .B(G233gat), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n310), .A2(new_n388), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n442), .B1(new_n445), .B2(new_n405), .ZN(new_n446));
  OAI211_X1 g245(.A(G228gat), .B(G233gat), .C1(new_n442), .C2(KEYINPUT82), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  XOR2_X1   g247(.A(KEYINPUT83), .B(G22gat), .Z(new_n449));
  AND3_X1   g248(.A1(new_n444), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n449), .B1(new_n444), .B2(new_n448), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n433), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT84), .ZN(new_n453));
  INV_X1    g252(.A(new_n449), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n446), .A2(new_n447), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n446), .A2(new_n447), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n444), .A2(new_n448), .A3(new_n449), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT84), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(new_n460), .A3(new_n433), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n453), .A2(new_n461), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n444), .A2(G22gat), .A3(new_n448), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n463), .A2(new_n451), .A3(new_n433), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n429), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  AOI211_X1 g265(.A(KEYINPUT85), .B(new_n464), .C1(new_n453), .C2(new_n461), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n428), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n460), .B1(new_n459), .B2(new_n433), .ZN(new_n469));
  INV_X1    g268(.A(new_n433), .ZN(new_n470));
  AOI211_X1 g269(.A(KEYINPUT84), .B(new_n470), .C1(new_n457), .C2(new_n458), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n465), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT85), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n462), .A2(new_n429), .A3(new_n465), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(KEYINPUT86), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n427), .A2(new_n468), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT39), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n320), .A2(new_n321), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n292), .A2(KEYINPUT79), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n305), .A2(new_n303), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n311), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI211_X1 g280(.A(new_n477), .B(new_n478), .C1(new_n481), .C2(new_n321), .ZN(new_n482));
  XOR2_X1   g281(.A(KEYINPUT87), .B(KEYINPUT39), .Z(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n321), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n329), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT40), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n481), .A2(new_n321), .ZN(new_n487));
  INV_X1    g286(.A(new_n478), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(KEYINPUT39), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT40), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n489), .A2(new_n490), .A3(new_n329), .A4(new_n484), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n423), .A2(new_n424), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT30), .B1(new_n420), .B2(new_n421), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n495), .A2(new_n419), .B1(new_n325), .B2(new_n330), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n492), .A2(KEYINPUT88), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT88), .B1(new_n492), .B2(new_n496), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n410), .A2(new_n415), .A3(KEYINPUT37), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n418), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT90), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT37), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n420), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT90), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n500), .A2(new_n505), .A3(new_n418), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n502), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT38), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n389), .A2(new_n405), .A3(new_n403), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n509), .A2(KEYINPUT89), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n414), .A2(new_n402), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(KEYINPUT89), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI211_X1 g312(.A(KEYINPUT38), .B(new_n421), .C1(new_n513), .C2(KEYINPUT37), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n514), .A2(new_n504), .B1(new_n420), .B2(new_n421), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n508), .A2(new_n515), .A3(new_n334), .A4(new_n338), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n473), .A2(new_n474), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n499), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n377), .A2(new_n385), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n359), .A2(new_n360), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n349), .B1(new_n351), .B2(new_n352), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n521), .A2(KEYINPUT67), .A3(KEYINPUT28), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n353), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n520), .B1(new_n523), .B2(new_n346), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n291), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G227gat), .A2(G233gat), .ZN(new_n526));
  XOR2_X1   g325(.A(new_n526), .B(KEYINPUT64), .Z(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n302), .A2(new_n386), .A3(new_n362), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n525), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT32), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT33), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G15gat), .B(G43gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(G71gat), .B(G99gat), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n534), .B(new_n535), .Z(new_n536));
  NAND3_X1  g335(.A1(new_n531), .A2(new_n533), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n525), .A2(new_n529), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n526), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT34), .B1(new_n525), .B2(new_n529), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n539), .A2(KEYINPUT34), .B1(new_n540), .B2(new_n527), .ZN(new_n541));
  INV_X1    g340(.A(new_n536), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n530), .B(KEYINPUT32), .C1(new_n532), .C2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n537), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT71), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT71), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n537), .A2(new_n541), .A3(new_n546), .A4(new_n543), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n537), .A2(new_n543), .ZN(new_n549));
  INV_X1    g348(.A(new_n541), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(KEYINPUT36), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT36), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT70), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n537), .A2(KEYINPUT70), .A3(new_n543), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n550), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n554), .B1(new_n548), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n553), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n476), .A2(new_n518), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT35), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n548), .A2(new_n558), .ZN(new_n563));
  AOI211_X1 g362(.A(new_n562), .B(new_n563), .C1(new_n473), .C2(new_n474), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n339), .A2(new_n426), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n548), .A2(new_n426), .A3(new_n551), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n566), .B1(new_n334), .B2(new_n338), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n567), .B1(new_n466), .B2(new_n467), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n564), .A2(new_n565), .B1(new_n562), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n244), .B1(new_n561), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n571));
  XNOR2_X1  g370(.A(G15gat), .B(G22gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT16), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n573), .A2(G1gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n575), .B1(G1gat), .B2(new_n572), .ZN(new_n576));
  INV_X1    g375(.A(G8gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT21), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n578), .B1(new_n579), .B2(new_n224), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n580), .A2(G183gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(G183gat), .ZN(new_n582));
  INV_X1    g381(.A(G231gat), .ZN(new_n583));
  INV_X1    g382(.A(G233gat), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n581), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n585), .B1(new_n581), .B2(new_n582), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n571), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n588), .ZN(new_n590));
  INV_X1    g389(.A(new_n571), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n590), .A2(new_n586), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n224), .A2(new_n579), .ZN(new_n594));
  XNOR2_X1  g393(.A(G127gat), .B(G155gat), .ZN(new_n595));
  INV_X1    g394(.A(G211gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n594), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n593), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n593), .A2(new_n600), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G134gat), .B(G162gat), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(G29gat), .ZN(new_n606));
  INV_X1    g405(.A(G36gat), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n606), .A2(new_n607), .A3(KEYINPUT14), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT14), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n609), .B1(G29gat), .B2(G36gat), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n608), .B(new_n610), .C1(new_n606), .C2(new_n607), .ZN(new_n611));
  XOR2_X1   g410(.A(KEYINPUT93), .B(G50gat), .Z(new_n612));
  INV_X1    g411(.A(G43gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT94), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n613), .A2(G50gat), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n612), .A2(KEYINPUT94), .A3(new_n613), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT15), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G43gat), .B(G50gat), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT92), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT15), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n611), .B1(new_n621), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n611), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  AND2_X1   g428(.A1(G232gat), .A2(G233gat), .ZN(new_n630));
  AOI22_X1  g429(.A1(new_n629), .A2(new_n212), .B1(KEYINPUT41), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT17), .B1(new_n626), .B2(new_n628), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT17), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n624), .A2(KEYINPUT15), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n634), .B1(new_n620), .B2(new_n619), .ZN(new_n635));
  OAI211_X1 g434(.A(new_n633), .B(new_n627), .C1(new_n635), .C2(new_n611), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n225), .B(KEYINPUT99), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n632), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n631), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(G190gat), .B(G218gat), .Z(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n641), .A2(KEYINPUT100), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n630), .A2(KEYINPUT41), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT98), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(KEYINPUT100), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n639), .A2(new_n642), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n647), .B1(new_n639), .B2(new_n642), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n605), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n650), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n652), .A2(new_n604), .A3(new_n648), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n603), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n627), .B1(new_n635), .B2(new_n611), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n656), .A2(new_n578), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n632), .A2(new_n636), .A3(new_n578), .ZN(new_n658));
  NAND2_X1  g457(.A1(G229gat), .A2(G233gat), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT18), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n656), .B(new_n578), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n659), .B(KEYINPUT13), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n657), .A2(new_n658), .A3(KEYINPUT18), .A4(new_n659), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n662), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(G113gat), .B(G141gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(G169gat), .B(G197gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT12), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n668), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n662), .A2(new_n666), .A3(new_n667), .A4(new_n674), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n655), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n570), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n339), .B(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT104), .B(G1gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1324gat));
  INV_X1    g485(.A(new_n426), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n573), .A2(new_n577), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n570), .A2(new_n687), .A3(new_n680), .A4(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n573), .A2(new_n577), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT42), .B1(new_n691), .B2(KEYINPUT106), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT106), .B1(new_n691), .B2(KEYINPUT105), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI211_X1 g493(.A(KEYINPUT106), .B(KEYINPUT42), .C1(new_n691), .C2(KEYINPUT105), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n681), .A2(new_n687), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n694), .B(new_n695), .C1(new_n577), .C2(new_n696), .ZN(G1325gat));
  INV_X1    g496(.A(new_n552), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n681), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(G15gat), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT107), .B1(new_n553), .B2(new_n559), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n563), .A2(KEYINPUT36), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n702), .B(new_n703), .C1(KEYINPUT36), .C2(new_n552), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(G15gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT108), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n699), .A2(new_n700), .B1(new_n681), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT109), .ZN(G1326gat));
  NAND2_X1  g509(.A1(new_n468), .A2(new_n475), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n681), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(KEYINPUT43), .B(G22gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1327gat));
  NAND2_X1  g514(.A1(new_n561), .A2(new_n569), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n651), .A2(new_n653), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n679), .A2(new_n603), .A3(new_n244), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n719), .A2(new_n606), .A3(new_n683), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT45), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n476), .A2(new_n518), .A3(new_n705), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n569), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n723), .A2(new_n724), .A3(new_n717), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n654), .B1(new_n561), .B2(new_n569), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(new_n683), .A3(new_n718), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n721), .B1(new_n606), .B2(new_n729), .ZN(G1328gat));
  AND2_X1   g529(.A1(new_n719), .A2(new_n607), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT111), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT46), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n731), .A2(new_n732), .A3(new_n733), .A4(new_n687), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n607), .A3(new_n687), .ZN(new_n735));
  OAI21_X1  g534(.A(KEYINPUT111), .B1(new_n735), .B2(KEYINPUT46), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n727), .A2(new_n687), .A3(new_n718), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(G36gat), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT110), .B1(new_n735), .B2(KEYINPUT46), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n735), .A2(KEYINPUT110), .A3(KEYINPUT46), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n737), .B(new_n739), .C1(new_n740), .C2(new_n741), .ZN(G1329gat));
  AOI21_X1  g541(.A(new_n724), .B1(new_n716), .B2(new_n717), .ZN(new_n743));
  AOI211_X1 g542(.A(KEYINPUT44), .B(new_n654), .C1(new_n722), .C2(new_n569), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n706), .B(new_n718), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G43gat), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n719), .A2(KEYINPUT112), .A3(new_n613), .A4(new_n698), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n726), .A2(new_n613), .A3(new_n698), .A4(new_n718), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n746), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT47), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n746), .A2(new_n751), .A3(KEYINPUT47), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(G1330gat));
  INV_X1    g555(.A(new_n517), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n727), .A2(new_n757), .A3(new_n718), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n612), .ZN(new_n759));
  INV_X1    g558(.A(new_n612), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n719), .A2(new_n712), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n759), .A2(KEYINPUT48), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n761), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n727), .A2(new_n712), .A3(new_n718), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n764), .B2(new_n612), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n762), .B1(KEYINPUT48), .B2(new_n765), .ZN(G1331gat));
  NOR2_X1   g565(.A1(new_n655), .A2(new_n678), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n723), .A2(new_n244), .A3(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n683), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XOR2_X1   g569(.A(new_n770), .B(G57gat), .Z(G1332gat));
  INV_X1    g570(.A(new_n244), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(new_n722), .B2(new_n569), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n773), .A2(new_n774), .A3(new_n767), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n774), .B1(new_n773), .B2(new_n767), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  AND2_X1   g577(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n777), .B(new_n687), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n777), .A2(new_n687), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n781), .B2(new_n778), .ZN(G1333gat));
  XNOR2_X1  g581(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n706), .B1(new_n775), .B2(new_n776), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G71gat), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n768), .A2(G71gat), .A3(new_n552), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n783), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n783), .ZN(new_n789));
  AOI211_X1 g588(.A(new_n786), .B(new_n789), .C1(new_n784), .C2(G71gat), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n788), .A2(new_n790), .ZN(G1334gat));
  NAND2_X1  g590(.A1(new_n777), .A2(new_n712), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g592(.A1(new_n603), .A2(new_n678), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n244), .B(new_n794), .C1(new_n743), .C2(new_n744), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n795), .A2(new_n204), .A3(new_n769), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n723), .A2(new_n717), .A3(new_n794), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n654), .B1(new_n722), .B2(new_n569), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n801), .A2(KEYINPUT51), .A3(new_n794), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n799), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT51), .B1(new_n801), .B2(new_n794), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n772), .B1(new_n804), .B2(KEYINPUT115), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n803), .A2(new_n805), .A3(new_n683), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n796), .B1(new_n806), .B2(new_n204), .ZN(G1336gat));
  NOR2_X1   g606(.A1(new_n426), .A2(G92gat), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n803), .A2(new_n805), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(G92gat), .B1(new_n795), .B2(new_n426), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n727), .A2(new_n244), .A3(new_n687), .A4(new_n794), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n772), .B1(new_n799), .B2(new_n802), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n813), .A2(G92gat), .B1(new_n814), .B2(new_n808), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n812), .B1(new_n811), .B2(new_n815), .ZN(G1337gat));
  INV_X1    g615(.A(new_n794), .ZN(new_n817));
  INV_X1    g616(.A(new_n743), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n817), .B1(new_n818), .B2(new_n725), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n819), .A2(KEYINPUT116), .A3(new_n244), .A4(new_n706), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n821), .B1(new_n795), .B2(new_n705), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n822), .A3(G99gat), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n552), .A2(G99gat), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n803), .A2(new_n805), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(G1338gat));
  NOR2_X1   g625(.A1(new_n517), .A2(G106gat), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n803), .A2(new_n805), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(G106gat), .B1(new_n795), .B2(new_n517), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n727), .A2(new_n244), .A3(new_n712), .A4(new_n794), .ZN(new_n832));
  AOI22_X1  g631(.A1(new_n832), .A2(G106gat), .B1(new_n814), .B2(new_n827), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n831), .B1(new_n830), .B2(new_n833), .ZN(G1339gat));
  INV_X1    g633(.A(new_n241), .ZN(new_n835));
  INV_X1    g634(.A(new_n233), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n242), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n235), .A2(new_n238), .A3(new_n226), .ZN(new_n839));
  INV_X1    g638(.A(new_n202), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(KEYINPUT54), .A3(new_n239), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT55), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n838), .A2(new_n842), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n835), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n663), .A2(new_n665), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n659), .B1(new_n657), .B2(new_n658), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n673), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n677), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n717), .A2(new_n847), .A3(new_n851), .ZN(new_n852));
  AOI22_X1  g651(.A1(new_n678), .A2(new_n847), .B1(new_n851), .B2(new_n244), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n717), .ZN(new_n854));
  INV_X1    g653(.A(new_n603), .ZN(new_n855));
  AOI22_X1  g654(.A1(new_n854), .A2(new_n855), .B1(new_n767), .B2(new_n772), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n769), .A2(new_n856), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n757), .A2(new_n563), .A3(new_n687), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n278), .A3(new_n678), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n712), .A2(new_n566), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(G113gat), .B1(new_n862), .B2(new_n679), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n860), .A2(new_n863), .ZN(G1340gat));
  NAND3_X1  g663(.A1(new_n859), .A2(new_n280), .A3(new_n244), .ZN(new_n865));
  OAI21_X1  g664(.A(G120gat), .B1(new_n862), .B2(new_n772), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n866), .A2(KEYINPUT117), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n866), .A2(KEYINPUT117), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n865), .B1(new_n867), .B2(new_n868), .ZN(G1341gat));
  INV_X1    g668(.A(new_n862), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(G127gat), .A3(new_n603), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(KEYINPUT118), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(KEYINPUT118), .ZN(new_n873));
  AOI21_X1  g672(.A(G127gat), .B1(new_n859), .B2(new_n603), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(G1342gat));
  INV_X1    g674(.A(G134gat), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n859), .A2(new_n876), .A3(new_n717), .ZN(new_n877));
  OR3_X1    g676(.A1(new_n877), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n876), .B1(new_n870), .B2(new_n717), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n879), .B1(KEYINPUT56), .B2(new_n877), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT119), .B1(new_n877), .B2(KEYINPUT56), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n878), .A2(new_n880), .A3(new_n881), .ZN(G1343gat));
  NAND2_X1  g681(.A1(new_n767), .A2(new_n772), .ZN(new_n883));
  AND4_X1   g682(.A1(new_n653), .A2(new_n851), .A3(new_n847), .A4(new_n651), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n851), .A2(new_n244), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n886));
  INV_X1    g685(.A(new_n846), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n845), .B1(new_n838), .B2(new_n842), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n886), .B(new_n241), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n678), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n847), .A2(new_n886), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n885), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n884), .B1(new_n892), .B2(new_n654), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n883), .B1(new_n893), .B2(new_n603), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n894), .A2(KEYINPUT121), .A3(KEYINPUT57), .A4(new_n712), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n683), .A2(new_n426), .A3(new_n705), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n894), .A2(KEYINPUT57), .A3(new_n712), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n856), .A2(new_n517), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n899), .B(new_n900), .C1(KEYINPUT57), .C2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n898), .A2(new_n902), .A3(new_n678), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(G141gat), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT58), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n678), .A2(new_n247), .ZN(new_n906));
  XOR2_X1   g705(.A(new_n906), .B(KEYINPUT122), .Z(new_n907));
  INV_X1    g706(.A(new_n901), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n683), .A2(new_n705), .ZN(new_n909));
  OR3_X1    g708(.A1(new_n908), .A2(KEYINPUT123), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT123), .B1(new_n908), .B2(new_n909), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(new_n426), .A3(new_n911), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n904), .B(new_n905), .C1(new_n907), .C2(new_n912), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n908), .A2(new_n896), .A3(new_n907), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n914), .B1(new_n903), .B2(G141gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n913), .B1(new_n915), .B2(new_n905), .ZN(G1344gat));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT57), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n894), .A2(new_n918), .A3(new_n712), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT57), .B1(new_n856), .B2(new_n517), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n919), .A2(new_n920), .A3(new_n244), .A4(new_n897), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n917), .B1(new_n921), .B2(G148gat), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n922), .A2(KEYINPUT124), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n898), .A2(new_n902), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n917), .B(G148gat), .C1(new_n924), .C2(new_n772), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n922), .A2(KEYINPUT124), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  OR3_X1    g726(.A1(new_n912), .A2(G148gat), .A3(new_n772), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1345gat));
  NAND2_X1  g728(.A1(new_n269), .A2(new_n270), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n924), .A2(new_n930), .A3(new_n855), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n912), .A2(new_n855), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(new_n932), .B2(new_n930), .ZN(G1346gat));
  NOR3_X1   g732(.A1(new_n924), .A2(new_n257), .A3(new_n654), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n912), .A2(new_n654), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n935), .B2(new_n257), .ZN(G1347gat));
  NAND2_X1  g735(.A1(new_n854), .A2(new_n855), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n883), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(new_n769), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n757), .A2(new_n563), .A3(new_n426), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n943), .A2(new_n358), .A3(new_n678), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n940), .A2(new_n698), .A3(new_n687), .A4(new_n711), .ZN(new_n945));
  OAI21_X1  g744(.A(G169gat), .B1(new_n945), .B2(new_n679), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(G1348gat));
  AOI21_X1  g746(.A(G176gat), .B1(new_n943), .B2(new_n244), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n945), .A2(new_n230), .A3(new_n772), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(G1349gat));
  NAND3_X1  g749(.A1(new_n943), .A2(new_n348), .A3(new_n603), .ZN(new_n951));
  OAI21_X1  g750(.A(G183gat), .B1(new_n945), .B2(new_n855), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT60), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n954), .A2(KEYINPUT125), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n953), .B(new_n955), .ZN(G1350gat));
  OAI21_X1  g755(.A(G190gat), .B1(new_n945), .B2(new_n654), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT61), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n943), .A2(new_n349), .A3(new_n717), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1351gat));
  AND2_X1   g759(.A1(new_n919), .A2(new_n920), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n706), .A2(new_n683), .A3(new_n426), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(G197gat), .B1(new_n963), .B2(new_n679), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n757), .A2(new_n687), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n939), .A2(new_n706), .A3(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(G197gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n966), .A2(new_n967), .A3(new_n678), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n964), .A2(new_n968), .ZN(G1352gat));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n966), .A2(new_n232), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n971), .B1(new_n972), .B2(new_n244), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n966), .A2(new_n232), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n974), .A2(KEYINPUT126), .A3(new_n772), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n970), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n961), .A2(new_n244), .A3(new_n962), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(G204gat), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n972), .A2(new_n971), .A3(new_n244), .ZN(new_n979));
  OAI21_X1  g778(.A(KEYINPUT126), .B1(new_n974), .B2(new_n772), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n979), .A2(KEYINPUT62), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n976), .A2(new_n978), .A3(new_n981), .ZN(G1353gat));
  OAI21_X1  g781(.A(G211gat), .B1(new_n963), .B2(new_n855), .ZN(new_n983));
  NAND2_X1  g782(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n984));
  OR2_X1    g783(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n966), .A2(new_n596), .A3(new_n603), .ZN(new_n987));
  OAI211_X1 g786(.A(new_n986), .B(new_n987), .C1(new_n983), .C2(new_n985), .ZN(G1354gat));
  OAI21_X1  g787(.A(G218gat), .B1(new_n963), .B2(new_n654), .ZN(new_n989));
  INV_X1    g788(.A(G218gat), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n966), .A2(new_n990), .A3(new_n717), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n989), .A2(new_n991), .ZN(G1355gat));
endmodule


