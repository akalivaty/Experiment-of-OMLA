//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n557, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1170, new_n1171, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  OR2_X1    g032(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n458));
  NAND2_X1  g033(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n460), .A2(G137), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  OR3_X1    g037(.A1(new_n462), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT68), .ZN(new_n467));
  AND3_X1   g042(.A1(new_n463), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n462), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n461), .A2(new_n468), .B1(G101), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n464), .A2(new_n466), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT67), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n464), .A2(new_n466), .A3(new_n474), .A4(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n460), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n470), .A2(new_n479), .ZN(G160));
  OAI221_X1 g055(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n460), .C2(G112), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n468), .A2(new_n478), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G2105), .ZN(new_n485));
  AOI21_X1  g060(.A(KEYINPUT69), .B1(new_n468), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n463), .A2(new_n467), .A3(new_n464), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n488));
  NOR3_X1   g063(.A1(new_n487), .A2(new_n488), .A3(G2105), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n484), .B1(new_n491), .B2(G136), .ZN(G162));
  NAND3_X1  g067(.A1(new_n460), .A2(KEYINPUT4), .A3(G138), .ZN(new_n493));
  NAND2_X1  g068(.A1(G126), .A2(G2105), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n487), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n458), .A2(G138), .A3(new_n459), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(new_n471), .ZN(new_n497));
  AND2_X1   g072(.A1(G114), .A2(G2105), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(G102), .B2(new_n485), .ZN(new_n499));
  OAI22_X1  g074(.A1(new_n497), .A2(KEYINPUT4), .B1(new_n462), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n495), .A2(new_n500), .ZN(G164));
  NAND2_X1  g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  OR2_X1    g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT70), .B(KEYINPUT6), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT71), .B1(new_n510), .B2(new_n508), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n513), .A2(KEYINPUT70), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(KEYINPUT70), .ZN(new_n515));
  OAI211_X1 g090(.A(new_n512), .B(G651), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n517), .A2(G88), .A3(new_n506), .A4(new_n518), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n517), .A2(G50), .A3(G543), .A4(new_n518), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT72), .ZN(new_n521));
  AOI21_X1  g096(.A(KEYINPUT72), .B1(new_n519), .B2(new_n520), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n509), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT73), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n525));
  OAI211_X1 g100(.A(new_n525), .B(new_n509), .C1(new_n521), .C2(new_n522), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(G166));
  NAND2_X1  g102(.A1(new_n517), .A2(new_n518), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n505), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT74), .B(G89), .Z(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AND3_X1   g106(.A1(new_n517), .A2(G543), .A3(new_n518), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G51), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n506), .A2(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n531), .A2(new_n533), .A3(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n505), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n529), .A2(G90), .B1(G651), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n532), .A2(G52), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  XOR2_X1   g122(.A(KEYINPUT75), .B(G81), .Z(new_n548));
  NAND2_X1  g123(.A1(new_n529), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n532), .A2(G43), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n508), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT76), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(new_n532), .A2(G53), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n532), .A2(new_n564), .A3(G53), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(KEYINPUT77), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n508), .B1(new_n567), .B2(KEYINPUT77), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n529), .A2(G91), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G166), .ZN(G303));
  INV_X1    g147(.A(G74), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n508), .B1(new_n505), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n532), .B2(G49), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n529), .A2(G87), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(G288));
  AND2_X1   g152(.A1(new_n517), .A2(new_n518), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n578), .A2(G86), .A3(new_n506), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(KEYINPUT78), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n529), .A2(new_n581), .A3(G86), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n505), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n532), .A2(G48), .B1(G651), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n580), .A2(new_n582), .A3(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(G72), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G60), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n505), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n529), .A2(G85), .B1(G651), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n532), .A2(G47), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(new_n529), .A2(G92), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n529), .A2(KEYINPUT10), .A3(G92), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n505), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n532), .A2(G54), .B1(G651), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n603), .A2(new_n604), .B1(new_n605), .B2(KEYINPUT79), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(KEYINPUT79), .B2(new_n605), .ZN(G284));
  OAI21_X1  g182(.A(new_n606), .B1(KEYINPUT79), .B2(new_n605), .ZN(G321));
  NOR2_X1   g183(.A1(G286), .A2(new_n604), .ZN(new_n609));
  INV_X1    g184(.A(G299), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n604), .ZN(G297));
  XNOR2_X1  g186(.A(G297), .B(KEYINPUT80), .ZN(G280));
  AND2_X1   g187(.A1(new_n598), .A2(new_n602), .ZN(new_n613));
  XOR2_X1   g188(.A(KEYINPUT81), .B(G559), .Z(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(G860), .B2(new_n614), .ZN(G148));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n554), .A2(new_n604), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT11), .Z(G282));
  INV_X1    g196(.A(new_n620), .ZN(G323));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  INV_X1    g198(.A(G111), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n623), .B1(new_n478), .B2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(new_n482), .ZN(new_n626));
  AND2_X1   g201(.A1(new_n626), .A2(G123), .ZN(new_n627));
  AOI211_X1 g202(.A(new_n625), .B(new_n627), .C1(new_n491), .C2(G135), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(G2096), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(G2096), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n485), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT12), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT82), .B(G2100), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n630), .A2(new_n631), .A3(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XOR2_X1   g214(.A(G2443), .B(G2446), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G1341), .B(G1348), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT83), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2427), .B(G2430), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n646), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(KEYINPUT14), .A3(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n643), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n643), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(G401));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2072), .B(G2078), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT18), .Z(new_n660));
  INV_X1    g235(.A(new_n656), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n657), .A2(KEYINPUT17), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(new_n658), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n661), .B2(new_n662), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n656), .A2(new_n658), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n657), .B1(new_n666), .B2(KEYINPUT17), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n660), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT84), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2096), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2100), .ZN(G227));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n674), .A2(new_n675), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n673), .A2(new_n678), .A3(new_n676), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n673), .A2(new_n678), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n681));
  AOI211_X1 g256(.A(new_n677), .B(new_n679), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(new_n680), .B2(new_n681), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n685), .B(new_n688), .ZN(G229));
  NAND3_X1  g264(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT94), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT25), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n491), .A2(G139), .ZN(new_n693));
  NAND2_X1  g268(.A1(G115), .A2(G2104), .ZN(new_n694));
  INV_X1    g269(.A(G127), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n694), .B1(new_n471), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(new_n478), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT95), .Z(new_n698));
  NAND3_X1  g273(.A1(new_n692), .A2(new_n693), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT96), .ZN(new_n700));
  MUX2_X1   g275(.A(G33), .B(new_n700), .S(G29), .Z(new_n701));
  NOR2_X1   g276(.A1(new_n701), .A2(G2072), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT97), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT101), .B(KEYINPUT23), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT102), .ZN(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G20), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n705), .B(new_n707), .Z(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G299), .B2(G16), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1956), .ZN(new_n710));
  INV_X1    g285(.A(G2090), .ZN(new_n711));
  NOR2_X1   g286(.A1(G29), .A2(G35), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G162), .B2(G29), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n710), .B1(new_n711), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT103), .ZN(new_n717));
  NOR2_X1   g292(.A1(G171), .A2(new_n706), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G5), .B2(new_n706), .ZN(new_n719));
  INV_X1    g294(.A(G1961), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT99), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n719), .A2(new_n720), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G26), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT28), .ZN(new_n726));
  OAI221_X1 g301(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n460), .C2(G116), .ZN(new_n727));
  INV_X1    g302(.A(G128), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n482), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n491), .B2(G140), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n726), .B1(new_n730), .B2(new_n724), .ZN(new_n731));
  INV_X1    g306(.A(G2067), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n706), .A2(G21), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G168), .B2(new_n706), .ZN(new_n735));
  INV_X1    g310(.A(G1966), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n723), .A2(new_n733), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n724), .A2(G32), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n491), .A2(G141), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n469), .A2(G105), .ZN(new_n741));
  NAND3_X1  g316(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT26), .Z(new_n743));
  INV_X1    g318(.A(G129), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n741), .B(new_n743), .C1(new_n482), .C2(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n739), .B1(new_n746), .B2(new_n724), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT27), .B(G1996), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n715), .A2(new_n711), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT31), .B(G11), .Z(new_n751));
  INV_X1    g326(.A(G28), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n752), .A2(KEYINPUT30), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT98), .ZN(new_n754));
  AOI21_X1  g329(.A(G29), .B1(new_n752), .B2(KEYINPUT30), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n751), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n629), .B2(new_n724), .ZN(new_n757));
  NOR2_X1   g332(.A1(G27), .A2(G29), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G164), .B2(G29), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G2078), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(G160), .A2(G29), .ZN(new_n762));
  AND2_X1   g337(.A1(KEYINPUT24), .A2(G34), .ZN(new_n763));
  NOR2_X1   g338(.A1(KEYINPUT24), .A2(G34), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n724), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G2084), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n749), .A2(new_n750), .A3(new_n761), .A4(new_n767), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n722), .A2(new_n738), .A3(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G4), .A2(G16), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT92), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n603), .B2(new_n706), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT93), .B(G1348), .Z(new_n773));
  AND2_X1   g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G16), .A2(G19), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n554), .B2(G16), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(G1341), .Z(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n772), .B2(new_n773), .ZN(new_n778));
  AOI211_X1 g353(.A(new_n774), .B(new_n778), .C1(G2072), .C2(new_n701), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n703), .A2(new_n717), .A3(new_n769), .A4(new_n779), .ZN(new_n780));
  MUX2_X1   g355(.A(G23), .B(G288), .S(G16), .Z(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT33), .B(G1976), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n781), .B(new_n782), .Z(new_n783));
  AND3_X1   g358(.A1(new_n580), .A2(new_n582), .A3(new_n586), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(G16), .ZN(new_n785));
  OR2_X1    g360(.A1(G6), .A2(G16), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT88), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n785), .A2(KEYINPUT88), .A3(new_n786), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT32), .B(G1981), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n792), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n789), .A2(new_n790), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n783), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n706), .A2(G22), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G166), .B2(new_n706), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT89), .B(G1971), .Z(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n798), .A2(new_n800), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n796), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(KEYINPUT34), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT34), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n796), .B(new_n805), .C1(new_n801), .C2(new_n802), .ZN(new_n806));
  NOR2_X1   g381(.A1(G25), .A2(G29), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n626), .A2(G119), .ZN(new_n808));
  OAI221_X1 g383(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n460), .C2(G107), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT86), .ZN(new_n810));
  AOI211_X1 g385(.A(new_n808), .B(new_n810), .C1(new_n491), .C2(G131), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n807), .B1(new_n811), .B2(G29), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT35), .B(G1991), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT87), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n812), .B(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(G16), .A2(G24), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G290), .B2(new_n706), .ZN(new_n817));
  INV_X1    g392(.A(G1986), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n815), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AND3_X1   g396(.A1(new_n806), .A2(KEYINPUT90), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(KEYINPUT90), .B1(new_n806), .B2(new_n821), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n804), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT91), .B(KEYINPUT36), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n825), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n804), .B(new_n827), .C1(new_n822), .C2(new_n823), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n780), .B1(new_n826), .B2(new_n828), .ZN(G311));
  NAND2_X1  g404(.A1(new_n826), .A2(new_n828), .ZN(new_n830));
  INV_X1    g405(.A(new_n780), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(G150));
  NAND2_X1  g407(.A1(new_n613), .A2(G559), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT38), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n529), .A2(G93), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n532), .A2(G55), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(new_n508), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n835), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT104), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n835), .A2(KEYINPUT104), .A3(new_n836), .A4(new_n838), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n841), .A2(new_n553), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n554), .A2(new_n839), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n834), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n847));
  AOI21_X1  g422(.A(G860), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n847), .B2(new_n846), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n841), .A2(new_n842), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G860), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT37), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n852), .ZN(G145));
  INV_X1    g428(.A(KEYINPUT106), .ZN(new_n854));
  INV_X1    g429(.A(G164), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n730), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n746), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n856), .A2(new_n857), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n699), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n700), .B2(new_n860), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n811), .A2(new_n633), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n810), .A2(new_n808), .ZN(new_n864));
  INV_X1    g439(.A(G131), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n864), .B1(new_n865), .B2(new_n490), .ZN(new_n866));
  INV_X1    g441(.A(new_n633), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n626), .A2(G130), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT105), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n491), .A2(G142), .ZN(new_n872));
  OAI221_X1 g447(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n460), .C2(G118), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n869), .B(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n862), .A2(new_n875), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n869), .B(new_n874), .Z(new_n877));
  OAI211_X1 g452(.A(new_n877), .B(new_n861), .C1(new_n700), .C2(new_n860), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(G162), .B(G160), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n629), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n854), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n881), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n876), .A2(new_n878), .A3(KEYINPUT106), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(G37), .B1(new_n879), .B2(new_n881), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g463(.A(KEYINPUT111), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n613), .A2(new_n610), .ZN(new_n890));
  AOI22_X1  g465(.A1(new_n598), .A2(new_n602), .B1(new_n566), .B2(new_n570), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT107), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n890), .A2(KEYINPUT107), .A3(new_n892), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n617), .A2(new_n845), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n616), .B1(new_n844), .B2(new_n843), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n895), .B(new_n896), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n616), .B(new_n845), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n890), .A2(new_n892), .A3(KEYINPUT41), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT41), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n603), .A2(G299), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n902), .B1(new_n903), .B2(new_n891), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n899), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT109), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n524), .A2(new_n784), .A3(new_n526), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n784), .B1(new_n524), .B2(new_n526), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(G290), .A2(G288), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n591), .A2(new_n575), .A3(new_n576), .A4(new_n592), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n519), .A2(new_n520), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT72), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT72), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n525), .B1(new_n920), .B2(new_n509), .ZN(new_n921));
  INV_X1    g496(.A(new_n526), .ZN(new_n922));
  OAI21_X1  g497(.A(G305), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n524), .A2(new_n784), .A3(new_n526), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n914), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT108), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n928));
  AOI211_X1 g503(.A(new_n928), .B(new_n914), .C1(new_n923), .C2(new_n924), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n908), .B(new_n915), .C1(new_n927), .C2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n926), .B1(new_n909), .B2(new_n910), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n928), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n925), .A2(KEYINPUT108), .A3(new_n926), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n936), .A2(new_n908), .A3(KEYINPUT42), .A4(new_n915), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n907), .B1(new_n932), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n932), .A2(new_n937), .A3(new_n907), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n932), .A2(new_n937), .A3(new_n907), .A4(KEYINPUT110), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n604), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n850), .A2(new_n604), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n889), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n940), .A2(new_n939), .ZN(new_n947));
  INV_X1    g522(.A(new_n938), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n947), .A2(new_n948), .A3(new_n942), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(G868), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(KEYINPUT111), .A3(new_n944), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n946), .A2(new_n951), .ZN(G295));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n944), .ZN(G331));
  AND2_X1   g528(.A1(G301), .A2(G286), .ZN(new_n954));
  NOR2_X1   g529(.A1(G301), .A2(G286), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n845), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n843), .B(new_n844), .C1(new_n954), .C2(new_n955), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(new_n893), .ZN(new_n960));
  INV_X1    g535(.A(new_n905), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n960), .B1(new_n961), .B2(new_n959), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n936), .A2(new_n915), .ZN(new_n963));
  AOI21_X1  g538(.A(G37), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n936), .A2(new_n915), .ZN(new_n965));
  INV_X1    g540(.A(new_n959), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n966), .A2(new_n905), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n965), .B1(new_n967), .B2(new_n960), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n964), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT44), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n961), .A2(new_n972), .A3(new_n959), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT112), .B1(new_n966), .B2(new_n905), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n895), .A2(new_n896), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n966), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n973), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n965), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n969), .B1(new_n978), .B2(new_n964), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT113), .B1(new_n971), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n977), .A2(new_n965), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n962), .A2(new_n963), .ZN(new_n982));
  INV_X1    g557(.A(G37), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT43), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n985), .A2(new_n986), .A3(KEYINPUT44), .A4(new_n970), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n980), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n969), .B1(new_n981), .B2(new_n984), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n964), .A2(new_n968), .A3(KEYINPUT43), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n988), .A2(new_n992), .ZN(G397));
  AND3_X1   g568(.A1(new_n470), .A2(new_n479), .A3(G40), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n995));
  INV_X1    g570(.A(G1384), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(new_n495), .B2(new_n500), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n994), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n998), .A2(KEYINPUT114), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(KEYINPUT114), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1002), .A2(G1996), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n1003), .B(KEYINPUT46), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n730), .B(G2067), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1002), .B1(new_n746), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n730), .A2(new_n732), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n746), .B(G1996), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n1005), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n811), .A2(new_n813), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1010), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n1001), .ZN(new_n1015));
  NOR2_X1   g590(.A1(G290), .A2(G1986), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1001), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT48), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n811), .B(new_n813), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1012), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1018), .B1(new_n1020), .B2(new_n1002), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n1009), .A2(new_n1015), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G8), .ZN(new_n1023));
  INV_X1    g598(.A(new_n997), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1023), .B1(new_n994), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1976), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n575), .A2(new_n576), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n586), .A2(new_n579), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(G1981), .ZN(new_n1029));
  INV_X1    g604(.A(G1981), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n580), .A2(new_n1030), .A3(new_n582), .A4(new_n586), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n1031), .A3(KEYINPUT49), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1032), .B(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT49), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1025), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1027), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1031), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1025), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(G288), .B2(new_n1026), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n575), .A2(new_n576), .A3(KEYINPUT116), .A4(G1976), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1042), .A2(new_n1025), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT52), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT52), .B1(G288), .B2(new_n1026), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1042), .A2(new_n1046), .A3(new_n1025), .A4(new_n1043), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1048), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1049));
  NAND3_X1  g624(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1051), .B1(G166), .B2(new_n1023), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n997), .A2(new_n995), .ZN(new_n1054));
  OAI211_X1 g629(.A(KEYINPUT45), .B(new_n996), .C1(new_n495), .C2(new_n500), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(new_n994), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1057), .A2(G1971), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1060), .B(new_n996), .C1(new_n495), .C2(new_n500), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1059), .A2(new_n994), .A3(new_n1061), .ZN(new_n1062));
  OR2_X1    g637(.A1(new_n1062), .A2(G2090), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1023), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1049), .A2(new_n1053), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1040), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1053), .A2(new_n1064), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1059), .A2(new_n994), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1059), .A2(new_n994), .A3(KEYINPUT118), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1061), .A3(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1058), .B1(new_n1072), .B2(G2090), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G8), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1074), .A2(new_n1052), .A3(new_n1050), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1056), .A2(new_n736), .ZN(new_n1076));
  INV_X1    g651(.A(G2084), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1059), .A2(new_n994), .A3(new_n1077), .A4(new_n1061), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1023), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(G168), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT119), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1079), .A2(new_n1082), .A3(G168), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1067), .A2(new_n1049), .A3(new_n1075), .A4(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT63), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1053), .A2(new_n1064), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1086), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1088), .A2(new_n1067), .A3(new_n1049), .A4(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1066), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G2078), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1054), .A2(new_n994), .A3(new_n1092), .A4(new_n1055), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1093), .A2(new_n1094), .B1(new_n1062), .B2(new_n720), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n470), .A2(new_n479), .A3(G40), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1096), .B1(new_n995), .B2(new_n997), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1097), .A2(KEYINPUT53), .A3(new_n1092), .A4(new_n1055), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1095), .A2(G301), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(G301), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT54), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G171), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1095), .A2(G301), .A3(new_n1098), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1107));
  AND4_X1   g682(.A1(new_n1075), .A2(new_n1107), .A3(new_n1067), .A4(new_n1049), .ZN(new_n1108));
  INV_X1    g683(.A(G1956), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT56), .B(G2072), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1110), .B(KEYINPUT121), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1072), .A2(new_n1109), .B1(new_n1057), .B2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1113), .B1(new_n566), .B2(new_n570), .ZN(new_n1114));
  NOR2_X1   g689(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1114), .B1(new_n610), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n994), .A2(new_n1024), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1119), .A2(G2067), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1120), .B1(new_n773), .B2(new_n1062), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(new_n603), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1117), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT58), .B(G1341), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1124), .B(KEYINPUT122), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1119), .A2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(G1996), .B2(new_n1056), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n554), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT59), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1127), .A2(new_n1130), .A3(new_n554), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT60), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1121), .A2(new_n1133), .A3(new_n613), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1121), .B(new_n613), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1132), .B(new_n1134), .C1(new_n1135), .C2(new_n1133), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1112), .A2(KEYINPUT61), .A3(new_n1116), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT61), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1123), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(G168), .A2(new_n1023), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT51), .B1(new_n1079), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g719(.A(KEYINPUT123), .B(KEYINPUT51), .C1(new_n1079), .C2(new_n1141), .ZN(new_n1145));
  OR3_X1    g720(.A1(new_n1079), .A2(KEYINPUT51), .A3(new_n1141), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1079), .A2(G286), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT124), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1147), .A2(KEYINPUT124), .A3(new_n1148), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1108), .B(new_n1140), .C1(new_n1149), .C2(new_n1151), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1091), .A2(new_n1152), .A3(KEYINPUT125), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT125), .B1(new_n1091), .B2(new_n1152), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT62), .B1(new_n1151), .B2(new_n1149), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1149), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(new_n1157), .A3(new_n1150), .ZN(new_n1158));
  AND4_X1   g733(.A1(new_n1075), .A2(new_n1067), .A3(new_n1049), .A4(new_n1100), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1155), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1153), .A2(new_n1154), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1016), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT115), .ZN(new_n1163));
  NAND2_X1  g738(.A1(G290), .A2(G1986), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1162), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1165), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1002), .B1(new_n1020), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1022), .B1(new_n1161), .B2(new_n1167), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g743(.A1(new_n654), .A2(G319), .ZN(new_n1170));
  NOR3_X1   g744(.A1(G229), .A2(G227), .A3(new_n1170), .ZN(new_n1171));
  XOR2_X1   g745(.A(new_n1171), .B(KEYINPUT127), .Z(new_n1172));
  NAND4_X1  g746(.A1(new_n887), .A2(new_n989), .A3(new_n991), .A4(new_n1172), .ZN(G225));
  INV_X1    g747(.A(G225), .ZN(G308));
endmodule


