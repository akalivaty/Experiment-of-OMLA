

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596;

  INV_X1 U326 ( .A(KEYINPUT100), .ZN(n413) );
  XNOR2_X1 U327 ( .A(n318), .B(n317), .ZN(n326) );
  XNOR2_X1 U328 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U329 ( .A(n402), .B(n358), .ZN(n359) );
  NOR2_X1 U330 ( .A1(n420), .A2(n419), .ZN(n509) );
  XNOR2_X1 U331 ( .A(n414), .B(n413), .ZN(n420) );
  XNOR2_X1 U332 ( .A(n482), .B(KEYINPUT48), .ZN(n483) );
  XOR2_X1 U333 ( .A(n335), .B(n334), .Z(n555) );
  XNOR2_X1 U334 ( .A(n367), .B(n366), .ZN(n294) );
  INV_X1 U335 ( .A(KEYINPUT23), .ZN(n356) );
  XNOR2_X1 U336 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U337 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U338 ( .A(n427), .B(n426), .ZN(n429) );
  INV_X1 U339 ( .A(n434), .ZN(n435) );
  XNOR2_X1 U340 ( .A(n466), .B(KEYINPUT64), .ZN(n467) );
  NOR2_X1 U341 ( .A1(n490), .A2(n422), .ZN(n423) );
  XNOR2_X1 U342 ( .A(n440), .B(n294), .ZN(n368) );
  XNOR2_X1 U343 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U344 ( .A(n590), .B(n467), .ZN(n494) );
  XNOR2_X1 U345 ( .A(n369), .B(n368), .ZN(n373) );
  XNOR2_X1 U346 ( .A(n438), .B(n437), .ZN(n442) );
  XNOR2_X1 U347 ( .A(n387), .B(KEYINPUT26), .ZN(n561) );
  INV_X1 U348 ( .A(G218GAT), .ZN(n491) );
  INV_X1 U349 ( .A(G106GAT), .ZN(n500) );
  XNOR2_X1 U350 ( .A(n491), .B(KEYINPUT62), .ZN(n492) );
  XNOR2_X1 U351 ( .A(n504), .B(G197GAT), .ZN(n505) );
  XNOR2_X1 U352 ( .A(n500), .B(KEYINPUT44), .ZN(n501) );
  XNOR2_X1 U353 ( .A(n497), .B(KEYINPUT114), .ZN(n498) );
  XNOR2_X1 U354 ( .A(n460), .B(G43GAT), .ZN(n461) );
  XNOR2_X1 U355 ( .A(n493), .B(n492), .ZN(G1355GAT) );
  XNOR2_X1 U356 ( .A(n506), .B(n505), .ZN(G1352GAT) );
  XNOR2_X1 U357 ( .A(n499), .B(n498), .ZN(G1338GAT) );
  XOR2_X1 U358 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n296) );
  XNOR2_X1 U359 ( .A(KEYINPUT20), .B(KEYINPUT86), .ZN(n295) );
  XNOR2_X1 U360 ( .A(n296), .B(n295), .ZN(n314) );
  XNOR2_X1 U361 ( .A(G183GAT), .B(KEYINPUT19), .ZN(n297) );
  XNOR2_X1 U362 ( .A(n297), .B(KEYINPUT17), .ZN(n298) );
  XOR2_X1 U363 ( .A(n298), .B(KEYINPUT18), .Z(n300) );
  XNOR2_X1 U364 ( .A(G169GAT), .B(G190GAT), .ZN(n299) );
  XOR2_X1 U365 ( .A(n300), .B(n299), .Z(n383) );
  XOR2_X1 U366 ( .A(G71GAT), .B(G120GAT), .Z(n302) );
  XNOR2_X1 U367 ( .A(G99GAT), .B(G176GAT), .ZN(n301) );
  XNOR2_X1 U368 ( .A(n302), .B(n301), .ZN(n427) );
  XOR2_X1 U369 ( .A(n383), .B(n427), .Z(n312) );
  XOR2_X1 U370 ( .A(G43GAT), .B(G134GAT), .Z(n316) );
  XOR2_X1 U371 ( .A(KEYINPUT65), .B(KEYINPUT83), .Z(n304) );
  XNOR2_X1 U372 ( .A(G15GAT), .B(KEYINPUT87), .ZN(n303) );
  XNOR2_X1 U373 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U374 ( .A(n316), .B(n305), .Z(n307) );
  NAND2_X1 U375 ( .A1(G227GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U376 ( .A(n307), .B(n306), .ZN(n310) );
  XOR2_X1 U377 ( .A(G127GAT), .B(KEYINPUT82), .Z(n309) );
  XNOR2_X1 U378 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n308) );
  XNOR2_X1 U379 ( .A(n309), .B(n308), .ZN(n391) );
  XOR2_X1 U380 ( .A(n310), .B(n391), .Z(n311) );
  XNOR2_X1 U381 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X2 U382 ( .A(n314), .B(n313), .ZN(n574) );
  XOR2_X1 U383 ( .A(G50GAT), .B(G162GAT), .Z(n366) );
  XOR2_X1 U384 ( .A(G85GAT), .B(KEYINPUT73), .Z(n439) );
  XNOR2_X1 U385 ( .A(n366), .B(n439), .ZN(n318) );
  AND2_X1 U386 ( .A1(G232GAT), .A2(G233GAT), .ZN(n315) );
  XOR2_X1 U387 ( .A(KEYINPUT76), .B(KEYINPUT9), .Z(n320) );
  XNOR2_X1 U388 ( .A(G218GAT), .B(KEYINPUT75), .ZN(n319) );
  XNOR2_X1 U389 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U390 ( .A(KEYINPUT11), .B(G92GAT), .Z(n322) );
  XNOR2_X1 U391 ( .A(G99GAT), .B(KEYINPUT74), .ZN(n321) );
  XNOR2_X1 U392 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U393 ( .A(n324), .B(n323), .Z(n325) );
  XNOR2_X1 U394 ( .A(n326), .B(n325), .ZN(n330) );
  XOR2_X1 U395 ( .A(KEYINPUT10), .B(KEYINPUT66), .Z(n328) );
  XNOR2_X1 U396 ( .A(G190GAT), .B(G106GAT), .ZN(n327) );
  XNOR2_X1 U397 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U398 ( .A(n330), .B(n329), .ZN(n335) );
  XOR2_X1 U399 ( .A(KEYINPUT7), .B(KEYINPUT68), .Z(n332) );
  XNOR2_X1 U400 ( .A(G36GAT), .B(G29GAT), .ZN(n331) );
  XNOR2_X1 U401 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U402 ( .A(KEYINPUT8), .B(n333), .ZN(n453) );
  INV_X1 U403 ( .A(n453), .ZN(n334) );
  XNOR2_X1 U404 ( .A(KEYINPUT36), .B(n555), .ZN(n490) );
  XOR2_X1 U405 ( .A(G57GAT), .B(KEYINPUT13), .Z(n434) );
  XNOR2_X1 U406 ( .A(G15GAT), .B(G1GAT), .ZN(n336) );
  XNOR2_X1 U407 ( .A(n336), .B(G8GAT), .ZN(n446) );
  XOR2_X1 U408 ( .A(n434), .B(n446), .Z(n338) );
  NAND2_X1 U409 ( .A1(G231GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U410 ( .A(n338), .B(n337), .ZN(n354) );
  XOR2_X1 U411 ( .A(KEYINPUT12), .B(KEYINPUT78), .Z(n340) );
  XNOR2_X1 U412 ( .A(KEYINPUT15), .B(KEYINPUT77), .ZN(n339) );
  XNOR2_X1 U413 ( .A(n340), .B(n339), .ZN(n352) );
  XOR2_X1 U414 ( .A(G78GAT), .B(G127GAT), .Z(n342) );
  XNOR2_X1 U415 ( .A(G183GAT), .B(G71GAT), .ZN(n341) );
  XNOR2_X1 U416 ( .A(n342), .B(n341), .ZN(n350) );
  XOR2_X1 U417 ( .A(KEYINPUT14), .B(KEYINPUT79), .Z(n344) );
  XNOR2_X1 U418 ( .A(KEYINPUT81), .B(KEYINPUT80), .ZN(n343) );
  XNOR2_X1 U419 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U420 ( .A(G64GAT), .B(G155GAT), .Z(n346) );
  XNOR2_X1 U421 ( .A(G22GAT), .B(G211GAT), .ZN(n345) );
  XNOR2_X1 U422 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U423 ( .A(n348), .B(n347), .Z(n349) );
  XNOR2_X1 U424 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U425 ( .A(n352), .B(n351), .Z(n353) );
  XOR2_X1 U426 ( .A(n354), .B(n353), .Z(n550) );
  INV_X1 U427 ( .A(n550), .ZN(n594) );
  XOR2_X1 U428 ( .A(G141GAT), .B(G22GAT), .Z(n445) );
  XNOR2_X1 U429 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n355) );
  XNOR2_X1 U430 ( .A(n355), .B(KEYINPUT2), .ZN(n402) );
  NAND2_X1 U431 ( .A1(G228GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U432 ( .A(n445), .B(n359), .ZN(n369) );
  XNOR2_X1 U433 ( .A(G148GAT), .B(KEYINPUT72), .ZN(n360) );
  XNOR2_X1 U434 ( .A(n360), .B(KEYINPUT71), .ZN(n361) );
  XOR2_X1 U435 ( .A(n361), .B(G204GAT), .Z(n363) );
  XNOR2_X1 U436 ( .A(G78GAT), .B(G106GAT), .ZN(n362) );
  XNOR2_X1 U437 ( .A(n363), .B(n362), .ZN(n440) );
  XOR2_X1 U438 ( .A(KEYINPUT90), .B(KEYINPUT24), .Z(n365) );
  XNOR2_X1 U439 ( .A(KEYINPUT89), .B(KEYINPUT22), .ZN(n364) );
  XNOR2_X1 U440 ( .A(n365), .B(n364), .ZN(n367) );
  XOR2_X1 U441 ( .A(KEYINPUT91), .B(G218GAT), .Z(n371) );
  XNOR2_X1 U442 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n370) );
  XNOR2_X1 U443 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U444 ( .A(G197GAT), .B(n372), .Z(n380) );
  XNOR2_X1 U445 ( .A(n373), .B(n380), .ZN(n571) );
  XOR2_X1 U446 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n375) );
  NAND2_X1 U447 ( .A1(G226GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U448 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U449 ( .A(G204GAT), .B(G176GAT), .Z(n377) );
  XNOR2_X1 U450 ( .A(G36GAT), .B(G8GAT), .ZN(n376) );
  XNOR2_X1 U451 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U452 ( .A(n379), .B(n378), .Z(n382) );
  XOR2_X1 U453 ( .A(G92GAT), .B(G64GAT), .Z(n433) );
  XNOR2_X1 U454 ( .A(n380), .B(n433), .ZN(n381) );
  XNOR2_X1 U455 ( .A(n382), .B(n381), .ZN(n384) );
  XOR2_X1 U456 ( .A(n384), .B(n383), .Z(n539) );
  NOR2_X1 U457 ( .A1(n574), .A2(n539), .ZN(n385) );
  NOR2_X1 U458 ( .A1(n571), .A2(n385), .ZN(n386) );
  XOR2_X1 U459 ( .A(KEYINPUT25), .B(n386), .Z(n389) );
  NAND2_X1 U460 ( .A1(n571), .A2(n574), .ZN(n387) );
  XNOR2_X1 U461 ( .A(n539), .B(KEYINPUT27), .ZN(n415) );
  NOR2_X1 U462 ( .A1(n561), .A2(n415), .ZN(n388) );
  NOR2_X1 U463 ( .A1(n389), .A2(n388), .ZN(n390) );
  XNOR2_X1 U464 ( .A(n390), .B(KEYINPUT99), .ZN(n412) );
  XOR2_X1 U465 ( .A(n391), .B(G1GAT), .Z(n393) );
  NAND2_X1 U466 ( .A1(G225GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U467 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U468 ( .A(KEYINPUT92), .B(G57GAT), .Z(n395) );
  XNOR2_X1 U469 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n394) );
  XNOR2_X1 U470 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U471 ( .A(n397), .B(n396), .ZN(n401) );
  XOR2_X1 U472 ( .A(KEYINPUT93), .B(G148GAT), .Z(n399) );
  XNOR2_X1 U473 ( .A(G141GAT), .B(G120GAT), .ZN(n398) );
  XNOR2_X1 U474 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U475 ( .A(n401), .B(n400), .ZN(n406) );
  XOR2_X1 U476 ( .A(G85GAT), .B(G162GAT), .Z(n404) );
  XNOR2_X1 U477 ( .A(G29GAT), .B(n402), .ZN(n403) );
  XNOR2_X1 U478 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U479 ( .A(n406), .B(n405), .Z(n411) );
  XOR2_X1 U480 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n408) );
  XNOR2_X1 U481 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n407) );
  XNOR2_X1 U482 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U483 ( .A(G134GAT), .B(n409), .ZN(n410) );
  XNOR2_X1 U484 ( .A(n411), .B(n410), .ZN(n537) );
  NAND2_X1 U485 ( .A1(n412), .A2(n537), .ZN(n414) );
  NOR2_X1 U486 ( .A1(n415), .A2(n537), .ZN(n416) );
  XNOR2_X1 U487 ( .A(n416), .B(KEYINPUT98), .ZN(n559) );
  XNOR2_X1 U488 ( .A(KEYINPUT28), .B(KEYINPUT67), .ZN(n417) );
  XNOR2_X1 U489 ( .A(n417), .B(n571), .ZN(n534) );
  NAND2_X1 U490 ( .A1(n559), .A2(n534), .ZN(n543) );
  XOR2_X1 U491 ( .A(KEYINPUT88), .B(n574), .Z(n418) );
  NOR2_X1 U492 ( .A1(n543), .A2(n418), .ZN(n419) );
  NOR2_X1 U493 ( .A1(n594), .A2(n509), .ZN(n421) );
  XNOR2_X1 U494 ( .A(n421), .B(KEYINPUT103), .ZN(n422) );
  XOR2_X1 U495 ( .A(KEYINPUT37), .B(n423), .Z(n495) );
  NAND2_X1 U496 ( .A1(G230GAT), .A2(G233GAT), .ZN(n425) );
  INV_X1 U497 ( .A(KEYINPUT32), .ZN(n424) );
  INV_X1 U498 ( .A(KEYINPUT31), .ZN(n428) );
  NAND2_X1 U499 ( .A1(n429), .A2(n428), .ZN(n432) );
  INV_X1 U500 ( .A(n429), .ZN(n430) );
  NAND2_X1 U501 ( .A1(n430), .A2(KEYINPUT31), .ZN(n431) );
  NAND2_X1 U502 ( .A1(n432), .A2(n431), .ZN(n438) );
  XNOR2_X1 U503 ( .A(n433), .B(KEYINPUT33), .ZN(n436) );
  XNOR2_X1 U504 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U505 ( .A(n442), .B(n441), .ZN(n590) );
  XOR2_X1 U506 ( .A(KEYINPUT69), .B(G197GAT), .Z(n444) );
  XNOR2_X1 U507 ( .A(G169GAT), .B(G113GAT), .ZN(n443) );
  XNOR2_X1 U508 ( .A(n444), .B(n443), .ZN(n457) );
  XOR2_X1 U509 ( .A(n446), .B(n445), .Z(n448) );
  XNOR2_X1 U510 ( .A(G50GAT), .B(G43GAT), .ZN(n447) );
  XNOR2_X1 U511 ( .A(n448), .B(n447), .ZN(n452) );
  XOR2_X1 U512 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n450) );
  NAND2_X1 U513 ( .A1(G229GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U514 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U515 ( .A(n452), .B(n451), .Z(n455) );
  XOR2_X1 U516 ( .A(n453), .B(KEYINPUT29), .Z(n454) );
  XNOR2_X1 U517 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U518 ( .A(n457), .B(n456), .ZN(n546) );
  NOR2_X1 U519 ( .A1(n590), .A2(n546), .ZN(n510) );
  NAND2_X1 U520 ( .A1(n495), .A2(n510), .ZN(n459) );
  XNOR2_X1 U521 ( .A(KEYINPUT38), .B(KEYINPUT104), .ZN(n458) );
  XNOR2_X1 U522 ( .A(n459), .B(n458), .ZN(n522) );
  NOR2_X1 U523 ( .A1(n574), .A2(n522), .ZN(n462) );
  XNOR2_X1 U524 ( .A(KEYINPUT40), .B(KEYINPUT105), .ZN(n460) );
  XNOR2_X1 U525 ( .A(n462), .B(n461), .ZN(G1330GAT) );
  NOR2_X1 U526 ( .A1(n534), .A2(n522), .ZN(n465) );
  XNOR2_X1 U527 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n463) );
  XNOR2_X1 U528 ( .A(n463), .B(G50GAT), .ZN(n464) );
  XNOR2_X1 U529 ( .A(n465), .B(n464), .ZN(G1331GAT) );
  INV_X1 U530 ( .A(n539), .ZN(n485) );
  INV_X1 U531 ( .A(KEYINPUT41), .ZN(n466) );
  INV_X1 U532 ( .A(n546), .ZN(n575) );
  NAND2_X1 U533 ( .A1(n494), .A2(n575), .ZN(n468) );
  XOR2_X1 U534 ( .A(n468), .B(KEYINPUT46), .Z(n469) );
  NOR2_X1 U535 ( .A1(n594), .A2(n469), .ZN(n470) );
  NAND2_X1 U536 ( .A1(n470), .A2(n555), .ZN(n472) );
  XOR2_X1 U537 ( .A(KEYINPUT115), .B(KEYINPUT47), .Z(n471) );
  XNOR2_X1 U538 ( .A(n472), .B(n471), .ZN(n481) );
  INV_X1 U539 ( .A(KEYINPUT117), .ZN(n479) );
  NOR2_X1 U540 ( .A1(n490), .A2(n550), .ZN(n474) );
  INV_X1 U541 ( .A(KEYINPUT45), .ZN(n473) );
  XNOR2_X1 U542 ( .A(n474), .B(n473), .ZN(n475) );
  NOR2_X1 U543 ( .A1(n475), .A2(n590), .ZN(n476) );
  XOR2_X1 U544 ( .A(KEYINPUT116), .B(n476), .Z(n477) );
  NOR2_X1 U545 ( .A1(n575), .A2(n477), .ZN(n478) );
  XNOR2_X1 U546 ( .A(n479), .B(n478), .ZN(n480) );
  NOR2_X1 U547 ( .A1(n481), .A2(n480), .ZN(n484) );
  INV_X1 U548 ( .A(KEYINPUT118), .ZN(n482) );
  XNOR2_X1 U549 ( .A(n484), .B(n483), .ZN(n544) );
  NAND2_X1 U550 ( .A1(n485), .A2(n544), .ZN(n487) );
  XOR2_X1 U551 ( .A(KEYINPUT54), .B(KEYINPUT122), .Z(n486) );
  XNOR2_X1 U552 ( .A(n487), .B(n486), .ZN(n488) );
  NAND2_X1 U553 ( .A1(n537), .A2(n488), .ZN(n570) );
  NOR2_X1 U554 ( .A1(n561), .A2(n570), .ZN(n489) );
  XOR2_X1 U555 ( .A(KEYINPUT126), .B(n489), .Z(n503) );
  NOR2_X1 U556 ( .A1(n490), .A2(n503), .ZN(n493) );
  XOR2_X1 U557 ( .A(KEYINPUT108), .B(n494), .Z(n581) );
  NOR2_X1 U558 ( .A1(n575), .A2(n581), .ZN(n527) );
  NAND2_X1 U559 ( .A1(n527), .A2(n495), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n496), .B(KEYINPUT112), .ZN(n540) );
  NOR2_X1 U561 ( .A1(n540), .A2(n574), .ZN(n499) );
  INV_X1 U562 ( .A(G99GAT), .ZN(n497) );
  NOR2_X1 U563 ( .A1(n540), .A2(n534), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(G1339GAT) );
  INV_X1 U565 ( .A(n503), .ZN(n593) );
  NAND2_X1 U566 ( .A1(n575), .A2(n593), .ZN(n506) );
  XOR2_X1 U567 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n504) );
  INV_X1 U568 ( .A(n555), .ZN(n587) );
  NOR2_X1 U569 ( .A1(n587), .A2(n550), .ZN(n507) );
  XOR2_X1 U570 ( .A(KEYINPUT16), .B(n507), .Z(n508) );
  NOR2_X1 U571 ( .A1(n509), .A2(n508), .ZN(n526) );
  NAND2_X1 U572 ( .A1(n510), .A2(n526), .ZN(n518) );
  NOR2_X1 U573 ( .A1(n537), .A2(n518), .ZN(n512) );
  XNOR2_X1 U574 ( .A(KEYINPUT34), .B(KEYINPUT101), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U576 ( .A(G1GAT), .B(n513), .ZN(G1324GAT) );
  NOR2_X1 U577 ( .A1(n539), .A2(n518), .ZN(n514) );
  XOR2_X1 U578 ( .A(KEYINPUT102), .B(n514), .Z(n515) );
  XNOR2_X1 U579 ( .A(G8GAT), .B(n515), .ZN(G1325GAT) );
  NOR2_X1 U580 ( .A1(n574), .A2(n518), .ZN(n517) );
  XNOR2_X1 U581 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(G1326GAT) );
  NOR2_X1 U583 ( .A1(n534), .A2(n518), .ZN(n519) );
  XOR2_X1 U584 ( .A(G22GAT), .B(n519), .Z(G1327GAT) );
  NOR2_X1 U585 ( .A1(n537), .A2(n522), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(G1328GAT) );
  NOR2_X1 U588 ( .A1(n539), .A2(n522), .ZN(n523) );
  XOR2_X1 U589 ( .A(G36GAT), .B(n523), .Z(G1329GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n525) );
  XNOR2_X1 U591 ( .A(G57GAT), .B(KEYINPUT110), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(n530) );
  NAND2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U594 ( .A(KEYINPUT109), .B(n528), .Z(n533) );
  NOR2_X1 U595 ( .A1(n537), .A2(n533), .ZN(n529) );
  XOR2_X1 U596 ( .A(n530), .B(n529), .Z(G1332GAT) );
  NOR2_X1 U597 ( .A1(n539), .A2(n533), .ZN(n531) );
  XOR2_X1 U598 ( .A(G64GAT), .B(n531), .Z(G1333GAT) );
  NOR2_X1 U599 ( .A1(n574), .A2(n533), .ZN(n532) );
  XOR2_X1 U600 ( .A(G71GAT), .B(n532), .Z(G1334GAT) );
  NOR2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n536) );
  XNOR2_X1 U602 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(G1335GAT) );
  NOR2_X1 U604 ( .A1(n537), .A2(n540), .ZN(n538) );
  XOR2_X1 U605 ( .A(G85GAT), .B(n538), .Z(G1336GAT) );
  NOR2_X1 U606 ( .A1(n540), .A2(n539), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G92GAT), .B(KEYINPUT113), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(G1337GAT) );
  NOR2_X1 U609 ( .A1(n574), .A2(n543), .ZN(n545) );
  NAND2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n554) );
  NOR2_X1 U611 ( .A1(n546), .A2(n554), .ZN(n547) );
  XOR2_X1 U612 ( .A(G113GAT), .B(n547), .Z(G1340GAT) );
  NOR2_X1 U613 ( .A1(n581), .A2(n554), .ZN(n549) );
  XNOR2_X1 U614 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(G1341GAT) );
  NOR2_X1 U616 ( .A1(n550), .A2(n554), .ZN(n552) );
  XNOR2_X1 U617 ( .A(KEYINPUT119), .B(KEYINPUT50), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G127GAT), .B(n553), .ZN(G1342GAT) );
  NOR2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n557) );
  XNOR2_X1 U621 ( .A(KEYINPUT120), .B(KEYINPUT51), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(G134GAT), .B(n558), .ZN(G1343GAT) );
  NAND2_X1 U624 ( .A1(n544), .A2(n559), .ZN(n560) );
  NOR2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n568) );
  NAND2_X1 U626 ( .A1(n568), .A2(n575), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT52), .B(KEYINPUT121), .Z(n564) );
  NAND2_X1 U629 ( .A1(n568), .A2(n494), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n566) );
  XOR2_X1 U631 ( .A(G148GAT), .B(KEYINPUT53), .Z(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1345GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n594), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U635 ( .A1(n568), .A2(n587), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U637 ( .A(G169GAT), .B(KEYINPUT123), .Z(n577) );
  NOR2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n572), .B(KEYINPUT55), .ZN(n573) );
  NOR2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n586) );
  NAND2_X1 U641 ( .A1(n586), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1348GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n579) );
  XNOR2_X1 U644 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XOR2_X1 U646 ( .A(KEYINPUT124), .B(n580), .Z(n584) );
  INV_X1 U647 ( .A(n581), .ZN(n582) );
  NAND2_X1 U648 ( .A1(n582), .A2(n586), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1349GAT) );
  NAND2_X1 U650 ( .A1(n586), .A2(n594), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n585), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U652 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n589) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(G1351GAT) );
  XOR2_X1 U655 ( .A(G204GAT), .B(KEYINPUT61), .Z(n592) );
  NAND2_X1 U656 ( .A1(n590), .A2(n593), .ZN(n591) );
  XNOR2_X1 U657 ( .A(n592), .B(n591), .ZN(G1353GAT) );
  XOR2_X1 U658 ( .A(G211GAT), .B(KEYINPUT127), .Z(n596) );
  NAND2_X1 U659 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U660 ( .A(n596), .B(n595), .ZN(G1354GAT) );
endmodule

