//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT66), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  AND2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND3_X1   g034(.A1(new_n459), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n460));
  AOI21_X1  g035(.A(KEYINPUT67), .B1(new_n459), .B2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(G101), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n459), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g041(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n459), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(G160));
  OR2_X1    g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n459), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  OR2_X1    g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(new_n459), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n477), .B1(G136), .B2(new_n480), .ZN(G162));
  OAI211_X1 g056(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n482));
  OR2_X1    g057(.A1(G102), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n483), .A2(new_n485), .A3(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n463), .B2(new_n464), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n489), .B(new_n492), .C1(new_n464), .C2(new_n463), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n487), .B1(new_n491), .B2(new_n493), .ZN(G164));
  OR2_X1    g069(.A1(KEYINPUT5), .A2(G543), .ZN(new_n495));
  NAND2_X1  g070(.A1(KEYINPUT5), .A2(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n497), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n498));
  INV_X1    g073(.A(G651), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g075(.A(KEYINPUT6), .B(G651), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G50), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  OAI22_X1  g082(.A1(new_n504), .A2(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n502), .A2(new_n503), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n500), .A2(new_n510), .ZN(G166));
  NAND3_X1  g086(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n512), .B(KEYINPUT7), .ZN(new_n513));
  INV_X1    g088(.A(G89), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n513), .B1(new_n514), .B2(new_n508), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT68), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n497), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n505), .A2(new_n504), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT68), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n521));
  INV_X1    g096(.A(new_n502), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G51), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT69), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT69), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n521), .A2(new_n526), .A3(new_n523), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n515), .B1(new_n525), .B2(new_n527), .ZN(G168));
  NAND2_X1  g103(.A1(G77), .A2(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n517), .A2(new_n519), .ZN(new_n530));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G651), .ZN(new_n533));
  INV_X1    g108(.A(new_n508), .ZN(new_n534));
  AOI22_X1  g109(.A1(G52), .A2(new_n522), .B1(new_n534), .B2(G90), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT70), .B(G81), .Z(new_n539));
  OAI22_X1  g114(.A1(new_n502), .A2(new_n538), .B1(new_n508), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n530), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n540), .B1(new_n543), .B2(G651), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  NAND2_X1  g124(.A1(new_n534), .A2(G91), .ZN(new_n550));
  OAI211_X1 g125(.A(G53), .B(G543), .C1(new_n506), .C2(new_n507), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(KEYINPUT9), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT9), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n501), .A2(new_n553), .A3(G53), .A4(G543), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g130(.A(G65), .B1(new_n505), .B2(new_n504), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n556), .A2(KEYINPUT71), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G651), .ZN(new_n559));
  AOI21_X1  g134(.A(KEYINPUT71), .B1(new_n556), .B2(new_n557), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n550), .B(new_n555), .C1(new_n559), .C2(new_n560), .ZN(G299));
  INV_X1    g136(.A(new_n515), .ZN(new_n562));
  INV_X1    g137(.A(new_n527), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n526), .B1(new_n521), .B2(new_n523), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(G286));
  INV_X1    g140(.A(G166), .ZN(G303));
  INV_X1    g141(.A(G74), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n499), .B1(new_n530), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(G49), .ZN(new_n569));
  INV_X1    g144(.A(G87), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n502), .A2(new_n569), .B1(new_n508), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G288));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n495), .B2(new_n496), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n497), .A2(new_n501), .A3(G86), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n501), .A2(G48), .A3(G543), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n582), .A2(new_n499), .ZN(new_n583));
  AOI22_X1  g158(.A1(G47), .A2(new_n522), .B1(new_n534), .B2(G85), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n534), .A2(G92), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT10), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G66), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n518), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(G54), .A2(new_n522), .B1(new_n592), .B2(G651), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n586), .B1(new_n595), .B2(G868), .ZN(G284));
  OAI21_X1  g171(.A(new_n586), .B1(new_n595), .B2(G868), .ZN(G321));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(G299), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(G168), .B2(new_n598), .ZN(G297));
  OAI21_X1  g175(.A(new_n599), .B1(G168), .B2(new_n598), .ZN(G280));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n595), .B1(new_n602), .B2(G860), .ZN(G148));
  NAND2_X1  g178(.A1(new_n595), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n605), .A2(KEYINPUT72), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(KEYINPUT72), .ZN(new_n607));
  OAI211_X1 g182(.A(new_n606), .B(new_n607), .C1(G868), .C2(new_n544), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g184(.A1(new_n460), .A2(new_n461), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(new_n478), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  INV_X1    g188(.A(G2100), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n473), .A2(G123), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n459), .A2(G111), .ZN(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n619));
  INV_X1    g194(.A(G135), .ZN(new_n620));
  OAI221_X1 g195(.A(new_n617), .B1(new_n618), .B2(new_n619), .C1(new_n620), .C2(new_n479), .ZN(new_n621));
  INV_X1    g196(.A(G2096), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n615), .A2(new_n616), .A3(new_n623), .ZN(G156));
  XNOR2_X1  g199(.A(G2427), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2430), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2435), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n628), .A2(KEYINPUT14), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2451), .B(G2454), .Z(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n632), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT74), .Z(new_n640));
  OAI21_X1  g215(.A(KEYINPUT75), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT75), .ZN(new_n642));
  INV_X1    g217(.A(new_n640), .ZN(new_n643));
  NAND4_X1  g218(.A1(new_n636), .A2(new_n642), .A3(new_n643), .A4(new_n637), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(G14), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(new_n638), .B2(new_n640), .ZN(new_n647));
  AND2_X1   g222(.A1(new_n645), .A2(new_n647), .ZN(G401));
  INV_X1    g223(.A(KEYINPUT18), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(new_n614), .ZN(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n652), .B2(KEYINPUT18), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(new_n622), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(G227));
  XNOR2_X1  g235(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT76), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT19), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  AND2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT20), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n666), .A2(new_n667), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  MUX2_X1   g248(.A(new_n673), .B(new_n672), .S(new_n665), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(G1981), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(G1986), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n675), .B(G1981), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n680), .A2(G1986), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n662), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1991), .B(G1996), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(G1986), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n677), .A2(new_n678), .ZN(new_n685));
  INV_X1    g260(.A(new_n662), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  AND3_X1   g262(.A1(new_n682), .A2(new_n683), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n683), .B1(new_n682), .B2(new_n687), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(G229));
  MUX2_X1   g265(.A(G6), .B(G305), .S(G16), .Z(new_n691));
  XOR2_X1   g266(.A(KEYINPUT32), .B(G1981), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G22), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G166), .B2(new_n694), .ZN(new_n696));
  INV_X1    g271(.A(G1971), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n693), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT33), .B(G1976), .Z(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n694), .A2(G23), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(new_n572), .B2(new_n694), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT79), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n699), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n701), .B2(new_n704), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n706), .A2(KEYINPUT34), .ZN(new_n707));
  INV_X1    g282(.A(G290), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G16), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G16), .B2(G24), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n710), .A2(new_n678), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n678), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n473), .A2(G119), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n459), .A2(G107), .ZN(new_n714));
  OAI21_X1  g289(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n715));
  INV_X1    g290(.A(G131), .ZN(new_n716));
  OAI221_X1 g291(.A(new_n713), .B1(new_n714), .B2(new_n715), .C1(new_n716), .C2(new_n479), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT78), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT77), .B(G29), .Z(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G25), .B2(new_n720), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT35), .B(G1991), .Z(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  NOR4_X1   g300(.A1(new_n711), .A2(new_n712), .A3(new_n724), .A4(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n706), .A2(KEYINPUT34), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n707), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT80), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(KEYINPUT36), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT36), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n694), .A2(G21), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G168), .B2(new_n694), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT84), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1966), .ZN(new_n737));
  AOI22_X1  g312(.A1(G141), .A2(new_n480), .B1(new_n610), .B2(G105), .ZN(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT26), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G129), .B2(new_n473), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G29), .ZN(new_n743));
  OR3_X1    g318(.A1(new_n742), .A2(KEYINPUT82), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  OAI21_X1  g320(.A(KEYINPUT82), .B1(G29), .B2(G32), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT27), .B(G1996), .Z(new_n748));
  NOR2_X1   g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT83), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n747), .A2(new_n748), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT31), .B(G11), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT30), .B(G28), .Z(new_n753));
  OAI221_X1 g328(.A(new_n752), .B1(G29), .B2(new_n753), .C1(new_n621), .C2(new_n719), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n743), .A2(G33), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT25), .ZN(new_n756));
  NAND2_X1  g331(.A1(G103), .A2(G2104), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(G2105), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n459), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n478), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(new_n459), .ZN(new_n762));
  AOI211_X1 g337(.A(new_n760), .B(new_n762), .C1(G139), .C2(new_n480), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n755), .B1(new_n763), .B2(new_n743), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n754), .B1(new_n764), .B2(G2072), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT24), .B(G34), .ZN(new_n766));
  AOI22_X1  g341(.A1(G160), .A2(G29), .B1(new_n719), .B2(new_n766), .ZN(new_n767));
  OAI221_X1 g342(.A(new_n765), .B1(G2072), .B2(new_n764), .C1(G2084), .C2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(G2084), .ZN(new_n769));
  NAND2_X1  g344(.A1(G164), .A2(new_n720), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G27), .B2(new_n720), .ZN(new_n771));
  INV_X1    g346(.A(G2078), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n769), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n772), .B2(new_n771), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n694), .A2(G5), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G171), .B2(new_n694), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n774), .B1(G1961), .B2(new_n776), .ZN(new_n777));
  NOR4_X1   g352(.A1(new_n750), .A2(new_n751), .A3(new_n768), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(G1961), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT85), .Z(new_n780));
  NAND3_X1  g355(.A1(new_n737), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n781), .A2(KEYINPUT86), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(KEYINPUT86), .ZN(new_n783));
  NOR2_X1   g358(.A1(G4), .A2(G16), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n595), .B2(G16), .ZN(new_n785));
  INV_X1    g360(.A(G1348), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n719), .A2(G26), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT28), .Z(new_n789));
  NAND2_X1  g364(.A1(new_n473), .A2(G128), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT81), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n793));
  INV_X1    g368(.A(G116), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(G2105), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n480), .B2(G140), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n789), .B1(new_n797), .B2(G29), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2067), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n720), .A2(G35), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G162), .B2(new_n720), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT29), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n787), .B(new_n799), .C1(G2090), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(G2090), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT87), .Z(new_n805));
  NAND2_X1  g380(.A1(new_n694), .A2(G19), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n544), .B2(new_n694), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1341), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT88), .B(KEYINPUT23), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n694), .A2(G20), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G299), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(new_n694), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1956), .ZN(new_n814));
  NOR4_X1   g389(.A1(new_n803), .A2(new_n805), .A3(new_n808), .A4(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n782), .A2(new_n783), .A3(new_n815), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n731), .A2(new_n733), .A3(new_n816), .ZN(G311));
  NOR2_X1   g392(.A1(new_n733), .A2(new_n816), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(KEYINPUT36), .B2(new_n730), .ZN(G150));
  NAND2_X1  g394(.A1(new_n595), .A2(G559), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT89), .B(G55), .ZN(new_n822));
  INV_X1    g397(.A(G93), .ZN(new_n823));
  OAI22_X1  g398(.A1(new_n502), .A2(new_n822), .B1(new_n508), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(G80), .A2(G543), .ZN(new_n825));
  INV_X1    g400(.A(G67), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n530), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n824), .B1(new_n827), .B2(G651), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n544), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n544), .A2(new_n828), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n821), .B(new_n831), .Z(new_n832));
  AND2_X1   g407(.A1(new_n832), .A2(KEYINPUT39), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(KEYINPUT39), .ZN(new_n834));
  NOR3_X1   g409(.A1(new_n833), .A2(new_n834), .A3(G860), .ZN(new_n835));
  INV_X1    g410(.A(new_n828), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G860), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT90), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  OR2_X1    g414(.A1(new_n835), .A2(new_n839), .ZN(G145));
  XNOR2_X1  g415(.A(new_n797), .B(new_n742), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G164), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n763), .A2(KEYINPUT92), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT91), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n473), .A2(G130), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n459), .A2(G118), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(G142), .B2(new_n480), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n612), .B(new_n850), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n717), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n842), .A2(new_n844), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n845), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n854), .A2(KEYINPUT94), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(KEYINPUT94), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n842), .B(new_n844), .ZN(new_n857));
  INV_X1    g432(.A(new_n852), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n621), .B(G160), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(G162), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n855), .A2(new_n856), .A3(new_n859), .A4(new_n862), .ZN(new_n863));
  XOR2_X1   g438(.A(KEYINPUT93), .B(G37), .Z(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n859), .A2(new_n854), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n865), .B1(new_n866), .B2(new_n861), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g444(.A(KEYINPUT98), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n831), .B(new_n604), .ZN(new_n871));
  NAND2_X1  g446(.A1(G299), .A2(KEYINPUT95), .ZN(new_n872));
  OR2_X1    g447(.A1(G299), .A2(KEYINPUT95), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n595), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n594), .A2(KEYINPUT95), .A3(G299), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT96), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(KEYINPUT41), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT41), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n876), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n884), .A2(new_n871), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n870), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n572), .B(KEYINPUT97), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(G305), .ZN(new_n888));
  XNOR2_X1  g463(.A(G290), .B(G166), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT42), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n880), .A2(new_n885), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n892), .A2(KEYINPUT98), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n886), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n891), .A2(new_n870), .A3(new_n885), .A4(new_n880), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(G868), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n894), .A2(KEYINPUT99), .A3(new_n896), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n894), .A2(new_n896), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT99), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n899), .B1(new_n836), .B2(new_n598), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n897), .B1(new_n898), .B2(new_n900), .ZN(G295));
  AOI21_X1  g476(.A(new_n897), .B1(new_n898), .B2(new_n900), .ZN(G331));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT102), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n905));
  NAND2_X1  g480(.A1(G301), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n831), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n829), .A2(new_n830), .A3(new_n906), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(G301), .A2(new_n905), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT101), .B1(G286), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(G171), .A2(KEYINPUT100), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT101), .ZN(new_n914));
  NAND3_X1  g489(.A1(G168), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n910), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n908), .A2(new_n912), .A3(new_n915), .A4(new_n909), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n876), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n917), .A2(new_n881), .A3(new_n883), .A4(new_n918), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n904), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n904), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n922), .A2(new_n924), .A3(new_n890), .ZN(new_n925));
  INV_X1    g500(.A(new_n921), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n890), .B1(new_n926), .B2(new_n919), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n864), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n903), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n890), .B1(new_n922), .B2(new_n924), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT102), .B1(new_n926), .B2(new_n919), .ZN(new_n931));
  INV_X1    g506(.A(new_n890), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n932), .A3(new_n923), .ZN(new_n933));
  INV_X1    g508(.A(G37), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n930), .A2(new_n933), .A3(KEYINPUT43), .A4(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT44), .B1(new_n929), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n925), .A2(G37), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n937), .A2(KEYINPUT103), .A3(new_n903), .A4(new_n930), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT43), .B1(new_n925), .B2(new_n928), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n930), .A2(new_n933), .A3(new_n903), .A4(new_n934), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT103), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n938), .A2(new_n939), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n936), .B1(new_n943), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g519(.A(KEYINPUT45), .ZN(new_n945));
  XOR2_X1   g520(.A(KEYINPUT104), .B(G1384), .Z(new_n946));
  OAI21_X1  g521(.A(new_n945), .B1(G164), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n469), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n948), .A2(G40), .A3(new_n462), .A4(new_n465), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n797), .A2(G2067), .ZN(new_n952));
  INV_X1    g527(.A(G2067), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n792), .A2(new_n953), .A3(new_n796), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G1996), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n742), .B(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n955), .A2(new_n723), .A3(new_n718), .A4(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n951), .B1(new_n958), .B2(new_n954), .ZN(new_n959));
  XOR2_X1   g534(.A(new_n959), .B(KEYINPUT125), .Z(new_n960));
  NAND3_X1  g535(.A1(new_n708), .A2(new_n678), .A3(new_n950), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT48), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n717), .B(KEYINPUT105), .ZN(new_n963));
  XOR2_X1   g538(.A(new_n963), .B(new_n723), .Z(new_n964));
  NAND2_X1  g539(.A1(new_n955), .A2(new_n957), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n962), .B1(new_n951), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n955), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n950), .B1(new_n968), .B2(new_n742), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n950), .A2(new_n956), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT46), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g547(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n973));
  OAI21_X1  g548(.A(new_n967), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AOI211_X1 g549(.A(new_n960), .B(new_n974), .C1(new_n972), .C2(new_n973), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT61), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n977));
  INV_X1    g552(.A(new_n560), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n978), .A2(G651), .A3(new_n558), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n552), .A2(new_n554), .B1(new_n534), .B2(G91), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n982), .B1(new_n979), .B2(new_n980), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT57), .ZN(new_n984));
  OAI22_X1  g559(.A1(KEYINPUT113), .A2(new_n981), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT113), .B1(G299), .B2(KEYINPUT112), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT57), .ZN(new_n987));
  INV_X1    g562(.A(G1384), .ZN(new_n988));
  INV_X1    g563(.A(new_n493), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n492), .B1(new_n478), .B2(new_n489), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n988), .B1(new_n991), .B2(new_n487), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n949), .B1(new_n992), .B2(KEYINPUT50), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT50), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n994), .B(new_n988), .C1(new_n991), .C2(new_n487), .ZN(new_n995));
  AOI21_X1  g570(.A(G1956), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G40), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n466), .A2(new_n469), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n945), .B1(G164), .B2(G1384), .ZN(new_n999));
  INV_X1    g574(.A(new_n946), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT45), .B(new_n1000), .C1(new_n991), .C2(new_n487), .ZN(new_n1001));
  XNOR2_X1  g576(.A(KEYINPUT56), .B(G2072), .ZN(new_n1002));
  AND4_X1   g577(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n985), .B(new_n987), .C1(new_n996), .C2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(new_n998), .A3(new_n995), .ZN(new_n1006));
  INV_X1    g581(.A(G1956), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n949), .B1(new_n992), .B2(new_n945), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1009), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n984), .B1(G299), .B2(KEYINPUT113), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n986), .A2(new_n1011), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n981), .A2(KEYINPUT113), .A3(new_n984), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1008), .B(new_n1010), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n976), .B1(new_n1004), .B2(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1004), .A2(new_n1014), .A3(new_n976), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT59), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n999), .A2(new_n1001), .A3(new_n956), .A4(new_n998), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n491), .A2(new_n493), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n482), .A2(new_n486), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1384), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n998), .ZN(new_n1022));
  XOR2_X1   g597(.A(KEYINPUT58), .B(G1341), .Z(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1018), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1018), .A2(KEYINPUT116), .A3(new_n1024), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1017), .B1(new_n1029), .B2(new_n544), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1018), .A2(KEYINPUT116), .A3(new_n1024), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT116), .B1(new_n1018), .B2(new_n1024), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1017), .B(new_n544), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  OAI22_X1  g609(.A1(new_n1015), .A2(new_n1016), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1021), .A2(new_n998), .A3(new_n953), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1036), .B1(new_n1006), .B2(new_n786), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(KEYINPUT60), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n998), .B1(new_n1021), .B2(new_n994), .ZN(new_n1041));
  NOR3_X1   g616(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n786), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1036), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(KEYINPUT60), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT117), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n595), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(KEYINPUT117), .A3(new_n594), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1040), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1037), .A2(KEYINPUT60), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT118), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI211_X1 g626(.A(new_n1038), .B(new_n595), .C1(new_n1037), .C2(KEYINPUT60), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n594), .B1(new_n1045), .B2(KEYINPUT117), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1039), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1050), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1035), .B1(new_n1051), .B2(new_n1057), .ZN(new_n1058));
  OR3_X1    g633(.A1(new_n1037), .A2(KEYINPUT114), .A3(new_n594), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT114), .B1(new_n1037), .B2(new_n594), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(new_n1004), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT115), .B1(new_n1061), .B2(new_n1014), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1061), .A2(KEYINPUT115), .A3(new_n1014), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT119), .B1(new_n1058), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1030), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1015), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1004), .A2(new_n1014), .A3(new_n976), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1067), .A2(new_n1033), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1055), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1064), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(new_n1062), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G8), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1078), .B1(new_n1021), .B2(new_n998), .ZN(new_n1079));
  INV_X1    g654(.A(G1976), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1079), .B1(G288), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT52), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n572), .B2(G1976), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1082), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n578), .A2(new_n676), .A3(new_n579), .A4(new_n580), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT107), .ZN(new_n1087));
  OAI21_X1  g662(.A(G61), .B1(new_n505), .B2(new_n504), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n499), .B1(new_n1088), .B2(new_n576), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n579), .A2(new_n580), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1089), .B1(new_n1090), .B2(KEYINPUT106), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT106), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n579), .A2(new_n580), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1087), .B1(new_n1094), .B2(G1981), .ZN(new_n1095));
  AOI211_X1 g670(.A(KEYINPUT107), .B(new_n676), .C1(new_n1091), .C2(new_n1093), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT49), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT108), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT108), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1099), .B(KEYINPUT49), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1095), .A2(new_n1096), .A3(KEYINPUT49), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1079), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1085), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n999), .A2(new_n1001), .A3(new_n772), .A4(new_n998), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT121), .B(G1961), .Z(new_n1109));
  AOI22_X1  g684(.A1(new_n1107), .A2(new_n1108), .B1(new_n1006), .B2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(KEYINPUT45), .B(new_n988), .C1(new_n991), .C2(new_n487), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT111), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1021), .A2(new_n1113), .A3(KEYINPUT45), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT110), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n482), .B(new_n486), .C1(new_n989), .C2(new_n990), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT45), .B1(new_n1117), .B2(new_n988), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1116), .B1(new_n1118), .B2(new_n949), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n999), .A2(KEYINPUT110), .A3(new_n998), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1107), .A2(G2078), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1115), .A2(new_n1119), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(G301), .B1(new_n1110), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1108), .A2(new_n1107), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1006), .A2(new_n1109), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1121), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n946), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1126), .B1(new_n1127), .B2(KEYINPUT45), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n949), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n998), .A2(KEYINPUT122), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1128), .A2(new_n1130), .A3(new_n1131), .A4(new_n947), .ZN(new_n1132));
  AND4_X1   g707(.A1(G301), .A2(new_n1124), .A3(new_n1125), .A4(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1106), .B1(new_n1123), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(G1971), .B1(new_n1009), .B2(new_n1001), .ZN(new_n1135));
  INV_X1    g710(.A(G2090), .ZN(new_n1136));
  AND4_X1   g711(.A1(new_n1136), .A2(new_n1005), .A3(new_n998), .A4(new_n995), .ZN(new_n1137));
  OAI21_X1  g712(.A(G8), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(G8), .B1(new_n500), .B2(new_n510), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT55), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1139), .B(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1138), .A2(KEYINPUT109), .A3(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(G8), .B(new_n1141), .C1(new_n1135), .C2(new_n1137), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT109), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1105), .A2(new_n1134), .A3(new_n1143), .A4(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1110), .A2(new_n1122), .A3(G301), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT54), .ZN(new_n1150));
  AOI21_X1  g725(.A(KEYINPUT123), .B1(new_n1110), .B2(new_n1132), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1151), .A2(G301), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1110), .A2(KEYINPUT123), .A3(new_n1132), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1150), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1148), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT51), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1115), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1157));
  INV_X1    g732(.A(G1966), .ZN(new_n1158));
  INV_X1    g733(.A(G2084), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1006), .ZN(new_n1160));
  AOI22_X1  g735(.A1(new_n1157), .A2(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1078), .B1(new_n1161), .B2(G168), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1160), .A2(new_n1159), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(G286), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1156), .B1(new_n1162), .B2(new_n1166), .ZN(new_n1167));
  AOI211_X1 g742(.A(KEYINPUT51), .B(new_n1078), .C1(new_n1161), .C2(G168), .ZN(new_n1168));
  OAI21_X1  g743(.A(KEYINPUT120), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1163), .A2(G168), .A3(new_n1164), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(G8), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1161), .A2(G168), .ZN(new_n1172));
  OAI21_X1  g747(.A(KEYINPUT51), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT120), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1162), .A2(new_n1156), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  AND3_X1   g751(.A1(new_n1155), .A2(new_n1169), .A3(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1066), .A2(new_n1077), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1169), .A2(new_n1176), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT62), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1169), .A2(new_n1176), .A3(KEYINPUT62), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1105), .A2(new_n1143), .A3(new_n1147), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n1183), .A2(new_n1123), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1181), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1144), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1105), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1086), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1189));
  NOR2_X1   g764(.A1(G288), .A2(G1976), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1187), .B1(new_n1191), .B2(new_n1103), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1161), .A2(new_n1078), .A3(G286), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1183), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT63), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1186), .A2(new_n1195), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1105), .A2(new_n1193), .A3(new_n1197), .A4(new_n1146), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1192), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1178), .A2(new_n1185), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT124), .ZN(new_n1201));
  INV_X1    g776(.A(new_n966), .ZN(new_n1202));
  XNOR2_X1  g777(.A(G290), .B(G1986), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n950), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  AND3_X1   g779(.A1(new_n1200), .A2(new_n1201), .A3(new_n1204), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1201), .B1(new_n1200), .B2(new_n1204), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n975), .B1(new_n1205), .B2(new_n1206), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g782(.A(G319), .ZN(new_n1209));
  OR2_X1    g783(.A1(G227), .A2(new_n1209), .ZN(new_n1210));
  NOR3_X1   g784(.A1(G229), .A2(G401), .A3(new_n1210), .ZN(new_n1211));
  NAND4_X1  g785(.A1(new_n929), .A2(new_n935), .A3(new_n868), .A4(new_n1211), .ZN(new_n1212));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n1213));
  XNOR2_X1  g787(.A(new_n1212), .B(new_n1213), .ZN(G308));
  XNOR2_X1  g788(.A(new_n1212), .B(KEYINPUT127), .ZN(G225));
endmodule


