//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 1 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n570, new_n571, new_n572, new_n573, new_n575,
    new_n576, new_n577, new_n578, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT64), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  INV_X1    g034(.A(new_n455), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n459), .A2(G2106), .B1(G567), .B2(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n463), .B(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G101), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(new_n462), .ZN(new_n469));
  OAI22_X1  g044(.A1(new_n465), .A2(new_n466), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n471), .B1(new_n468), .B2(G125), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(new_n462), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n468), .A2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n476), .A2(G124), .B1(new_n480), .B2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT66), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT67), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND3_X1  g062(.A1(new_n462), .A2(G102), .A3(G2104), .ZN(new_n488));
  AOI22_X1  g063(.A1(new_n468), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(new_n462), .ZN(new_n490));
  OAI211_X1 g065(.A(G138), .B(new_n462), .C1(new_n477), .C2(new_n478), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n468), .A2(KEYINPUT4), .A3(G138), .A4(new_n462), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n490), .A2(new_n495), .ZN(G164));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(G651), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(KEYINPUT68), .A3(KEYINPUT6), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n499), .A2(new_n501), .B1(new_n498), .B2(G651), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OR2_X1    g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n500), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G62), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n499), .A2(new_n501), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n498), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n506), .A2(new_n507), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n509), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n505), .A2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT7), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT7), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n520), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n508), .A2(G63), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n510), .A2(G89), .A3(new_n512), .A4(new_n511), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n510), .A2(G51), .A3(G543), .A4(new_n511), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(G168));
  INV_X1    g101(.A(G64), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n527), .B1(new_n506), .B2(new_n507), .ZN(new_n528));
  AND2_X1   g103(.A1(G77), .A2(G543), .ZN(new_n529));
  OAI21_X1  g104(.A(G651), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n510), .A2(G90), .A3(new_n512), .A4(new_n511), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n510), .A2(G52), .A3(G543), .A4(new_n511), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(G171));
  NAND3_X1  g109(.A1(new_n502), .A2(G81), .A3(new_n512), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n502), .A2(G43), .A3(G543), .ZN(new_n536));
  INV_X1    g111(.A(G56), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(new_n506), .B2(new_n507), .ZN(new_n538));
  AND2_X1   g113(.A1(G68), .A2(G543), .ZN(new_n539));
  OAI21_X1  g114(.A(G651), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n535), .A2(new_n536), .A3(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  NAND4_X1  g122(.A1(new_n510), .A2(G53), .A3(G543), .A4(new_n511), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT9), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g125(.A1(new_n502), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT69), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT70), .ZN(new_n555));
  INV_X1    g130(.A(G91), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n513), .B2(new_n556), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n502), .A2(KEYINPUT70), .A3(G91), .A4(new_n512), .ZN(new_n558));
  AND2_X1   g133(.A1(KEYINPUT5), .A2(G543), .ZN(new_n559));
  NOR2_X1   g134(.A1(KEYINPUT5), .A2(G543), .ZN(new_n560));
  OAI21_X1  g135(.A(G65), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT71), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n500), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n561), .A2(KEYINPUT71), .A3(new_n562), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n557), .A2(new_n558), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n550), .A2(KEYINPUT69), .A3(new_n551), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n554), .A2(new_n567), .A3(new_n568), .ZN(G299));
  NAND2_X1  g144(.A1(new_n533), .A2(KEYINPUT72), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT72), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n530), .A2(new_n531), .A3(new_n532), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G301));
  INV_X1    g149(.A(KEYINPUT73), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n525), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n522), .A2(new_n523), .A3(new_n524), .A4(KEYINPUT73), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G286));
  AND2_X1   g154(.A1(new_n502), .A2(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G49), .ZN(new_n581));
  INV_X1    g156(.A(new_n513), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G87), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(G288));
  NAND2_X1  g160(.A1(new_n580), .A2(G48), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(new_n500), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n582), .A2(G86), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n500), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT74), .ZN(new_n593));
  AOI22_X1  g168(.A1(G47), .A2(new_n580), .B1(new_n582), .B2(G85), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(new_n512), .A2(G66), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n500), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(new_n580), .B2(G54), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  INV_X1    g175(.A(G92), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n513), .B2(new_n601), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n502), .A2(KEYINPUT10), .A3(G92), .A4(new_n512), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(G868), .B2(new_n573), .ZN(G321));
  XNOR2_X1  g182(.A(G321), .B(KEYINPUT75), .ZN(G284));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  MUX2_X1   g184(.A(G286), .B(G299), .S(new_n609), .Z(G297));
  XNOR2_X1  g185(.A(G297), .B(KEYINPUT76), .ZN(G280));
  INV_X1    g186(.A(new_n605), .ZN(new_n612));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n541), .A2(new_n609), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n605), .A2(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(new_n609), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n476), .A2(G123), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT77), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n480), .A2(G135), .ZN(new_n621));
  NOR2_X1   g196(.A1(G99), .A2(G2105), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n620), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(G2096), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n463), .B(KEYINPUT65), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(new_n468), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  INV_X1    g205(.A(G2100), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n626), .A2(new_n632), .A3(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n640), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT78), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n648), .B(G14), .C1(new_n646), .C2(new_n645), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT79), .ZN(G401));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT80), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  NOR2_X1   g229(.A1(G2072), .A2(G2078), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n444), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n653), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT18), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(KEYINPUT17), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n660), .A2(new_n652), .A3(new_n654), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT81), .Z(new_n662));
  INV_X1    g237(.A(new_n660), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n654), .B1(new_n663), .B2(new_n653), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n653), .B2(new_n657), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n659), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(new_n625), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2100), .ZN(G227));
  XOR2_X1   g243(.A(G1971), .B(G1976), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n673), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT20), .Z(new_n677));
  AOI211_X1 g252(.A(new_n675), .B(new_n677), .C1(new_n670), .C2(new_n674), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  INV_X1    g254(.A(G1981), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n678), .B(new_n683), .Z(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT82), .B(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(G229));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n688), .A2(G24), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(G290), .B2(G16), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT85), .ZN(new_n691));
  INV_X1    g266(.A(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(KEYINPUT86), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n691), .B(G1986), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT86), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G25), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n476), .A2(G119), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(G95), .A2(G2105), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n702), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT83), .Z(new_n704));
  AOI211_X1 g279(.A(new_n701), .B(new_n704), .C1(G131), .C2(new_n480), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n699), .B1(new_n705), .B2(new_n698), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT84), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT35), .B(G1991), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n694), .A2(new_n697), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n688), .A2(G6), .ZN(new_n711));
  INV_X1    g286(.A(G305), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(new_n688), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT87), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT32), .B(G1981), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT88), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n714), .A2(new_n717), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n688), .A2(G22), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G166), .B2(new_n688), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT90), .B(G1971), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(G16), .A2(G23), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT89), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G288), .B2(new_n688), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT33), .B(G1976), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n718), .A2(new_n719), .A3(new_n723), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT34), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n710), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT36), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT99), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n688), .A2(G4), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n612), .B2(new_n688), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1348), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n688), .A2(G19), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n542), .B2(new_n688), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1341), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n476), .A2(G128), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n480), .A2(G140), .ZN(new_n742));
  NOR2_X1   g317(.A1(G104), .A2(G2105), .ZN(new_n743));
  OAI21_X1  g318(.A(G2104), .B1(new_n462), .B2(G116), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n741), .B(new_n742), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n698), .A2(G26), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT28), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G2067), .ZN(new_n750));
  NOR3_X1   g325(.A1(new_n737), .A2(new_n740), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT91), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n698), .A2(G32), .ZN(new_n753));
  NAND3_X1  g328(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT26), .Z(new_n755));
  INV_X1    g330(.A(G129), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n475), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n480), .A2(G141), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT93), .ZN(new_n759));
  AOI211_X1 g334(.A(new_n757), .B(new_n759), .C1(G105), .C2(new_n627), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n753), .B1(new_n760), .B2(new_n698), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT27), .B(G1996), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT31), .B(G11), .Z(new_n764));
  INV_X1    g339(.A(KEYINPUT30), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n698), .B1(new_n765), .B2(G28), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT95), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n766), .A2(new_n767), .B1(new_n765), .B2(G28), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n764), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n624), .B2(new_n698), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT96), .ZN(new_n772));
  NOR2_X1   g347(.A1(G171), .A2(new_n688), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G5), .B2(new_n688), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G168), .A2(new_n688), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n688), .B2(G21), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT94), .B(G1966), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n775), .A2(G1961), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n763), .A2(new_n772), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n698), .A2(G35), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G162), .B2(new_n698), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT29), .B(G2090), .Z(new_n783));
  XOR2_X1   g358(.A(new_n782), .B(new_n783), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n480), .A2(G139), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT92), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT25), .Z(new_n788));
  AOI22_X1  g363(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(new_n462), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(new_n698), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n698), .B2(G33), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n793), .A2(new_n442), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n442), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT24), .ZN(new_n796));
  INV_X1    g371(.A(G34), .ZN(new_n797));
  AOI21_X1  g372(.A(G29), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n796), .B2(new_n797), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G160), .B2(new_n698), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G2084), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n794), .A2(new_n795), .A3(new_n801), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n780), .A2(new_n784), .A3(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT98), .B(KEYINPUT23), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n688), .A2(G20), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G299), .B2(G16), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1956), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n800), .A2(G2084), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT97), .ZN(new_n810));
  OAI22_X1  g385(.A1(new_n775), .A2(G1961), .B1(new_n777), .B2(new_n778), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n698), .A2(G27), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G164), .B2(new_n698), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G2078), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n810), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  AND4_X1   g390(.A1(new_n752), .A2(new_n803), .A3(new_n808), .A4(new_n815), .ZN(new_n816));
  AND3_X1   g391(.A1(new_n733), .A2(new_n734), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n734), .B1(new_n733), .B2(new_n816), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(G311));
  NAND2_X1  g394(.A1(new_n733), .A2(new_n816), .ZN(G150));
  NAND4_X1  g395(.A1(new_n510), .A2(G55), .A3(G543), .A4(new_n511), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n510), .A2(G93), .A3(new_n512), .A4(new_n511), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT101), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(G67), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n506), .B2(new_n507), .ZN(new_n826));
  AND2_X1   g401(.A1(G80), .A2(G543), .ZN(new_n827));
  OAI21_X1  g402(.A(G651), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT100), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g405(.A(KEYINPUT100), .B(G651), .C1(new_n826), .C2(new_n827), .ZN(new_n831));
  AND3_X1   g406(.A1(new_n824), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT102), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n823), .B1(new_n821), .B2(new_n822), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n832), .A2(new_n833), .A3(new_n542), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n541), .A2(KEYINPUT102), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n535), .A2(new_n536), .A3(new_n833), .A4(new_n540), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n824), .A2(new_n830), .A3(new_n831), .ZN(new_n839));
  OAI211_X1 g414(.A(new_n837), .B(new_n838), .C1(new_n839), .C2(new_n834), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT38), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n612), .A2(G559), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n844), .A2(KEYINPUT39), .ZN(new_n845));
  INV_X1    g420(.A(G860), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(KEYINPUT39), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n846), .B1(new_n832), .B2(new_n835), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT37), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT103), .ZN(G145));
  INV_X1    g427(.A(KEYINPUT104), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n853), .B(new_n488), .C1(new_n489), .C2(new_n462), .ZN(new_n854));
  OAI21_X1  g429(.A(G126), .B1(new_n477), .B2(new_n478), .ZN(new_n855));
  NAND2_X1  g430(.A1(G114), .A2(G2104), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n462), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n488), .ZN(new_n858));
  OAI21_X1  g433(.A(KEYINPUT104), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n493), .A2(new_n494), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n854), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n745), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n791), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(new_n760), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n705), .B(new_n629), .ZN(new_n865));
  INV_X1    g440(.A(G130), .ZN(new_n866));
  NOR2_X1   g441(.A1(G106), .A2(G2105), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n868));
  OAI22_X1  g443(.A1(new_n475), .A2(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(G142), .B2(new_n480), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n865), .B(new_n870), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n871), .A2(KEYINPUT105), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(KEYINPUT105), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n864), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(new_n864), .B2(new_n873), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n624), .B(G160), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(G162), .ZN(new_n877));
  AOI21_X1  g452(.A(G37), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(new_n877), .B2(new_n875), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g455(.A(new_n609), .B1(new_n839), .B2(new_n834), .ZN(new_n881));
  XNOR2_X1  g456(.A(G290), .B(G305), .ZN(new_n882));
  XOR2_X1   g457(.A(G303), .B(G288), .Z(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n884), .B(KEYINPUT42), .Z(new_n885));
  XOR2_X1   g460(.A(new_n841), .B(new_n616), .Z(new_n886));
  NAND2_X1  g461(.A1(G299), .A2(new_n612), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT106), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n605), .A2(new_n568), .A3(new_n567), .A4(new_n554), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(G299), .A2(new_n612), .A3(KEYINPUT106), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n890), .A2(KEYINPUT107), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT107), .B1(new_n890), .B2(new_n891), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n886), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n890), .A2(new_n891), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT41), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n897));
  OR3_X1    g472(.A1(G299), .A2(new_n612), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n887), .A2(new_n897), .A3(new_n889), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n896), .B1(new_n900), .B2(KEYINPUT41), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n894), .B1(new_n902), .B2(new_n886), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n885), .B(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n881), .B1(new_n904), .B2(new_n609), .ZN(G295));
  OAI21_X1  g480(.A(new_n881), .B1(new_n904), .B2(new_n609), .ZN(G331));
  NAND3_X1  g481(.A1(new_n576), .A2(G171), .A3(new_n577), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n570), .A2(G168), .A3(new_n572), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n841), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n836), .A3(new_n840), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n913), .A2(new_n895), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT109), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n911), .A2(new_n915), .A3(new_n912), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n909), .A2(new_n836), .A3(KEYINPUT109), .A4(new_n840), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n914), .B1(new_n901), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n884), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(G37), .B1(new_n920), .B2(new_n921), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n920), .A2(new_n921), .ZN(new_n925));
  INV_X1    g500(.A(G37), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n918), .B1(new_n892), .B2(new_n893), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n895), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT41), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n930), .A2(KEYINPUT110), .A3(new_n913), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n895), .A2(new_n929), .B1(new_n912), .B2(new_n911), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT110), .B1(new_n934), .B2(new_n931), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n884), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g513(.A(KEYINPUT111), .B(new_n884), .C1(new_n933), .C2(new_n935), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n927), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  MUX2_X1   g516(.A(new_n924), .B(new_n940), .S(new_n941), .Z(new_n942));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT112), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(new_n940), .B2(new_n941), .ZN(new_n946));
  INV_X1    g521(.A(new_n939), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n930), .A2(new_n913), .A3(new_n931), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(new_n928), .A3(new_n932), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT111), .B1(new_n951), .B2(new_n884), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n923), .B1(new_n947), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n953), .A2(KEYINPUT112), .A3(KEYINPUT43), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n946), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n922), .A2(new_n923), .A3(new_n941), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT44), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT113), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT113), .ZN(new_n960));
  AOI211_X1 g535(.A(new_n960), .B(new_n957), .C1(new_n946), .C2(new_n954), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n944), .B1(new_n959), .B2(new_n961), .ZN(G397));
  INV_X1    g537(.A(KEYINPUT127), .ZN(new_n963));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT45), .B1(new_n861), .B2(new_n964), .ZN(new_n965));
  XOR2_X1   g540(.A(KEYINPUT114), .B(G40), .Z(new_n966));
  NOR3_X1   g541(.A1(new_n470), .A2(new_n473), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  OR3_X1    g543(.A1(new_n968), .A2(KEYINPUT115), .A3(G1996), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT115), .B1(new_n968), .B2(G1996), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n968), .ZN(new_n972));
  XOR2_X1   g547(.A(new_n745), .B(G2067), .Z(new_n973));
  INV_X1    g548(.A(G1996), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n973), .B1(new_n760), .B2(new_n974), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n971), .A2(new_n760), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n705), .A2(new_n708), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n705), .A2(new_n708), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n972), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n976), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(G290), .A2(G1986), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n692), .B1(new_n593), .B2(new_n594), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n972), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n967), .A2(new_n861), .A3(new_n964), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G8), .ZN(new_n988));
  INV_X1    g563(.A(G1976), .ZN(new_n989));
  NOR2_X1   g564(.A1(G288), .A2(new_n989), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n987), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT52), .B1(G288), .B2(new_n989), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n993), .B1(new_n994), .B2(new_n991), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n712), .A2(G1981), .ZN(new_n996));
  NAND2_X1  g571(.A1(G305), .A2(new_n680), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(KEYINPUT118), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT49), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n987), .A2(new_n988), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT49), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n996), .A2(new_n997), .A3(KEYINPUT118), .A4(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT119), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n999), .A2(KEYINPUT119), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n995), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n861), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n857), .A2(new_n858), .ZN(new_n1009));
  AOI21_X1  g584(.A(G1384), .B1(new_n860), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n967), .B1(new_n1010), .B2(KEYINPUT45), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT116), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  AOI22_X1  g587(.A1(G101), .A2(new_n627), .B1(new_n480), .B2(G137), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n468), .A2(G125), .ZN(new_n1014));
  OAI21_X1  g589(.A(G2105), .B1(new_n1014), .B2(new_n471), .ZN(new_n1015));
  INV_X1    g590(.A(new_n966), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n964), .B1(new_n490), .B2(new_n495), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n861), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(KEYINPUT117), .B(G1971), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1012), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1017), .B1(KEYINPUT50), .B2(new_n1019), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n861), .A2(new_n1027), .A3(new_n964), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n1029), .A2(G2090), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n988), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(G303), .A2(G8), .ZN(new_n1032));
  XOR2_X1   g607(.A(new_n1032), .B(KEYINPUT55), .Z(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1027), .B1(new_n861), .B2(new_n964), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1027), .B(new_n964), .C1(new_n490), .C2(new_n495), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n967), .ZN(new_n1037));
  OR3_X1    g612(.A1(new_n1035), .A2(new_n1037), .A3(G2090), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n988), .B1(new_n1025), .B2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1007), .B(new_n1034), .C1(new_n1033), .C2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1023), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1021), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n443), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g621(.A(KEYINPUT123), .B(G1961), .Z(new_n1047));
  AND3_X1   g622(.A1(new_n1026), .A2(KEYINPUT122), .A3(new_n1028), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT122), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n965), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1013), .B(KEYINPUT124), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1045), .A2(G2078), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1015), .A2(G40), .A3(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1051), .A2(new_n1022), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1046), .A2(G301), .A3(new_n1050), .A4(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n495), .B1(new_n490), .B2(KEYINPUT104), .ZN(new_n1057));
  AOI21_X1  g632(.A(G1384), .B1(new_n1057), .B2(new_n854), .ZN(new_n1058));
  OAI211_X1 g633(.A(KEYINPUT120), .B(new_n967), .C1(new_n1058), .C2(KEYINPUT45), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT120), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(new_n965), .B2(new_n1017), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1019), .A2(new_n1018), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1059), .A2(new_n1061), .A3(new_n1053), .A4(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(G2078), .B1(new_n1012), .B2(new_n1023), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1050), .B(new_n1064), .C1(new_n1065), .C2(KEYINPUT53), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n573), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1056), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1050), .B(new_n1055), .C1(new_n1065), .C2(KEYINPUT53), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G171), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT125), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n1066), .A2(new_n573), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1069), .B1(new_n1076), .B2(KEYINPUT54), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1059), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n778), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1029), .A2(G2084), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(G168), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(G8), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1080), .B1(new_n1078), .B2(new_n778), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(G168), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT51), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  AOI211_X1 g661(.A(KEYINPUT51), .B(new_n988), .C1(new_n1084), .C2(G168), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1956), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT56), .B(G2072), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1020), .A2(new_n1022), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n550), .A2(KEYINPUT121), .A3(new_n551), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT121), .B1(new_n550), .B2(new_n551), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n567), .B(new_n1095), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1091), .A2(new_n1093), .A3(new_n1094), .A4(new_n1098), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1099), .A2(new_n612), .ZN(new_n1100));
  INV_X1    g675(.A(G1348), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n986), .A2(G2067), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1100), .A2(new_n1105), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n605), .A4(new_n1104), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1020), .A2(new_n974), .A3(new_n1022), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT58), .B(G1341), .Z(new_n1111));
  NAND2_X1  g686(.A1(new_n986), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n542), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT59), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(new_n1116), .A3(new_n542), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1107), .A2(new_n1106), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT61), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1119), .A2(new_n1120), .A3(new_n1099), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1120), .B1(new_n1119), .B2(new_n1099), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1109), .B(new_n1118), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT60), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1028), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n967), .B1(new_n1010), .B2(new_n1027), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1026), .A2(KEYINPUT122), .A3(new_n1028), .ZN(new_n1129));
  AOI21_X1  g704(.A(G1348), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1124), .B1(new_n1130), .B2(new_n1103), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n1104), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1131), .A2(new_n1132), .A3(new_n612), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1108), .B1(new_n1123), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1089), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1077), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1086), .A2(new_n1088), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT51), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n988), .B1(new_n1084), .B2(G168), .ZN(new_n1140));
  INV_X1    g715(.A(new_n778), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n965), .A2(new_n1017), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1062), .B1(new_n1142), .B2(KEYINPUT120), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1141), .B1(new_n1143), .B2(new_n1061), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n525), .B1(new_n1144), .B2(new_n1080), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1139), .B1(new_n1140), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT62), .B1(new_n1146), .B2(new_n1087), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1067), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1138), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1041), .B1(new_n1136), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n1151));
  OAI211_X1 g726(.A(G8), .B(new_n578), .C1(new_n1144), .C2(new_n1080), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1151), .B1(new_n1040), .B2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1152), .A2(new_n1151), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1154), .A2(new_n1034), .A3(new_n1007), .A4(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1007), .A2(new_n1033), .A3(new_n1031), .ZN(new_n1158));
  AOI211_X1 g733(.A(G1976), .B(G288), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1159));
  NOR2_X1   g734(.A1(G305), .A2(G1981), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1000), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1157), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n985), .B1(new_n1150), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT46), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n971), .B(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n760), .A2(new_n973), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(new_n972), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT47), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1168), .B(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1170), .A2(KEYINPUT126), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n972), .A2(new_n982), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1172), .B(KEYINPUT48), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n981), .A2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n745), .A2(G2067), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1175), .B1(new_n976), .B2(new_n978), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1174), .B1(new_n968), .B2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1171), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1170), .A2(KEYINPUT126), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n963), .B1(new_n1163), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1179), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1182), .A2(new_n1171), .A3(new_n1177), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1157), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1138), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1185), .B1(new_n1077), .B2(new_n1135), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1184), .B1(new_n1041), .B2(new_n1186), .ZN(new_n1187));
  OAI211_X1 g762(.A(new_n1183), .B(KEYINPUT127), .C1(new_n1187), .C2(new_n985), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1181), .A2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g764(.A1(new_n686), .A2(G319), .ZN(new_n1191));
  NOR3_X1   g765(.A1(G401), .A2(G227), .A3(new_n1191), .ZN(new_n1192));
  NAND3_X1  g766(.A1(new_n1192), .A2(new_n879), .A3(new_n942), .ZN(G225));
  INV_X1    g767(.A(G225), .ZN(G308));
endmodule


