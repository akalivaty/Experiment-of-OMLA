//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n809, new_n810, new_n812, new_n813, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  INV_X1    g003(.A(G8gat), .ZN(new_n205));
  OAI221_X1 g004(.A(new_n204), .B1(KEYINPUT93), .B2(new_n205), .C1(G1gat), .C2(new_n202), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(KEYINPUT93), .ZN(new_n207));
  XOR2_X1   g006(.A(new_n206), .B(new_n207), .Z(new_n208));
  OR2_X1    g007(.A1(KEYINPUT91), .A2(G43gat), .ZN(new_n209));
  INV_X1    g008(.A(G50gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(KEYINPUT91), .A2(G43gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n210), .A2(G43gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT90), .B(KEYINPUT15), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OR3_X1    g016(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT15), .B1(new_n210), .B2(G43gat), .ZN(new_n221));
  INV_X1    g020(.A(G43gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(G50gat), .ZN(new_n223));
  INV_X1    g022(.A(G29gat), .ZN(new_n224));
  INV_X1    g023(.A(G36gat), .ZN(new_n225));
  OAI22_X1  g024(.A1(new_n221), .A2(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n217), .A2(new_n220), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT92), .ZN(new_n229));
  INV_X1    g028(.A(new_n223), .ZN(new_n230));
  INV_X1    g029(.A(new_n221), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n220), .A2(KEYINPUT89), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT89), .ZN(new_n233));
  OAI22_X1  g032(.A1(new_n218), .A2(new_n233), .B1(new_n224), .B2(new_n225), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n230), .B(new_n231), .C1(new_n232), .C2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT92), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n217), .A2(new_n236), .A3(new_n227), .A4(new_n220), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n229), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  AND2_X1   g037(.A1(new_n238), .A2(KEYINPUT17), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(KEYINPUT17), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n208), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n208), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(new_n238), .ZN(new_n243));
  NAND2_X1  g042(.A1(G229gat), .A2(G233gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n241), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT18), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n208), .B(new_n238), .Z(new_n248));
  XNOR2_X1  g047(.A(new_n244), .B(KEYINPUT13), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n241), .A2(KEYINPUT18), .A3(new_n243), .A4(new_n244), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n247), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(KEYINPUT87), .B(KEYINPUT11), .Z(new_n254));
  XNOR2_X1  g053(.A(G113gat), .B(G141gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G169gat), .B(G197gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT88), .B(KEYINPUT12), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n253), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n247), .A2(new_n260), .A3(new_n251), .A4(new_n252), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n262), .A2(KEYINPUT94), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT94), .B1(new_n262), .B2(new_n263), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G57gat), .B(G64gat), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G71gat), .B(G78gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT21), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n208), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G183gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  AND2_X1   g074(.A1(G231gat), .A2(G233gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n275), .A2(new_n276), .ZN(new_n279));
  XOR2_X1   g078(.A(G127gat), .B(G155gat), .Z(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT20), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n278), .A2(new_n279), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n282), .B1(new_n278), .B2(new_n279), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n271), .A2(KEYINPUT21), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(G211gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n287), .B(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n286), .B(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n239), .A2(new_n240), .ZN(new_n292));
  XOR2_X1   g091(.A(G99gat), .B(G106gat), .Z(new_n293));
  NAND2_X1  g092(.A1(G99gat), .A2(G106gat), .ZN(new_n294));
  INV_X1    g093(.A(G85gat), .ZN(new_n295));
  INV_X1    g094(.A(G92gat), .ZN(new_n296));
  AOI22_X1  g095(.A1(KEYINPUT8), .A2(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(KEYINPUT98), .ZN(new_n298));
  NAND2_X1  g097(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n299), .A2(G85gat), .A3(G92gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n293), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT99), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT98), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n297), .B(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n301), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n300), .B(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n293), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n306), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n303), .A2(new_n304), .A3(new_n310), .ZN(new_n311));
  OAI211_X1 g110(.A(KEYINPUT99), .B(new_n293), .C1(new_n298), .C2(new_n302), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n292), .A2(new_n313), .ZN(new_n314));
  AND3_X1   g113(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n313), .A2(new_n238), .ZN(new_n316));
  NOR3_X1   g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(G190gat), .B(G218gat), .Z(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT100), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n321), .B(KEYINPUT96), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n322), .B(G134gat), .ZN(new_n323));
  INV_X1    g122(.A(G162gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n317), .B(new_n318), .ZN(new_n327));
  XOR2_X1   g126(.A(new_n326), .B(new_n327), .Z(new_n328));
  NAND2_X1  g127(.A1(new_n291), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n271), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n311), .A2(new_n312), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n271), .A2(new_n303), .A3(new_n310), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G230gat), .A2(G233gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n334), .B(KEYINPUT103), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n313), .A2(KEYINPUT10), .A3(new_n271), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT10), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n331), .A2(new_n339), .A3(new_n332), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT101), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n331), .A2(KEYINPUT101), .A3(new_n339), .A4(new_n332), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n338), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n336), .B1(new_n344), .B2(new_n335), .ZN(new_n345));
  XNOR2_X1  g144(.A(G120gat), .B(G148gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(G176gat), .B(G204gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT102), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  AOI211_X1 g150(.A(KEYINPUT102), .B(new_n338), .C1(new_n342), .C2(new_n343), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n351), .A2(new_n352), .A3(new_n335), .ZN(new_n353));
  INV_X1    g152(.A(new_n348), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n354), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n353), .A2(KEYINPUT104), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT104), .ZN(new_n357));
  INV_X1    g156(.A(new_n344), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT102), .ZN(new_n359));
  INV_X1    g158(.A(new_n335), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n350), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n355), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n357), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n349), .B1(new_n356), .B2(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n329), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT31), .B(G50gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G197gat), .B(G204gat), .ZN(new_n369));
  INV_X1    g168(.A(G211gat), .ZN(new_n370));
  INV_X1    g169(.A(G218gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n369), .B1(KEYINPUT22), .B2(new_n372), .ZN(new_n373));
  XOR2_X1   g172(.A(G211gat), .B(G218gat), .Z(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT75), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n373), .B(new_n374), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n376), .B1(new_n378), .B2(KEYINPUT75), .ZN(new_n379));
  XOR2_X1   g178(.A(G155gat), .B(G162gat), .Z(new_n380));
  XNOR2_X1  g179(.A(G141gat), .B(G148gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT77), .B(KEYINPUT2), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT78), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(G141gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(G148gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT79), .B(G148gat), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n387), .B1(new_n388), .B2(new_n386), .ZN(new_n389));
  NAND2_X1  g188(.A1(G155gat), .A2(G162gat), .ZN(new_n390));
  INV_X1    g189(.A(G155gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n324), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n390), .B1(new_n392), .B2(KEYINPUT2), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n385), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT3), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT29), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n379), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OR2_X1    g198(.A1(new_n399), .A2(KEYINPUT81), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n396), .B1(new_n378), .B2(KEYINPUT29), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n394), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n401), .A2(new_n402), .B1(G228gat), .B2(G233gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(KEYINPUT81), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n400), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n379), .A2(new_n398), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n395), .B1(new_n406), .B2(new_n396), .ZN(new_n407));
  OAI211_X1 g206(.A(G228gat), .B(G233gat), .C1(new_n407), .C2(new_n399), .ZN(new_n408));
  XNOR2_X1  g207(.A(G78gat), .B(G106gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(G22gat), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n405), .A2(new_n408), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n411), .B1(new_n405), .B2(new_n408), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n368), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n414), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n416), .A2(new_n367), .A3(new_n412), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT85), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT71), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n422));
  NOR2_X1   g221(.A1(G169gat), .A2(G176gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT23), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n424), .B(KEYINPUT66), .Z(new_n425));
  NAND2_X1  g224(.A1(G169gat), .A2(G176gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT23), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n427), .B1(G169gat), .B2(G176gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n430));
  OAI221_X1 g229(.A(new_n429), .B1(G183gat), .B2(G190gat), .C1(new_n430), .C2(KEYINPUT65), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n430), .A2(KEYINPUT65), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n428), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n422), .B1(new_n425), .B2(new_n433), .ZN(new_n434));
  OR2_X1    g233(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(G190gat), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n430), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n429), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n440), .A2(KEYINPUT25), .A3(new_n428), .A4(new_n424), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n434), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n443));
  AND2_X1   g242(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n444));
  NOR2_X1   g243(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n443), .B1(new_n446), .B2(KEYINPUT27), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT68), .B1(new_n447), .B2(G190gat), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT28), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n435), .A2(KEYINPUT27), .A3(new_n436), .ZN(new_n450));
  INV_X1    g249(.A(new_n443), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT68), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(new_n453), .A3(new_n438), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n448), .A2(new_n449), .A3(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(KEYINPUT27), .B(G183gat), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n456), .A2(KEYINPUT28), .A3(new_n438), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(G183gat), .A2(G190gat), .ZN(new_n459));
  INV_X1    g258(.A(G169gat), .ZN(new_n460));
  INV_X1    g259(.A(G176gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT26), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT26), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n426), .A2(new_n463), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n459), .B(new_n462), .C1(new_n464), .C2(new_n423), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(KEYINPUT69), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT70), .B1(new_n458), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT70), .ZN(new_n469));
  AOI211_X1 g268(.A(new_n469), .B(new_n466), .C1(new_n455), .C2(new_n457), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n442), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G113gat), .B(G120gat), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n472), .A2(KEYINPUT1), .ZN(new_n473));
  XOR2_X1   g272(.A(G127gat), .B(G134gat), .Z(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n475), .B(new_n442), .C1(new_n468), .C2(new_n470), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(G227gat), .A2(G233gat), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n421), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  AOI211_X1 g281(.A(KEYINPUT71), .B(new_n480), .C1(new_n477), .C2(new_n478), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT32), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  XOR2_X1   g283(.A(KEYINPUT72), .B(KEYINPUT33), .Z(new_n485));
  OAI21_X1  g284(.A(new_n485), .B1(new_n482), .B2(new_n483), .ZN(new_n486));
  XNOR2_X1  g285(.A(G15gat), .B(G43gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(G71gat), .ZN(new_n488));
  INV_X1    g287(.A(G99gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n484), .A2(new_n486), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n477), .A2(new_n480), .A3(new_n478), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT34), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT73), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n493), .B1(new_n480), .B2(new_n494), .ZN(new_n495));
  XOR2_X1   g294(.A(new_n492), .B(new_n495), .Z(new_n496));
  INV_X1    g295(.A(new_n490), .ZN(new_n497));
  OAI221_X1 g296(.A(KEYINPUT32), .B1(new_n485), .B2(new_n497), .C1(new_n482), .C2(new_n483), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n491), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n496), .B1(new_n491), .B2(new_n498), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT74), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n491), .A2(new_n501), .A3(new_n496), .A4(new_n498), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n420), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n491), .A2(new_n498), .ZN(new_n506));
  INV_X1    g305(.A(new_n496), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n496), .A3(new_n498), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(KEYINPUT74), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n510), .A2(KEYINPUT85), .A3(new_n503), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n419), .B1(new_n505), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G226gat), .ZN(new_n513));
  INV_X1    g312(.A(G233gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n442), .B(new_n515), .C1(new_n468), .C2(new_n470), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n458), .A2(new_n467), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n442), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n515), .A2(KEYINPUT29), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n379), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT76), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(KEYINPUT76), .A3(new_n379), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n517), .A2(new_n442), .A3(new_n515), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n527), .B1(new_n471), .B2(new_n519), .ZN(new_n528));
  INV_X1    g327(.A(new_n379), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G8gat), .B(G36gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(G64gat), .B(G92gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n526), .A2(KEYINPUT30), .A3(new_n530), .A4(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT30), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n524), .A2(new_n530), .A3(new_n525), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n536), .B1(new_n537), .B2(new_n533), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n533), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(KEYINPUT80), .B(KEYINPUT0), .Z(new_n542));
  XNOR2_X1  g341(.A(G1gat), .B(G29gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G57gat), .B(G85gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT5), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n475), .B1(new_n402), .B2(KEYINPUT3), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n385), .A2(new_n394), .A3(new_n475), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT4), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT4), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n385), .A2(new_n552), .A3(new_n394), .A4(new_n475), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n397), .A2(new_n549), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G225gat), .A2(G233gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n402), .A2(new_n476), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n555), .B1(new_n557), .B2(new_n550), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n548), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT5), .B1(new_n554), .B2(new_n555), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n547), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT6), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n556), .A2(new_n548), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n558), .B1(new_n554), .B2(new_n555), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n564), .B(new_n546), .C1(new_n548), .C2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n562), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n560), .A2(new_n561), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(KEYINPUT6), .A3(new_n546), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NOR3_X1   g369(.A1(new_n541), .A2(KEYINPUT35), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(new_n569), .ZN(new_n572));
  AND4_X1   g371(.A1(new_n572), .A2(new_n535), .A3(new_n540), .A4(new_n538), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n573), .A2(new_n508), .A3(new_n418), .A4(new_n509), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT35), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT86), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n574), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n512), .A2(new_n571), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n379), .B1(new_n516), .B2(new_n520), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n580), .B1(new_n528), .B2(new_n379), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT38), .B1(new_n581), .B2(KEYINPUT37), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT82), .B(KEYINPUT37), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n524), .A2(new_n530), .A3(new_n525), .A4(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n582), .A2(new_n584), .A3(new_n533), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT83), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n537), .A2(new_n533), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n582), .A2(new_n584), .A3(KEYINPUT83), .A4(new_n533), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n587), .A2(new_n570), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT84), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n537), .A2(KEYINPUT37), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n584), .A2(new_n533), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT38), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n588), .B1(new_n585), .B2(new_n586), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n597), .A2(KEYINPUT84), .A3(new_n570), .A4(new_n590), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n593), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n554), .A2(new_n555), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n557), .A2(new_n555), .A3(new_n550), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(KEYINPUT39), .A3(new_n601), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n602), .B(new_n547), .C1(KEYINPUT39), .C2(new_n600), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT40), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n541), .A2(new_n566), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n599), .A2(new_n418), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT36), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n510), .A2(new_n607), .A3(new_n503), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n508), .A2(KEYINPUT36), .A3(new_n509), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n573), .A2(new_n418), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n606), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n266), .B(new_n366), .C1(new_n579), .C2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT105), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n266), .ZN(new_n617));
  AND3_X1   g416(.A1(new_n510), .A2(KEYINPUT85), .A3(new_n503), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT85), .B1(new_n510), .B2(new_n503), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n418), .B(new_n571), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n577), .A2(new_n578), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n617), .B1(new_n622), .B2(new_n612), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n623), .A2(KEYINPUT105), .A3(new_n366), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n616), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n570), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(G1gat), .ZN(G1324gat));
  INV_X1    g426(.A(KEYINPUT106), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n541), .ZN(new_n629));
  XOR2_X1   g428(.A(KEYINPUT16), .B(G8gat), .Z(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n628), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(KEYINPUT42), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT42), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n628), .B(new_n634), .C1(new_n629), .C2(new_n631), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n629), .A2(G8gat), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n633), .A2(new_n635), .A3(new_n636), .ZN(G1325gat));
  NAND2_X1  g436(.A1(new_n505), .A2(new_n511), .ZN(new_n638));
  AOI21_X1  g437(.A(G15gat), .B1(new_n625), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n610), .A2(KEYINPUT107), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT107), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n608), .A2(new_n641), .A3(new_n609), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n643), .B1(new_n616), .B2(new_n624), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n639), .B1(G15gat), .B2(new_n644), .ZN(G1326gat));
  XNOR2_X1  g444(.A(KEYINPUT43), .B(G22gat), .ZN(new_n646));
  INV_X1    g445(.A(new_n624), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT105), .B1(new_n623), .B2(new_n366), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n419), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT108), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT108), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n625), .A2(new_n651), .A3(new_n419), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n646), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n651), .B1(new_n625), .B2(new_n419), .ZN(new_n654));
  AOI211_X1 g453(.A(KEYINPUT108), .B(new_n418), .C1(new_n616), .C2(new_n624), .ZN(new_n655));
  INV_X1    g454(.A(new_n646), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n653), .A2(new_n657), .ZN(G1327gat));
  INV_X1    g457(.A(new_n291), .ZN(new_n659));
  INV_X1    g458(.A(new_n365), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(new_n328), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n623), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n663), .A2(new_n224), .A3(new_n570), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT45), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n326), .B(new_n327), .ZN(new_n666));
  OAI211_X1 g465(.A(KEYINPUT44), .B(new_n666), .C1(new_n579), .C2(new_n613), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n262), .A2(new_n263), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n661), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n670), .B(KEYINPUT109), .Z(new_n671));
  AND3_X1   g470(.A1(new_n608), .A2(new_n641), .A3(new_n609), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n641), .B1(new_n608), .B2(new_n609), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n611), .B(new_n606), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n328), .B1(new_n674), .B2(new_n622), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n667), .B(new_n671), .C1(new_n675), .C2(KEYINPUT44), .ZN(new_n676));
  OAI21_X1  g475(.A(G29gat), .B1(new_n676), .B2(new_n572), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n665), .A2(new_n677), .ZN(G1328gat));
  NAND3_X1  g477(.A1(new_n663), .A2(new_n225), .A3(new_n541), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n679), .B(KEYINPUT46), .Z(new_n680));
  INV_X1    g479(.A(new_n541), .ZN(new_n681));
  OAI21_X1  g480(.A(G36gat), .B1(new_n676), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(G1329gat));
  NAND2_X1  g482(.A1(new_n209), .A2(new_n211), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(new_n676), .B2(new_n643), .ZN(new_n686));
  AND4_X1   g485(.A1(new_n638), .A2(new_n623), .A3(new_n684), .A4(new_n662), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT47), .B1(new_n689), .B2(KEYINPUT110), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n606), .A2(new_n611), .ZN(new_n692));
  AOI22_X1  g491(.A1(new_n643), .A2(new_n692), .B1(new_n621), .B2(new_n620), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n693), .B2(new_n328), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n672), .A2(new_n673), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n694), .A2(new_n695), .A3(new_n667), .A4(new_n671), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n687), .B1(new_n696), .B2(new_n685), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT110), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT47), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n690), .A2(new_n700), .ZN(G1330gat));
  OAI21_X1  g500(.A(G50gat), .B1(new_n676), .B2(new_n418), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT48), .B1(new_n702), .B2(KEYINPUT111), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n663), .A2(new_n210), .A3(new_n419), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n702), .B(new_n704), .C1(KEYINPUT111), .C2(KEYINPUT48), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(G1331gat));
  NOR2_X1   g507(.A1(new_n693), .A2(new_n668), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n329), .A2(new_n660), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n570), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g513(.A1(new_n711), .A2(new_n681), .ZN(new_n715));
  NOR2_X1   g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  AND2_X1   g515(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n718), .B1(new_n715), .B2(new_n716), .ZN(G1333gat));
  NAND3_X1  g518(.A1(new_n712), .A2(G71gat), .A3(new_n695), .ZN(new_n720));
  INV_X1    g519(.A(G71gat), .ZN(new_n721));
  INV_X1    g520(.A(new_n638), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n711), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT50), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT50), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n720), .A2(new_n726), .A3(new_n723), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(G1334gat));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n419), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g529(.A1(new_n291), .A2(new_n668), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n694), .A2(new_n365), .A3(new_n667), .A4(new_n731), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n732), .A2(new_n295), .A3(new_n572), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n675), .A2(new_n731), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT51), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n675), .A2(KEYINPUT51), .A3(new_n731), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n738), .A2(new_n570), .A3(new_n365), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n733), .B1(new_n295), .B2(new_n739), .ZN(G1336gat));
  NAND2_X1  g539(.A1(new_n674), .A2(new_n622), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT44), .B1(new_n741), .B2(new_n666), .ZN(new_n742));
  AOI211_X1 g541(.A(new_n691), .B(new_n328), .C1(new_n622), .C2(new_n612), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n744), .A2(new_n541), .A3(new_n365), .A4(new_n731), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G92gat), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n681), .A2(G92gat), .A3(new_n660), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT52), .B1(new_n738), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n736), .A2(new_n737), .B1(new_n750), .B2(new_n747), .ZN(new_n751));
  OR2_X1    g550(.A1(new_n747), .A2(new_n750), .ZN(new_n752));
  AOI22_X1  g551(.A1(new_n745), .A2(G92gat), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n749), .B1(new_n753), .B2(new_n754), .ZN(G1337gat));
  NOR3_X1   g554(.A1(new_n732), .A2(new_n489), .A3(new_n643), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n738), .A2(new_n638), .A3(new_n365), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n756), .B1(new_n489), .B2(new_n757), .ZN(G1338gat));
  OAI21_X1  g557(.A(G106gat), .B1(new_n732), .B2(new_n418), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n418), .A2(G106gat), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n675), .A2(KEYINPUT51), .A3(new_n731), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT51), .B1(new_n675), .B2(new_n731), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n365), .B(new_n760), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n765), .B1(new_n763), .B2(KEYINPUT113), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n759), .B(new_n763), .C1(KEYINPUT113), .C2(new_n765), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(G1339gat));
  INV_X1    g568(.A(new_n258), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n248), .A2(new_n250), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n244), .B1(new_n241), .B2(new_n243), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n263), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n365), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT104), .B1(new_n353), .B2(new_n355), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n362), .A2(new_n357), .A3(new_n363), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n344), .A2(KEYINPUT54), .A3(new_n335), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(new_n354), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT54), .B1(new_n358), .B2(new_n360), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n353), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n780), .B(KEYINPUT55), .C1(new_n353), .C2(new_n781), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n778), .A2(new_n784), .A3(new_n668), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n775), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n775), .A2(new_n786), .A3(KEYINPUT114), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(new_n328), .A3(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n778), .A2(new_n784), .A3(new_n774), .A4(new_n785), .ZN(new_n792));
  OR2_X1    g591(.A1(new_n792), .A2(new_n328), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n291), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n329), .A2(new_n668), .A3(new_n365), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(new_n419), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n541), .A2(new_n572), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(new_n638), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(G113gat), .B1(new_n799), .B2(new_n617), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n796), .A2(new_n572), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n419), .A2(new_n499), .A3(new_n500), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(new_n541), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n669), .A2(G113gat), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(KEYINPUT115), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n800), .B1(new_n805), .B2(new_n807), .ZN(G1340gat));
  OR3_X1    g607(.A1(new_n805), .A2(G120gat), .A3(new_n660), .ZN(new_n809));
  OAI21_X1  g608(.A(G120gat), .B1(new_n799), .B2(new_n660), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(G1341gat));
  AOI21_X1  g610(.A(G127gat), .B1(new_n804), .B2(new_n291), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n799), .A2(new_n659), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n812), .B1(G127gat), .B2(new_n813), .ZN(G1342gat));
  NAND2_X1  g613(.A1(new_n681), .A2(new_n666), .ZN(new_n815));
  XOR2_X1   g614(.A(new_n815), .B(KEYINPUT116), .Z(new_n816));
  NOR3_X1   g615(.A1(new_n803), .A2(G134gat), .A3(new_n816), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT56), .ZN(new_n818));
  OAI21_X1  g617(.A(G134gat), .B1(new_n799), .B2(new_n328), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(G1343gat));
  NAND4_X1  g619(.A1(new_n266), .A2(new_n778), .A3(new_n784), .A4(new_n785), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n666), .B1(new_n821), .B2(new_n775), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n328), .A2(new_n792), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n659), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n795), .ZN(new_n827));
  OAI211_X1 g626(.A(KEYINPUT117), .B(new_n659), .C1(new_n822), .C2(new_n823), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n418), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT118), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n830), .B1(new_n796), .B2(new_n418), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n829), .A2(KEYINPUT118), .A3(new_n831), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n643), .A2(new_n798), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(new_n668), .A3(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n840), .B1(new_n796), .B2(new_n572), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n695), .A2(new_n418), .ZN(new_n842));
  OAI211_X1 g641(.A(KEYINPUT119), .B(new_n570), .C1(new_n794), .C2(new_n795), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n841), .A2(new_n681), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(G141gat), .ZN(new_n845));
  AOI22_X1  g644(.A1(G141gat), .A2(new_n839), .B1(new_n845), .B2(new_n266), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n848), .A2(new_n386), .A3(new_n681), .A4(new_n266), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n847), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851));
  INV_X1    g650(.A(new_n831), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n795), .B1(new_n824), .B2(new_n825), .ZN(new_n853));
  AOI211_X1 g652(.A(new_n851), .B(new_n852), .C1(new_n853), .C2(new_n828), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(new_n832), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n837), .B1(new_n855), .B2(new_n834), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n386), .B1(new_n856), .B2(new_n266), .ZN(new_n857));
  OAI22_X1  g656(.A1(new_n846), .A2(new_n847), .B1(new_n850), .B2(new_n857), .ZN(G1344gat));
  OR3_X1    g657(.A1(new_n844), .A2(new_n388), .A3(new_n660), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860));
  INV_X1    g659(.A(G148gat), .ZN(new_n861));
  OAI211_X1 g660(.A(KEYINPUT57), .B(new_n419), .C1(new_n794), .C2(new_n795), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n821), .A2(new_n775), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n793), .B1(new_n863), .B2(new_n666), .ZN(new_n864));
  AOI22_X1  g663(.A1(new_n864), .A2(new_n659), .B1(new_n617), .B2(new_n366), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n830), .B1(new_n865), .B2(new_n418), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n660), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n837), .A2(KEYINPUT120), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n837), .A2(KEYINPUT120), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n861), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n867), .A2(KEYINPUT121), .A3(new_n868), .A4(new_n869), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n860), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n836), .A2(new_n365), .A3(new_n838), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n875), .A2(new_n860), .A3(new_n388), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n859), .B1(new_n874), .B2(new_n876), .ZN(G1345gat));
  NAND3_X1  g676(.A1(new_n856), .A2(G155gat), .A3(new_n291), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n391), .B1(new_n844), .B2(new_n659), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(G1346gat));
  AOI21_X1  g679(.A(new_n324), .B1(new_n856), .B2(new_n666), .ZN(new_n881));
  INV_X1    g680(.A(new_n816), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n848), .A2(new_n324), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT122), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n836), .A2(new_n666), .A3(new_n838), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(G162gat), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n848), .A2(new_n324), .A3(new_n882), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n884), .A2(new_n889), .ZN(G1347gat));
  AND2_X1   g689(.A1(new_n791), .A2(new_n793), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n827), .B1(new_n891), .B2(new_n291), .ZN(new_n892));
  AND4_X1   g691(.A1(new_n572), .A2(new_n892), .A3(new_n541), .A4(new_n802), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(new_n460), .A3(new_n668), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT123), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n681), .A2(new_n570), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n638), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n797), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n895), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n898), .A2(new_n617), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n894), .B1(new_n901), .B2(new_n460), .ZN(G1348gat));
  NOR2_X1   g701(.A1(new_n898), .A2(new_n900), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(G176gat), .A3(new_n365), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT124), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n893), .A2(new_n365), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n461), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n903), .A2(new_n908), .A3(G176gat), .A4(new_n365), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n905), .A2(new_n907), .A3(new_n909), .ZN(G1349gat));
  NAND3_X1  g709(.A1(new_n893), .A2(new_n456), .A3(new_n291), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n898), .A2(new_n659), .A3(new_n900), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n912), .B2(new_n437), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT60), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT60), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n911), .B(new_n915), .C1(new_n912), .C2(new_n437), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1350gat));
  NAND3_X1  g716(.A1(new_n893), .A2(new_n438), .A3(new_n666), .ZN(new_n918));
  AOI211_X1 g717(.A(KEYINPUT61), .B(new_n438), .C1(new_n903), .C2(new_n666), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n920));
  INV_X1    g719(.A(new_n898), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n666), .A3(new_n899), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n920), .B1(new_n922), .B2(G190gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n918), .B1(new_n919), .B2(new_n923), .ZN(G1351gat));
  NAND2_X1  g723(.A1(new_n862), .A2(new_n866), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n643), .A2(new_n896), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G197gat), .B1(new_n928), .B2(new_n617), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n892), .A2(new_n572), .A3(new_n541), .A4(new_n842), .ZN(new_n930));
  OR3_X1    g729(.A1(new_n930), .A2(G197gat), .A3(new_n669), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(G1352gat));
  OR3_X1    g734(.A1(new_n930), .A2(G204gat), .A3(new_n660), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n936), .A2(KEYINPUT62), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n867), .A2(new_n927), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(G204gat), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n936), .A2(KEYINPUT62), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(G1353gat));
  AOI211_X1 g740(.A(new_n659), .B(new_n926), .C1(new_n862), .C2(new_n866), .ZN(new_n942));
  OAI21_X1  g741(.A(KEYINPUT63), .B1(new_n942), .B2(new_n370), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n659), .A2(G211gat), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n944), .B1(new_n930), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n643), .A2(new_n419), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n796), .A2(new_n948), .A3(new_n570), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n949), .A2(KEYINPUT126), .A3(new_n541), .A4(new_n945), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT63), .ZN(new_n952));
  OAI211_X1 g751(.A(new_n952), .B(G211gat), .C1(new_n928), .C2(new_n659), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n943), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT127), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n943), .A2(new_n951), .A3(new_n953), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(G1354gat));
  NOR3_X1   g757(.A1(new_n928), .A2(new_n371), .A3(new_n328), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n949), .A2(new_n541), .A3(new_n666), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n959), .B1(new_n371), .B2(new_n960), .ZN(G1355gat));
endmodule


