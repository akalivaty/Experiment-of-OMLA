//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n772, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n187));
  INV_X1    g001(.A(G131), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT65), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G137), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(KEYINPUT65), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n189), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n189), .A2(new_n192), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n188), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT11), .A2(G134), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n199), .B1(new_n191), .B2(new_n193), .ZN(new_n200));
  NOR2_X1   g014(.A1(KEYINPUT11), .A2(G134), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n201), .B1(G137), .B2(new_n198), .ZN(new_n202));
  AOI21_X1  g016(.A(G131), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n187), .B1(new_n197), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G146), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n208));
  OAI21_X1  g022(.A(G143), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n207), .A2(G143), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n209), .A2(G128), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  AND2_X1   g028(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n215));
  NOR2_X1   g029(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n214), .B1(new_n209), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G143), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(G146), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT64), .B(G146), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(new_n219), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n213), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n192), .A2(KEYINPUT65), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n190), .A2(G137), .ZN(new_n225));
  AOI21_X1  g039(.A(G134), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(G131), .B1(new_n226), .B2(new_n195), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n198), .B1(new_n224), .B2(new_n225), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n198), .A2(G137), .ZN(new_n229));
  OR2_X1    g043(.A1(KEYINPUT11), .A2(G134), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n188), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n227), .A2(new_n232), .A3(KEYINPUT71), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n204), .A2(new_n223), .A3(new_n233), .ZN(new_n234));
  AND2_X1   g048(.A1(KEYINPUT70), .A2(G119), .ZN(new_n235));
  NOR2_X1   g049(.A1(KEYINPUT70), .A2(G119), .ZN(new_n236));
  OAI21_X1  g050(.A(G116), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G119), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n237), .B1(G116), .B2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT2), .B(G113), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n240), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n242), .B(new_n237), .C1(G116), .C2(new_n238), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n209), .A2(KEYINPUT0), .A3(G128), .A4(new_n211), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT0), .B(G128), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n188), .A2(KEYINPUT66), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(new_n200), .B2(new_n202), .ZN(new_n250));
  NOR3_X1   g064(.A1(new_n228), .A2(new_n231), .A3(new_n248), .ZN(new_n251));
  OAI221_X1 g065(.A(new_n246), .B1(new_n222), .B2(new_n247), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n234), .A2(new_n245), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n227), .A2(new_n232), .A3(KEYINPUT67), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n217), .B1(new_n221), .B2(new_n219), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n222), .B1(G128), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n205), .A2(G146), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n219), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NOR4_X1   g074(.A1(new_n260), .A2(new_n217), .A3(new_n214), .A4(new_n210), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n255), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT67), .B1(new_n227), .B2(new_n232), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n252), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT30), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n264), .A2(KEYINPUT69), .A3(new_n265), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n233), .B1(new_n257), .B2(new_n261), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT71), .B1(new_n227), .B2(new_n232), .ZN(new_n271));
  OAI211_X1 g085(.A(KEYINPUT30), .B(new_n252), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n234), .A2(KEYINPUT72), .A3(KEYINPUT30), .A4(new_n252), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n268), .A2(new_n269), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n254), .B1(new_n276), .B2(new_n244), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n278), .B(G101), .ZN(new_n279));
  NOR2_X1   g093(.A1(G237), .A2(G953), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G210), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n279), .B(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n263), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(new_n223), .A3(new_n255), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n245), .B1(new_n286), .B2(new_n252), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT28), .B1(new_n254), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT74), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n234), .A2(new_n289), .A3(new_n252), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n289), .B1(new_n234), .B2(new_n252), .ZN(new_n291));
  NOR3_X1   g105(.A1(new_n290), .A2(new_n291), .A3(new_n244), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n288), .B1(new_n292), .B2(KEYINPUT28), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n282), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT29), .B1(new_n284), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G902), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n234), .A2(new_n252), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT74), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n234), .A2(new_n289), .A3(new_n252), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n245), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT28), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n297), .A2(new_n244), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n253), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT28), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n282), .A2(KEYINPUT29), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n296), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G472), .B1(new_n295), .B2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(G472), .A2(G902), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n253), .A2(KEYINPUT73), .A3(new_n282), .ZN(new_n312));
  AOI21_X1  g126(.A(KEYINPUT31), .B1(new_n276), .B2(new_n244), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n274), .A2(new_n275), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT69), .B1(new_n264), .B2(new_n265), .ZN(new_n315));
  AOI211_X1 g129(.A(new_n267), .B(KEYINPUT30), .C1(new_n286), .C2(new_n252), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n314), .B(new_n244), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n312), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n312), .A2(new_n313), .B1(new_n318), .B2(KEYINPUT31), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT75), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n264), .A2(new_n244), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n301), .B1(new_n321), .B2(new_n253), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n322), .B1(new_n301), .B2(new_n300), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n320), .B1(new_n323), .B2(new_n282), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n293), .A2(KEYINPUT75), .A3(new_n283), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AOI211_X1 g140(.A(KEYINPUT32), .B(new_n311), .C1(new_n319), .C2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT32), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n318), .A2(KEYINPUT31), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT31), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n317), .A2(new_n330), .A3(new_n312), .ZN(new_n331));
  AOI211_X1 g145(.A(new_n320), .B(new_n282), .C1(new_n302), .C2(new_n288), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT75), .B1(new_n293), .B2(new_n283), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n329), .B(new_n331), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n328), .B1(new_n334), .B2(new_n310), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n309), .B1(new_n327), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(KEYINPUT76), .B(new_n309), .C1(new_n327), .C2(new_n335), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT94), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT16), .ZN(new_n341));
  INV_X1    g155(.A(G125), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n342), .A2(KEYINPUT78), .A3(G140), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G140), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G125), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(G140), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT78), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n341), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n346), .A2(KEYINPUT16), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n207), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n350), .ZN(new_n352));
  XNOR2_X1  g166(.A(G125), .B(G140), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n343), .B1(new_n353), .B2(KEYINPUT78), .ZN(new_n354));
  OAI211_X1 g168(.A(G146), .B(new_n352), .C1(new_n354), .C2(new_n341), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT17), .ZN(new_n357));
  INV_X1    g171(.A(G237), .ZN(new_n358));
  INV_X1    g172(.A(G953), .ZN(new_n359));
  AND4_X1   g173(.A1(G143), .A2(new_n358), .A3(new_n359), .A4(G214), .ZN(new_n360));
  AOI21_X1  g174(.A(G143), .B1(new_n280), .B2(G214), .ZN(new_n361));
  OAI21_X1  g175(.A(G131), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT93), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n358), .A2(new_n359), .A3(G214), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n219), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n280), .A2(G143), .A3(G214), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT93), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n368), .A3(G131), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n357), .B1(new_n363), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n340), .B1(new_n356), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n368), .B1(new_n367), .B2(G131), .ZN(new_n372));
  AOI211_X1 g186(.A(KEYINPUT93), .B(new_n188), .C1(new_n365), .C2(new_n366), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT17), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n374), .A2(KEYINPUT94), .A3(new_n355), .A4(new_n351), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n367), .A2(G131), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n372), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n357), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n371), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G113), .B(G122), .ZN(new_n380));
  INV_X1    g194(.A(G104), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n380), .B(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(KEYINPUT18), .A2(G131), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n367), .B(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n353), .B1(new_n206), .B2(new_n208), .ZN(new_n385));
  INV_X1    g199(.A(new_n354), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n385), .B1(new_n386), .B2(new_n207), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n379), .A2(new_n382), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n382), .B1(new_n379), .B2(new_n388), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n296), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT96), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI211_X1 g207(.A(KEYINPUT96), .B(new_n296), .C1(new_n389), .C2(new_n390), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(G475), .A3(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(G475), .A2(G902), .ZN(new_n396));
  XOR2_X1   g210(.A(new_n396), .B(KEYINPUT95), .Z(new_n397));
  NAND3_X1  g211(.A1(new_n379), .A2(new_n382), .A3(new_n388), .ZN(new_n398));
  MUX2_X1   g212(.A(new_n353), .B(new_n354), .S(KEYINPUT19), .Z(new_n399));
  OAI21_X1  g213(.A(new_n355), .B1(new_n399), .B2(new_n221), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n388), .B1(new_n400), .B2(new_n377), .ZN(new_n401));
  INV_X1    g215(.A(new_n382), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n397), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT20), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n404), .B(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n395), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT99), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT14), .ZN(new_n409));
  INV_X1    g223(.A(G116), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n409), .B1(new_n410), .B2(G122), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n410), .A2(G122), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G122), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G116), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n414), .A2(G116), .ZN(new_n416));
  OAI211_X1 g230(.A(KEYINPUT99), .B(new_n415), .C1(new_n416), .C2(new_n409), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(KEYINPUT100), .A3(new_n409), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT100), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n410), .A2(G122), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n419), .B1(new_n420), .B2(KEYINPUT14), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n413), .A2(new_n417), .A3(new_n418), .A4(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G107), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT97), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n424), .B1(new_n415), .B2(new_n420), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n415), .A2(new_n420), .A3(new_n424), .ZN(new_n427));
  AOI21_X1  g241(.A(G107), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n214), .A2(G143), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n219), .A2(G128), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(new_n189), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n423), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n189), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT13), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n436), .B1(new_n214), .B2(G143), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT98), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n431), .A2(KEYINPUT98), .A3(new_n436), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n219), .A2(KEYINPUT13), .A3(G128), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n439), .A2(new_n440), .A3(new_n430), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G134), .ZN(new_n443));
  INV_X1    g257(.A(new_n427), .ZN(new_n444));
  INV_X1    g258(.A(G107), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n444), .A2(new_n445), .A3(new_n425), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n435), .B(new_n443), .C1(new_n428), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n434), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT9), .B(G234), .ZN(new_n449));
  INV_X1    g263(.A(G217), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n449), .A2(new_n450), .A3(G953), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT101), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n434), .A2(new_n447), .A3(new_n451), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n448), .A2(KEYINPUT101), .A3(new_n452), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT102), .ZN(new_n459));
  INV_X1    g273(.A(G478), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(KEYINPUT15), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n458), .A2(new_n459), .A3(new_n296), .A4(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n456), .A2(new_n296), .A3(new_n457), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n461), .B1(new_n464), .B2(KEYINPUT102), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n464), .A2(KEYINPUT102), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n407), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(G234), .A2(G237), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(G952), .A3(new_n359), .ZN(new_n470));
  XOR2_X1   g284(.A(KEYINPUT21), .B(G898), .Z(new_n471));
  NAND3_X1  g285(.A1(new_n469), .A2(G902), .A3(G953), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT0), .ZN(new_n475));
  NOR4_X1   g289(.A1(new_n260), .A2(new_n475), .A3(new_n214), .A4(new_n210), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n221), .A2(new_n219), .ZN(new_n477));
  INV_X1    g291(.A(new_n220), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n247), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(G125), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n342), .B(new_n213), .C1(new_n218), .C2(new_n222), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT88), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n359), .A2(G224), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT88), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n483), .A2(KEYINPUT7), .A3(new_n484), .A4(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(G110), .B(G122), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT8), .ZN(new_n489));
  XOR2_X1   g303(.A(KEYINPUT85), .B(KEYINPUT5), .Z(new_n490));
  OR2_X1    g304(.A1(KEYINPUT70), .A2(G119), .ZN(new_n491));
  NAND2_X1  g305(.A1(KEYINPUT70), .A2(G119), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n490), .A2(G116), .A3(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n494), .B(G113), .C1(new_n239), .C2(new_n490), .ZN(new_n495));
  INV_X1    g309(.A(G101), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n445), .A2(G104), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n381), .A2(G107), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT3), .B1(new_n381), .B2(G107), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT83), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n445), .B2(G104), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT3), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(new_n445), .A3(G104), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n381), .A2(KEYINPUT83), .A3(G107), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n501), .A2(new_n503), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n500), .B1(new_n507), .B2(G101), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n495), .A2(new_n243), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n243), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n494), .A2(G113), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n237), .B(KEYINPUT5), .C1(G116), .C2(new_n238), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n489), .B(new_n509), .C1(new_n513), .C2(new_n508), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n487), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT90), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n359), .A2(G224), .B1(KEYINPUT89), .B2(KEYINPUT7), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n517), .B1(KEYINPUT89), .B2(KEYINPUT7), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n482), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n516), .B1(new_n482), .B2(new_n518), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT91), .B1(new_n515), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n521), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n519), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT91), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n525), .A2(new_n526), .A3(new_n487), .A4(new_n514), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n503), .A2(new_n506), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n528), .A2(new_n496), .A3(new_n501), .A4(new_n505), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n507), .A2(G101), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(KEYINPUT4), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT4), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n507), .A2(new_n532), .A3(G101), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(new_n244), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n507), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n499), .B1(new_n535), .B2(new_n496), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n495), .A2(new_n536), .A3(new_n243), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n534), .A2(new_n488), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n523), .A2(new_n527), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n483), .A2(new_n486), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(G224), .A3(new_n359), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n488), .B1(new_n534), .B2(new_n537), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT6), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT87), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT87), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n545), .A2(new_n549), .A3(new_n546), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT86), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n538), .A2(new_n545), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n552), .B1(new_n553), .B2(KEYINPUT6), .ZN(new_n554));
  NOR4_X1   g368(.A1(new_n538), .A2(new_n545), .A3(KEYINPUT86), .A4(new_n546), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n544), .B(new_n551), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n540), .A2(new_n556), .A3(new_n296), .ZN(new_n557));
  OAI21_X1  g371(.A(G210), .B1(G237), .B2(G902), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT92), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n540), .A2(new_n556), .A3(new_n296), .A4(new_n560), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(G214), .B1(G237), .B2(G902), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G221), .B1(new_n449), .B2(G902), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G469), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n250), .A2(new_n251), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(G128), .B1(new_n260), .B2(new_n212), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n477), .A2(new_n478), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n574), .A2(new_n213), .A3(new_n508), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT1), .ZN(new_n576));
  OAI21_X1  g390(.A(G128), .B1(new_n220), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n260), .B2(new_n210), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n508), .B1(new_n213), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n571), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT12), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT12), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n582), .B(new_n571), .C1(new_n575), .C2(new_n579), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT10), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n213), .A2(new_n578), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n584), .B1(new_n585), .B2(new_n508), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n476), .A2(new_n479), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(new_n531), .A3(new_n533), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n223), .A2(KEYINPUT10), .A3(new_n536), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n586), .A2(new_n588), .A3(new_n589), .A4(new_n570), .ZN(new_n590));
  XNOR2_X1  g404(.A(G110), .B(G140), .ZN(new_n591));
  INV_X1    g405(.A(G227), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(G953), .ZN(new_n593));
  XOR2_X1   g407(.A(new_n591), .B(new_n593), .Z(new_n594));
  NAND4_X1  g408(.A1(new_n581), .A2(new_n583), .A3(new_n590), .A4(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n571), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n594), .B1(new_n598), .B2(new_n590), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n569), .B(new_n296), .C1(new_n596), .C2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT84), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n598), .A2(new_n590), .ZN(new_n603));
  INV_X1    g417(.A(new_n594), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n595), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n606), .A2(KEYINPUT84), .A3(new_n569), .A4(new_n296), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n581), .A2(new_n590), .A3(new_n583), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n604), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n598), .A2(new_n590), .A3(new_n594), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n296), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(G469), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n568), .B1(new_n608), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n474), .A2(new_n566), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT23), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n618), .B1(new_n493), .B2(G128), .ZN(new_n619));
  INV_X1    g433(.A(G110), .ZN(new_n620));
  OAI21_X1  g434(.A(G128), .B1(new_n235), .B2(new_n236), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n214), .A2(KEYINPUT23), .A3(G119), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n619), .A2(new_n620), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT24), .B(G110), .Z(new_n625));
  INV_X1    g439(.A(KEYINPUT77), .ZN(new_n626));
  AOI22_X1  g440(.A1(new_n621), .A2(new_n626), .B1(G119), .B2(new_n214), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n493), .A2(KEYINPUT77), .A3(G128), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n355), .B(new_n385), .C1(new_n624), .C2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(KEYINPUT79), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n627), .A2(new_n628), .ZN(new_n632));
  INV_X1    g446(.A(new_n625), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n623), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT79), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n635), .A2(new_n636), .A3(new_n355), .A4(new_n385), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n627), .A2(new_n625), .A3(new_n628), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n619), .A2(new_n621), .A3(new_n622), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n356), .B(new_n638), .C1(new_n620), .C2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n631), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n359), .A2(G221), .A3(G234), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT22), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G137), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n631), .A2(new_n637), .A3(new_n640), .A4(new_n644), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n646), .A2(new_n296), .A3(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT25), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT80), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n646), .A2(new_n647), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT81), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n653), .A2(new_n654), .A3(KEYINPUT25), .A4(new_n296), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT81), .B1(new_n648), .B2(new_n649), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n648), .A2(KEYINPUT80), .A3(new_n649), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n652), .A2(new_n655), .A3(new_n656), .A4(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n450), .B1(G234), .B2(new_n296), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n659), .A2(G902), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n653), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT82), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n338), .A2(new_n339), .A3(new_n617), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G101), .ZN(G3));
  NAND2_X1  g481(.A1(new_n334), .A2(new_n310), .ZN(new_n668));
  AOI21_X1  g482(.A(G902), .B1(new_n319), .B2(new_n326), .ZN(new_n669));
  INV_X1    g483(.A(G472), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n671), .A2(new_n664), .A3(new_n616), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n557), .A2(new_n558), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n540), .A2(new_n556), .A3(new_n296), .A4(new_n559), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n673), .A2(new_n565), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT33), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n456), .A2(new_n676), .A3(new_n457), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n453), .A2(KEYINPUT33), .A3(new_n455), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n679), .A2(KEYINPUT103), .A3(G478), .A4(new_n296), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n464), .A2(new_n460), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n677), .A2(G478), .A3(new_n296), .A4(new_n678), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT103), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n680), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n407), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n675), .A2(new_n686), .A3(new_n473), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n672), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT34), .B(G104), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G6));
  XOR2_X1   g505(.A(new_n473), .B(KEYINPUT104), .Z(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n395), .A2(new_n406), .A3(new_n467), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n675), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n672), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT35), .B(G107), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G9));
  AOI21_X1  g513(.A(new_n670), .B1(new_n334), .B2(new_n296), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n310), .B2(new_n334), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n645), .A2(KEYINPUT36), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n641), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n661), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n660), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n617), .A2(new_n701), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT37), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n620), .ZN(G12));
  NAND4_X1  g522(.A1(new_n615), .A2(new_n565), .A3(new_n673), .A4(new_n674), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n470), .B1(new_n472), .B2(G900), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n395), .A2(new_n406), .A3(new_n467), .A4(new_n710), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n711), .A2(KEYINPUT105), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(KEYINPUT105), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n709), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n338), .A2(new_n714), .A3(new_n339), .A4(new_n705), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G128), .ZN(G30));
  XOR2_X1   g530(.A(new_n710), .B(KEYINPUT39), .Z(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n615), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(KEYINPUT107), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(KEYINPUT40), .ZN(new_n721));
  AOI22_X1  g535(.A1(new_n658), .A2(new_n659), .B1(new_n661), .B2(new_n703), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n407), .A2(new_n467), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n277), .A2(new_n283), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n296), .B1(new_n304), .B2(new_n282), .ZN(new_n726));
  OAI21_X1  g540(.A(G472), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(new_n727), .B(KEYINPUT106), .Z(new_n728));
  NAND2_X1  g542(.A1(new_n668), .A2(KEYINPUT32), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n334), .A2(new_n328), .A3(new_n310), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n564), .B(KEYINPUT38), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n732), .A2(new_n565), .A3(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n721), .A2(new_n722), .A3(new_n724), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G143), .ZN(G45));
  AOI21_X1  g550(.A(KEYINPUT76), .B1(new_n731), .B2(new_n309), .ZN(new_n737));
  INV_X1    g551(.A(new_n339), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n709), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n407), .A2(new_n685), .A3(new_n710), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n739), .A2(new_n705), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G146), .ZN(G48));
  INV_X1    g557(.A(new_n606), .ZN(new_n744));
  OAI21_X1  g558(.A(G469), .B1(new_n744), .B2(G902), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n608), .A2(new_n567), .A3(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n338), .A2(new_n339), .A3(new_n665), .A4(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n687), .ZN(new_n749));
  XOR2_X1   g563(.A(KEYINPUT41), .B(G113), .Z(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G15));
  NOR2_X1   g565(.A1(new_n748), .A2(new_n695), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n410), .ZN(G18));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n675), .A2(new_n747), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n673), .A2(new_n565), .A3(new_n674), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT108), .B1(new_n756), .B2(new_n746), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n474), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n758), .A2(new_n338), .A3(new_n339), .A4(new_n705), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G119), .ZN(G21));
  NAND2_X1  g574(.A1(new_n306), .A2(new_n283), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n311), .B1(new_n319), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n700), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n665), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n756), .A2(new_n723), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n747), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n764), .A2(new_n766), .A3(new_n692), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(new_n414), .ZN(G24));
  NAND2_X1  g582(.A1(new_n755), .A2(new_n757), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n700), .A2(new_n722), .A3(new_n762), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n741), .A3(new_n770), .ZN(new_n771));
  XOR2_X1   g585(.A(KEYINPUT109), .B(G125), .Z(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(G27));
  INV_X1    g587(.A(KEYINPUT42), .ZN(new_n774));
  INV_X1    g588(.A(new_n565), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n568), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n562), .A2(new_n563), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT110), .B1(new_n610), .B2(new_n611), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n611), .A2(KEYINPUT110), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n296), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AOI22_X1  g594(.A1(new_n780), .A2(G469), .B1(new_n602), .B2(new_n607), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n338), .A2(new_n339), .A3(new_n665), .A4(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n407), .A2(new_n685), .A3(new_n710), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n774), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n664), .B1(new_n731), .B2(new_n309), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n784), .A2(new_n777), .A3(new_n781), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n786), .A2(KEYINPUT42), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G131), .ZN(G33));
  AND4_X1   g604(.A1(new_n338), .A2(new_n339), .A3(new_n665), .A4(new_n782), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n712), .A2(new_n713), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G134), .ZN(G36));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n795));
  OR3_X1    g609(.A1(new_n778), .A2(new_n795), .A3(new_n779), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n612), .A2(new_n795), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(G469), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(G469), .A2(G902), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT46), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT111), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n800), .A2(KEYINPUT46), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n800), .A2(new_n804), .A3(KEYINPUT46), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n802), .A2(new_n803), .A3(new_n608), .A4(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n567), .A3(new_n718), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT112), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n671), .A2(new_n705), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT113), .ZN(new_n810));
  INV_X1    g624(.A(new_n685), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n407), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n812), .A2(KEYINPUT43), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(KEYINPUT43), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT44), .B1(new_n810), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n564), .A2(new_n775), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n810), .A2(KEYINPUT44), .A3(new_n815), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n808), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G137), .ZN(G39));
  NAND2_X1  g636(.A1(new_n806), .A2(new_n567), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT47), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n823), .B(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n739), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n818), .A2(new_n665), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n825), .A2(new_n826), .A3(new_n741), .A4(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G140), .ZN(G42));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n830));
  INV_X1    g644(.A(new_n732), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n608), .A2(new_n745), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(KEYINPUT49), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n831), .A2(new_n776), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n664), .B1(new_n834), .B2(KEYINPUT49), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n839), .B1(new_n833), .B2(new_n835), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n733), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n838), .A2(new_n812), .A3(new_n841), .ZN(new_n842));
  AOI211_X1 g656(.A(new_n470), .B(new_n764), .C1(new_n813), .C2(new_n814), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n733), .A2(new_n565), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n843), .A2(new_n747), .A3(new_n844), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n845), .B(KEYINPUT50), .Z(new_n846));
  NOR2_X1   g660(.A1(new_n832), .A2(new_n567), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n817), .B(new_n843), .C1(new_n825), .C2(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n777), .A2(new_n470), .A3(new_n832), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n815), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n770), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n831), .A2(new_n665), .A3(new_n849), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(new_n395), .A3(new_n406), .A4(new_n811), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n846), .A2(new_n848), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT51), .B1(new_n848), .B2(new_n855), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n854), .A2(new_n856), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n850), .A2(new_n786), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT48), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n843), .A2(new_n769), .ZN(new_n862));
  INV_X1    g676(.A(G952), .ZN(new_n863));
  AOI211_X1 g677(.A(new_n863), .B(G953), .C1(new_n852), .C2(new_n686), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n338), .A2(new_n339), .A3(new_n705), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n817), .A2(new_n468), .A3(new_n710), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT115), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n817), .A2(KEYINPUT115), .A3(new_n468), .A4(new_n710), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n616), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n792), .A2(new_n791), .B1(new_n866), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n759), .B1(new_n748), .B2(new_n695), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n748), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n767), .B1(new_n875), .B2(new_n688), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n872), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT116), .ZN(new_n878));
  INV_X1    g692(.A(new_n762), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n705), .B(new_n879), .C1(new_n670), .C2(new_n669), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n562), .A2(new_n563), .A3(new_n776), .ZN(new_n881));
  INV_X1    g695(.A(new_n781), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n741), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n878), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n770), .A2(new_n787), .A3(KEYINPUT116), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n686), .A2(new_n694), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(new_n566), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n672), .A2(new_n888), .A3(new_n693), .ZN(new_n889));
  AND4_X1   g703(.A1(new_n666), .A2(new_n886), .A3(new_n706), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n789), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n877), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n338), .A2(new_n339), .A3(new_n705), .A4(new_n741), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n715), .B(new_n771), .C1(new_n893), .C2(new_n709), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n765), .A2(new_n567), .A3(new_n710), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n732), .A2(new_n895), .A3(new_n722), .A4(new_n882), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT52), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n715), .A2(new_n771), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT52), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n899), .A2(new_n742), .A3(new_n900), .A4(new_n896), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n892), .A2(new_n902), .A3(KEYINPUT53), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT53), .ZN(new_n904));
  INV_X1    g718(.A(new_n767), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n905), .B1(new_n748), .B2(new_n687), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n906), .A2(new_n873), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n907), .A2(new_n789), .A3(new_n890), .A4(new_n872), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n898), .A2(new_n901), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n904), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n903), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT54), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n903), .A2(new_n910), .A3(KEYINPUT54), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n865), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n859), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(G952), .A2(G953), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT118), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n830), .B(new_n842), .C1(new_n916), .C2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n919), .B1(new_n859), .B2(new_n915), .ZN(new_n921));
  INV_X1    g735(.A(new_n842), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT119), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n920), .A2(new_n923), .ZN(G75));
  AOI21_X1  g738(.A(new_n296), .B1(new_n903), .B2(new_n910), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT56), .B1(new_n925), .B2(G210), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n551), .B1(new_n554), .B2(new_n555), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(new_n544), .Z(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT55), .ZN(new_n929));
  NOR2_X1   g743(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n926), .B(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n863), .A2(G953), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT121), .Z(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n932), .A2(new_n935), .ZN(G51));
  AND3_X1   g750(.A1(new_n903), .A2(KEYINPUT54), .A3(new_n910), .ZN(new_n937));
  AOI21_X1  g751(.A(KEYINPUT54), .B1(new_n903), .B2(new_n910), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n799), .B(KEYINPUT57), .Z(new_n940));
  AOI21_X1  g754(.A(new_n744), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n798), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n911), .A2(G902), .A3(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT122), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n925), .A2(KEYINPUT122), .A3(new_n942), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n934), .B1(new_n941), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT123), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g764(.A(KEYINPUT123), .B(new_n934), .C1(new_n941), .C2(new_n947), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(G54));
  NAND3_X1  g766(.A1(new_n925), .A2(KEYINPUT58), .A3(G475), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n398), .A2(new_n403), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n953), .B(new_n954), .Z(new_n955));
  NOR2_X1   g769(.A1(new_n955), .A2(new_n935), .ZN(G60));
  NAND2_X1  g770(.A1(G478), .A2(G902), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT59), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n939), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n679), .B(KEYINPUT124), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n959), .A2(new_n960), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n961), .A2(new_n962), .A3(new_n935), .ZN(G63));
  NAND2_X1  g777(.A1(G217), .A2(G902), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT60), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(new_n903), .B2(new_n910), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n935), .B1(new_n966), .B2(new_n703), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n653), .B2(new_n966), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g783(.A(new_n359), .B1(new_n471), .B2(G224), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n666), .A2(new_n889), .A3(new_n706), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n907), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n970), .B1(new_n972), .B2(new_n359), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n927), .B1(G898), .B2(new_n359), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n973), .B(new_n974), .Z(G69));
  XOR2_X1   g789(.A(new_n276), .B(new_n399), .Z(new_n976));
  NAND3_X1  g790(.A1(new_n592), .A2(G900), .A3(G953), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n808), .A2(new_n765), .A3(new_n786), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT125), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n821), .A2(new_n828), .A3(new_n789), .ZN(new_n980));
  INV_X1    g794(.A(new_n894), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n793), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n979), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n976), .B(new_n977), .C1(new_n984), .C2(G953), .ZN(new_n985));
  AND2_X1   g799(.A1(G227), .A2(G900), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n976), .B1(G953), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n735), .A2(new_n981), .ZN(new_n988));
  OR2_X1    g802(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n989), .A2(new_n821), .A3(new_n828), .A4(new_n990), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n739), .A2(new_n665), .A3(new_n720), .A4(new_n817), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n992), .A2(new_n887), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n359), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n987), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n985), .A2(new_n995), .ZN(G72));
  NAND2_X1  g810(.A1(G472), .A2(G902), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT63), .Z(new_n998));
  INV_X1    g812(.A(new_n972), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n993), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n998), .B1(new_n991), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n725), .ZN(new_n1002));
  INV_X1    g816(.A(new_n284), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n1003), .A2(new_n725), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n911), .A2(new_n998), .A3(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1002), .A2(new_n934), .A3(new_n1005), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n979), .A2(new_n999), .A3(new_n980), .A4(new_n983), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT126), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n1007), .A2(new_n1008), .A3(new_n998), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1008), .B1(new_n1007), .B2(new_n998), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n284), .B(KEYINPUT127), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1006), .B1(new_n1011), .B2(new_n1012), .ZN(G57));
endmodule


