//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1315,
    new_n1316, new_n1317, new_n1318, new_n1319, new_n1320, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT64), .Z(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n203), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n207), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n211), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT65), .Z(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n223), .A2(new_n224), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n211), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n202), .A2(new_n203), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n229), .B1(new_n232), .B2(new_n235), .ZN(new_n236));
  AND3_X1   g0036(.A1(new_n225), .A2(new_n226), .A3(new_n236), .ZN(G361));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT66), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G264), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n201), .A2(G68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n203), .A2(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n249), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  OAI21_X1  g0056(.A(KEYINPUT67), .B1(new_n211), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT67), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n258), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n257), .A2(new_n230), .A3(new_n259), .A4(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT68), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n231), .A2(G1), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n264), .B1(new_n265), .B2(new_n201), .ZN(new_n266));
  INV_X1    g0066(.A(new_n265), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(KEYINPUT68), .A3(G50), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n263), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n257), .A2(new_n230), .A3(new_n259), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT8), .B(G58), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n256), .A2(G20), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G150), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G20), .A2(G33), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  OAI22_X1  g0076(.A1(new_n271), .A2(new_n273), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n204), .A2(G20), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n270), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n269), .B(new_n279), .C1(G50), .C2(new_n261), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT9), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g0082(.A(new_n282), .B(KEYINPUT69), .Z(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n256), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(G222), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(G1698), .ZN(new_n290));
  INV_X1    g0090(.A(G223), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n289), .B1(new_n218), .B2(new_n287), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G41), .ZN(new_n295));
  INV_X1    g0095(.A(G45), .ZN(new_n296));
  AOI21_X1  g0096(.A(G1), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G33), .A2(G41), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n298), .A2(G1), .A3(G13), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n297), .A2(new_n299), .A3(G274), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n293), .A2(new_n297), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(G226), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n294), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G200), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  OAI221_X1 g0106(.A(new_n305), .B1(new_n281), .B2(new_n280), .C1(new_n306), .C2(new_n304), .ZN(new_n307));
  OR3_X1    g0107(.A1(new_n283), .A2(new_n307), .A3(KEYINPUT10), .ZN(new_n308));
  OAI21_X1  g0108(.A(KEYINPUT10), .B1(new_n283), .B2(new_n307), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n304), .ZN(new_n311));
  INV_X1    g0111(.A(G179), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n313), .B(new_n280), .C1(G169), .C2(new_n311), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n287), .A2(G232), .A3(new_n288), .ZN(new_n315));
  OAI221_X1 g0115(.A(new_n315), .B1(new_n207), .B2(new_n287), .C1(new_n290), .C2(new_n213), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n293), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n301), .B1(G244), .B2(new_n302), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n271), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n322), .A2(new_n275), .B1(G20), .B2(G77), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT15), .B(G87), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n273), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n261), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n325), .A2(new_n270), .B1(new_n218), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n263), .A2(G77), .A3(new_n267), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n321), .B(new_n329), .C1(G179), .C2(new_n319), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n319), .A2(G200), .ZN(new_n332));
  INV_X1    g0132(.A(new_n319), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n329), .B1(new_n333), .B2(G190), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n331), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n310), .A2(new_n314), .A3(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(KEYINPUT3), .A2(G33), .ZN(new_n337));
  NOR2_X1   g0137(.A1(KEYINPUT3), .A2(G33), .ZN(new_n338));
  OAI211_X1 g0138(.A(G226), .B(new_n288), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  OAI211_X1 g0139(.A(G232), .B(G1698), .C1(new_n337), .C2(new_n338), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G33), .A2(G97), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n293), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n299), .A2(G238), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT70), .ZN(new_n346));
  AND3_X1   g0146(.A1(new_n300), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n346), .B1(new_n300), .B2(new_n345), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n343), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT13), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT13), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n343), .B(new_n351), .C1(new_n347), .C2(new_n348), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n350), .A2(G179), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT71), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n350), .A2(new_n354), .A3(new_n352), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT73), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n349), .A2(KEYINPUT71), .A3(KEYINPUT13), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n355), .A2(new_n356), .A3(G169), .A4(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n353), .B1(new_n358), .B2(KEYINPUT14), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT72), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT14), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n355), .A2(G169), .A3(new_n357), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n362), .B1(new_n363), .B2(new_n360), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n359), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n275), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(new_n273), .B2(new_n218), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n270), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT11), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n326), .A2(new_n203), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n371), .B(KEYINPUT12), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n263), .A2(G68), .A3(new_n267), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n368), .B2(new_n369), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n365), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n306), .B1(new_n349), .B2(KEYINPUT13), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n376), .B1(new_n352), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n355), .A2(G200), .A3(new_n357), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT16), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n256), .A2(KEYINPUT74), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT74), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G33), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(new_n387), .A3(new_n284), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n286), .A2(KEYINPUT7), .A3(new_n231), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n285), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n203), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g0195(.A(G58), .B(G68), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(G20), .B1(G159), .B2(new_n275), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n384), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT75), .ZN(new_n400));
  XNOR2_X1  g0200(.A(KEYINPUT74), .B(G33), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n231), .B(new_n285), .C1(new_n401), .C2(new_n284), .ZN(new_n402));
  OAI21_X1  g0202(.A(G68), .B1(new_n402), .B2(KEYINPUT7), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n385), .A2(new_n387), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n338), .B1(new_n404), .B2(KEYINPUT3), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n393), .B1(new_n405), .B2(new_n231), .ZN(new_n406));
  OAI211_X1 g0206(.A(KEYINPUT16), .B(new_n397), .C1(new_n403), .C2(new_n406), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n388), .A2(new_n389), .B1(new_n392), .B2(new_n393), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n397), .B1(new_n408), .B2(new_n203), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT75), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n410), .A3(new_n384), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n400), .A2(new_n407), .A3(new_n270), .A4(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n271), .A2(new_n265), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n263), .A2(new_n413), .B1(new_n326), .B2(new_n271), .ZN(new_n414));
  INV_X1    g0214(.A(G200), .ZN(new_n415));
  MUX2_X1   g0215(.A(G223), .B(G226), .S(G1698), .Z(new_n416));
  AOI21_X1  g0216(.A(new_n284), .B1(new_n385), .B2(new_n387), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n416), .B1(new_n417), .B2(new_n338), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G87), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n299), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n302), .A2(G232), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n300), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n415), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n299), .A2(G274), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n297), .A2(new_n425), .B1(new_n302), .B2(G232), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n285), .B1(new_n401), .B2(new_n284), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n427), .A2(new_n416), .B1(G33), .B2(G87), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n426), .B1(new_n428), .B2(new_n299), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n423), .B1(G190), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n412), .A2(new_n414), .A3(new_n430), .ZN(new_n431));
  XOR2_X1   g0231(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(KEYINPUT76), .A2(KEYINPUT17), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n412), .A2(new_n414), .A3(new_n430), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n414), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n407), .A2(new_n270), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n286), .A2(KEYINPUT7), .A3(new_n231), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n440), .B1(new_n401), .B2(new_n284), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT7), .B1(new_n285), .B2(new_n391), .ZN(new_n442));
  OAI21_X1  g0242(.A(G68), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI211_X1 g0243(.A(KEYINPUT75), .B(KEYINPUT16), .C1(new_n443), .C2(new_n397), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n410), .B1(new_n409), .B2(new_n384), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n438), .B1(new_n439), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(G169), .B1(new_n420), .B2(new_n422), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n426), .B(G179), .C1(new_n428), .C2(new_n299), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(KEYINPUT18), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n450), .B1(new_n412), .B2(new_n414), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT18), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n437), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  NOR4_X1   g0255(.A1(new_n336), .A2(new_n378), .A3(new_n383), .A4(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(G238), .A2(G1698), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n457), .B1(new_n219), .B2(G1698), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(new_n417), .B2(new_n338), .ZN(new_n459));
  INV_X1    g0259(.A(G116), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n401), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n299), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n260), .A2(G45), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(new_n215), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n299), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n424), .B2(new_n464), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n320), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n425), .A2(new_n465), .B1(new_n466), .B2(new_n299), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n461), .B1(new_n427), .B2(new_n458), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n312), .B(new_n470), .C1(new_n471), .C2(new_n299), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n324), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(new_n261), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT19), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n231), .B1(new_n341), .B2(new_n476), .ZN(new_n477));
  OR2_X1    g0277(.A1(KEYINPUT77), .A2(G97), .ZN(new_n478));
  NAND2_X1  g0278(.A1(KEYINPUT77), .A2(G97), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n478), .A2(new_n214), .A3(new_n207), .A4(new_n479), .ZN(new_n480));
  AND2_X1   g0280(.A1(KEYINPUT77), .A2(G97), .ZN(new_n481));
  NOR2_X1   g0281(.A1(KEYINPUT77), .A2(G97), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n272), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n477), .A2(new_n480), .B1(new_n483), .B2(new_n476), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n231), .B(G68), .C1(new_n417), .C2(new_n338), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n475), .B1(new_n486), .B2(new_n270), .ZN(new_n487));
  AND2_X1   g0287(.A1(G1), .A2(G13), .ZN(new_n488));
  AND3_X1   g0288(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n488), .B1(new_n489), .B2(new_n258), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n256), .A2(G1), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n490), .A2(new_n257), .A3(new_n261), .A4(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(new_n324), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT81), .B1(new_n487), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n270), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n497), .B1(new_n484), .B2(new_n485), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT81), .ZN(new_n499));
  NOR4_X1   g0299(.A1(new_n498), .A2(new_n494), .A3(new_n499), .A4(new_n475), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n473), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n470), .B1(new_n471), .B2(new_n299), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G200), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n262), .A2(new_n491), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G87), .ZN(new_n505));
  OAI211_X1 g0305(.A(G190), .B(new_n470), .C1(new_n471), .C2(new_n299), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n503), .A2(new_n487), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT82), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n276), .A2(new_n218), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT6), .ZN(new_n511));
  AND2_X1   g0311(.A1(G97), .A2(G107), .ZN(new_n512));
  NOR2_X1   g0312(.A1(G97), .A2(G107), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n481), .A2(new_n482), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n207), .A2(KEYINPUT6), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n510), .B1(new_n517), .B2(G20), .ZN(new_n518));
  OAI21_X1  g0318(.A(G107), .B1(new_n441), .B2(new_n442), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n497), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n493), .A2(new_n206), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n261), .A2(G97), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  XOR2_X1   g0323(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n524));
  NOR2_X1   g0324(.A1(new_n219), .A2(G1698), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n524), .B1(new_n405), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G283), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT79), .ZN(new_n529));
  XNOR2_X1  g0329(.A(new_n528), .B(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(G250), .B(G1698), .C1(new_n337), .C2(new_n338), .ZN(new_n531));
  AND2_X1   g0331(.A1(KEYINPUT4), .A2(G244), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n288), .B(new_n532), .C1(new_n337), .C2(new_n338), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n299), .B1(new_n527), .B2(new_n535), .ZN(new_n536));
  OR2_X1    g0336(.A1(KEYINPUT5), .A2(G41), .ZN(new_n537));
  NAND2_X1  g0337(.A1(KEYINPUT5), .A2(G41), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n464), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n425), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g0340(.A(KEYINPUT5), .B(G41), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n541), .A2(new_n465), .B1(new_n488), .B2(new_n298), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(G257), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n540), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n536), .A2(G190), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n524), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(new_n427), .B2(new_n525), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n293), .B1(new_n548), .B2(new_n534), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n542), .A2(G257), .B1(new_n425), .B2(new_n539), .ZN(new_n550));
  AOI21_X1  g0350(.A(G200), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n523), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n320), .B1(new_n536), .B2(new_n545), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n516), .B1(new_n478), .B2(new_n479), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G97), .A2(G107), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT6), .B1(new_n208), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(G20), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n510), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n207), .B1(new_n390), .B2(new_n394), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n270), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n521), .ZN(new_n562));
  INV_X1    g0362(.A(new_n522), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n549), .A2(new_n312), .A3(new_n550), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n553), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n552), .A2(KEYINPUT80), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT80), .B1(new_n552), .B2(new_n566), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n508), .B(new_n509), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n508), .B1(new_n567), .B2(new_n568), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT82), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n460), .A2(G20), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n528), .A2(new_n529), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT79), .B1(G33), .B2(G283), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n231), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(G33), .B1(new_n478), .B2(new_n479), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n270), .B(new_n572), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT20), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n256), .B1(new_n481), .B2(new_n482), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n530), .A2(new_n231), .A3(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n581), .A2(KEYINPUT20), .A3(new_n270), .A4(new_n572), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n326), .A2(new_n460), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT83), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n493), .B2(new_n460), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n504), .A2(KEYINPUT83), .A3(G116), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n583), .A2(new_n584), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n541), .A2(new_n465), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n589), .A2(G270), .A3(new_n299), .ZN(new_n590));
  NOR2_X1   g0390(.A1(G257), .A2(G1698), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n220), .B2(G1698), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(G303), .ZN(new_n594));
  OAI22_X1  g0394(.A1(new_n405), .A2(new_n593), .B1(new_n594), .B2(new_n287), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n590), .B1(new_n595), .B2(new_n293), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n320), .B1(new_n596), .B2(new_n540), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n588), .A2(new_n597), .A3(KEYINPUT21), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n542), .A2(G270), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n337), .A2(new_n338), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n427), .A2(new_n592), .B1(G303), .B2(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n540), .B(new_n599), .C1(new_n601), .C2(new_n299), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n602), .A2(new_n312), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n588), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n598), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n602), .A2(G200), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n306), .B2(new_n602), .ZN(new_n608));
  OR2_X1    g0408(.A1(new_n608), .A2(new_n588), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n588), .A2(new_n597), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT21), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n606), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(G250), .A2(G1698), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n544), .B2(G1698), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n417), .B2(new_n338), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n404), .A2(G294), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n293), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n542), .A2(G264), .B1(new_n425), .B2(new_n539), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(G179), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT86), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n320), .B1(new_n619), .B2(new_n620), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT86), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n326), .A2(new_n207), .ZN(new_n628));
  XNOR2_X1  g0428(.A(new_n628), .B(KEYINPUT25), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(G107), .B2(new_n504), .ZN(new_n630));
  XOR2_X1   g0430(.A(KEYINPUT84), .B(KEYINPUT24), .Z(new_n631));
  NOR2_X1   g0431(.A1(new_n631), .A2(KEYINPUT85), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(KEYINPUT85), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT22), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(new_n214), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n231), .B(new_n636), .C1(new_n417), .C2(new_n338), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n231), .A2(G87), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n635), .B1(new_n600), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n404), .A2(new_n231), .A3(G116), .ZN(new_n641));
  OAI21_X1  g0441(.A(KEYINPUT23), .B1(new_n231), .B2(G107), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT23), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n643), .A2(new_n207), .A3(G20), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n640), .A2(new_n641), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n634), .B1(new_n638), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n645), .B1(new_n461), .B2(new_n231), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n649), .A2(new_n633), .A3(new_n637), .A4(new_n640), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n632), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n630), .B1(new_n651), .B2(new_n497), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n627), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n299), .B1(new_n616), .B2(new_n617), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n589), .A2(G264), .A3(new_n299), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n540), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n415), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n427), .A2(new_n615), .B1(G294), .B2(new_n404), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n620), .B(new_n306), .C1(new_n658), .C2(new_n299), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n660), .B(new_n630), .C1(new_n651), .C2(new_n497), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n653), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n613), .A2(new_n662), .ZN(new_n663));
  AND4_X1   g0463(.A1(new_n456), .A2(new_n569), .A3(new_n571), .A4(new_n663), .ZN(G372));
  AND3_X1   g0464(.A1(new_n553), .A2(new_n564), .A3(new_n565), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n501), .A2(new_n665), .A3(new_n507), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n501), .A2(new_n665), .A3(KEYINPUT26), .A4(new_n507), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n661), .A2(new_n552), .A3(new_n566), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n612), .A2(new_n604), .A3(new_n598), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n648), .A2(new_n650), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n270), .B1(new_n673), .B2(new_n632), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n674), .A2(new_n630), .B1(new_n623), .B2(new_n626), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n671), .B(new_n508), .C1(new_n672), .C2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n670), .A2(new_n676), .A3(new_n501), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n456), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n314), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n383), .A2(new_n330), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n437), .B1(new_n378), .B2(new_n680), .ZN(new_n681));
  AOI211_X1 g0481(.A(KEYINPUT18), .B(new_n450), .C1(new_n414), .C2(new_n412), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n412), .A2(new_n414), .ZN(new_n683));
  INV_X1    g0483(.A(new_n450), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n453), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n679), .B1(new_n687), .B2(new_n310), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n678), .A2(new_n688), .ZN(G369));
  NAND3_X1  g0489(.A1(new_n260), .A2(new_n231), .A3(G13), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT27), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n692), .A2(new_n260), .A3(new_n231), .A4(G13), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n691), .A2(G213), .A3(G343), .A4(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT87), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n693), .A2(G213), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT87), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n696), .A2(new_n697), .A3(G343), .A4(new_n691), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT21), .B1(new_n588), .B2(new_n597), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n700), .B1(new_n605), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT91), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n695), .A2(new_n698), .A3(KEYINPUT91), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI22_X1  g0506(.A1(new_n662), .A2(new_n702), .B1(new_n653), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(KEYINPUT88), .B1(new_n588), .B2(new_n699), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT88), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n579), .A2(new_n582), .B1(new_n460), .B2(new_n326), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n587), .A2(new_n586), .ZN(new_n711));
  AOI211_X1 g0511(.A(new_n709), .B(new_n700), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n605), .A2(new_n701), .B1(new_n708), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT89), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n712), .A2(new_n708), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n606), .A2(new_n715), .A3(new_n609), .A4(new_n612), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT89), .ZN(new_n717));
  OAI221_X1 g0517(.A(new_n717), .B1(new_n712), .B2(new_n708), .C1(new_n605), .C2(new_n701), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n714), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n719), .A2(KEYINPUT90), .A3(G330), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(KEYINPUT90), .B1(new_n719), .B2(G330), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n652), .A2(new_n699), .ZN(new_n725));
  OAI22_X1  g0525(.A1(new_n662), .A2(new_n725), .B1(new_n653), .B2(new_n700), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n707), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  XOR2_X1   g0527(.A(new_n727), .B(KEYINPUT92), .Z(G399));
  INV_X1    g0528(.A(new_n227), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G41), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n480), .A2(G116), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n731), .A2(G1), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(new_n234), .B2(new_n731), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT93), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT28), .ZN(new_n736));
  INV_X1    g0536(.A(new_n706), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n677), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT29), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT96), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(new_n677), .B2(new_n700), .ZN(new_n742));
  INV_X1    g0542(.A(new_n501), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n743), .B1(new_n668), .B2(new_n669), .ZN(new_n744));
  AOI211_X1 g0544(.A(KEYINPUT96), .B(new_n699), .C1(new_n744), .C2(new_n676), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n740), .B1(new_n746), .B2(new_n739), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT95), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n602), .B1(new_n536), .B2(new_n545), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n502), .B(new_n312), .C1(new_n654), .C2(new_n656), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n599), .B1(new_n601), .B2(new_n299), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n502), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n536), .A2(new_n545), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n622), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(KEYINPUT30), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT30), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n622), .A2(new_n753), .A3(new_n754), .A4(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n751), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  XOR2_X1   g0559(.A(KEYINPUT94), .B(KEYINPUT31), .Z(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n706), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n748), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n759), .A2(new_n700), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n763), .B1(new_n764), .B2(KEYINPUT31), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n759), .A2(new_n748), .A3(new_n762), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n571), .A2(new_n663), .A3(new_n569), .A4(new_n737), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G330), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n747), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n736), .B1(new_n772), .B2(G1), .ZN(G364));
  INV_X1    g0573(.A(new_n724), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n231), .A2(G13), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n260), .B1(new_n775), .B2(G45), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n774), .B1(G330), .B2(new_n719), .C1(new_n730), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n730), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT97), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n729), .A2(new_n600), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G355), .A2(new_n782), .B1(new_n460), .B2(new_n729), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n254), .A2(new_n296), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n427), .A2(new_n729), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(G45), .B2(new_n234), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n783), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G13), .A2(G33), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT98), .Z(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n230), .B1(G20), .B2(new_n320), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G179), .A2(G200), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(G20), .B1(new_n795), .B2(new_n306), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT102), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n796), .A2(new_n797), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n231), .A2(new_n312), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n803), .A2(G190), .A3(G200), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(KEYINPUT99), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n804), .A2(KEYINPUT99), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G294), .A2(new_n802), .B1(new_n809), .B2(G326), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n231), .A2(G190), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n794), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n812), .A2(KEYINPUT101), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(KEYINPUT101), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G329), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n231), .A2(new_n306), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n312), .A2(G200), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G322), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n811), .A2(new_n819), .ZN(new_n822));
  INV_X1    g0622(.A(G311), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n820), .A2(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n415), .A2(G179), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n818), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n803), .A2(new_n306), .A3(G200), .ZN(new_n827));
  XOR2_X1   g0627(.A(KEYINPUT33), .B(G317), .Z(new_n828));
  OAI221_X1 g0628(.A(new_n600), .B1(new_n826), .B2(new_n594), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n811), .A2(new_n825), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n824), .B(new_n829), .C1(G283), .C2(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n810), .A2(new_n817), .A3(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(G159), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n815), .A2(new_n834), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT32), .Z(new_n836));
  NOR2_X1   g0636(.A1(new_n826), .A2(new_n214), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n600), .B(new_n837), .C1(G107), .C2(new_n831), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n838), .B1(new_n203), .B2(new_n827), .C1(new_n206), .C2(new_n801), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n820), .A2(new_n202), .B1(new_n822), .B2(new_n218), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(new_n809), .B2(G50), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT100), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n833), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n781), .B(new_n793), .C1(new_n844), .C2(new_n791), .ZN(new_n845));
  INV_X1    g0645(.A(new_n790), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n845), .B1(new_n719), .B2(new_n846), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n778), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G396));
  INV_X1    g0649(.A(new_n791), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n789), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT103), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n780), .B1(new_n852), .B2(G77), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT104), .Z(new_n854));
  INV_X1    g0654(.A(new_n820), .ZN(new_n855));
  INV_X1    g0655(.A(new_n822), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G143), .A2(new_n855), .B1(new_n856), .B2(G159), .ZN(new_n857));
  INV_X1    g0657(.A(G137), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n857), .B1(new_n274), .B2(new_n827), .C1(new_n808), .C2(new_n858), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT34), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n427), .B1(new_n201), .B2(new_n826), .C1(new_n203), .C2(new_n830), .ZN(new_n861));
  INV_X1    g0661(.A(G132), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n815), .A2(new_n862), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n861), .B(new_n863), .C1(new_n802), .C2(G58), .ZN(new_n864));
  INV_X1    g0664(.A(G283), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n600), .B1(new_n822), .B2(new_n460), .C1(new_n827), .C2(new_n865), .ZN(new_n866));
  AOI22_X1  g0666(.A1(G294), .A2(new_n855), .B1(new_n831), .B2(G87), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n207), .B2(new_n826), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n866), .B(new_n868), .C1(G311), .C2(new_n816), .ZN(new_n869));
  AOI22_X1  g0669(.A1(G97), .A2(new_n802), .B1(new_n809), .B2(G303), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n860), .A2(new_n864), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n331), .A2(new_n700), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n334), .A2(new_n332), .B1(new_n329), .B2(new_n699), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n872), .B1(new_n873), .B2(new_n331), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  OAI221_X1 g0675(.A(new_n854), .B1(new_n850), .B2(new_n871), .C1(new_n875), .C2(new_n789), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n738), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n878), .A2(new_n875), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n706), .B(new_n874), .C1(new_n744), .C2(new_n676), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n882), .A2(new_n770), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n779), .B1(new_n882), .B2(new_n770), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n877), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(G384));
  OR2_X1    g0687(.A1(new_n517), .A2(KEYINPUT35), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n517), .A2(KEYINPUT35), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n888), .A2(G116), .A3(new_n232), .A4(new_n889), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n890), .B(KEYINPUT36), .Z(new_n891));
  OAI211_X1 g0691(.A(new_n235), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n260), .B(G13), .C1(new_n892), .C2(new_n250), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n696), .A2(new_n691), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n412), .B2(new_n414), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n451), .A2(new_n454), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT107), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n434), .B2(new_n436), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n434), .A2(new_n900), .A3(new_n436), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n898), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n412), .A2(new_n414), .A3(new_n430), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n905), .A2(new_n452), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n906), .A2(KEYINPUT106), .A3(KEYINPUT37), .A4(new_n898), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT37), .B1(new_n897), .B2(KEYINPUT106), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n431), .B1(new_n447), .B2(new_n450), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n908), .B1(new_n909), .B2(new_n897), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n895), .B1(new_n904), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n407), .A2(new_n270), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n405), .A2(new_n393), .A3(new_n231), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n402), .A2(KEYINPUT7), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(new_n915), .A3(G68), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT16), .B1(new_n916), .B2(new_n397), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n414), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n896), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n455), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n918), .A2(new_n684), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(new_n920), .A3(new_n431), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT37), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n897), .A2(KEYINPUT37), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n906), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n922), .A2(KEYINPUT38), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT39), .B1(new_n912), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n920), .B1(new_n686), .B2(new_n437), .ZN(new_n931));
  AOI22_X1  g0731(.A1(KEYINPUT37), .A2(new_n924), .B1(new_n906), .B2(new_n926), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n895), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n929), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT39), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n378), .A2(new_n700), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n930), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n364), .B1(new_n360), .B2(new_n358), .ZN(new_n939));
  INV_X1    g0739(.A(new_n359), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n376), .B(new_n699), .C1(new_n941), .C2(new_n383), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n376), .A2(new_n699), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n382), .B(new_n943), .C1(new_n365), .C2(new_n377), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n872), .B(KEYINPUT105), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n945), .B1(new_n880), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n934), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n947), .A2(new_n948), .B1(new_n686), .B2(new_n919), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n938), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n456), .B(new_n740), .C1(new_n746), .C2(new_n739), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n688), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n950), .B(new_n952), .Z(new_n953));
  INV_X1    g0753(.A(G330), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n874), .B1(new_n942), .B2(new_n944), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT108), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT31), .B1(new_n956), .B2(KEYINPUT94), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n759), .A2(new_n700), .A3(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n759), .A2(new_n700), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n761), .A2(new_n956), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n768), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n955), .A2(new_n934), .A3(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT40), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n437), .A2(KEYINPUT107), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n966), .A2(new_n686), .A3(new_n903), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n911), .B1(new_n897), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n929), .B1(new_n968), .B2(KEYINPUT38), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n969), .A2(KEYINPUT40), .A3(new_n962), .A4(new_n955), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n965), .A2(new_n970), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n456), .A2(new_n962), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n954), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n971), .B2(new_n972), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n953), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n260), .B2(new_n775), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n953), .A2(new_n974), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n894), .B1(new_n976), .B2(new_n977), .ZN(G367));
  INV_X1    g0778(.A(KEYINPUT111), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT42), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n662), .A2(new_n702), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n553), .A2(new_n565), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n564), .A2(new_n706), .ZN(new_n983));
  NOR3_X1   g0783(.A1(new_n982), .A2(new_n983), .A3(KEYINPUT110), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT110), .ZN(new_n985));
  INV_X1    g0785(.A(new_n983), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n553), .A2(new_n565), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n552), .A2(new_n566), .A3(new_n983), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n984), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n980), .B1(new_n981), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n986), .A2(new_n987), .A3(new_n985), .ZN(new_n992));
  AND3_X1   g0792(.A1(new_n552), .A2(new_n566), .A3(new_n983), .ZN(new_n993));
  OAI21_X1  g0793(.A(KEYINPUT110), .B1(new_n982), .B2(new_n983), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n675), .B(new_n992), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n706), .B1(new_n995), .B2(new_n566), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n979), .B1(new_n991), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n672), .A2(new_n653), .A3(new_n661), .A4(new_n700), .ZN(new_n999));
  OAI21_X1  g0799(.A(KEYINPUT42), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n665), .B1(new_n990), .B2(new_n675), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n1000), .B(KEYINPUT111), .C1(new_n706), .C2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  NOR3_X1   g0803(.A1(new_n998), .A2(new_n999), .A3(KEYINPUT42), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(KEYINPUT112), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT112), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1003), .A2(new_n1008), .A3(new_n1005), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n501), .A2(new_n507), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n700), .B1(new_n487), .B2(new_n505), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT109), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n743), .A2(new_n1011), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT43), .Z(new_n1018));
  NAND3_X1  g0818(.A1(new_n1007), .A2(new_n1009), .A3(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1017), .A2(KEYINPUT43), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1008), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1021));
  AOI211_X1 g0821(.A(KEYINPUT112), .B(new_n1004), .C1(new_n997), .C2(new_n1002), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n726), .B1(new_n720), .B2(new_n722), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1024), .A2(new_n998), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1019), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT113), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1019), .A2(new_n1023), .A3(KEYINPUT113), .A4(new_n1025), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1024), .A2(KEYINPUT114), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT114), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1032), .B(new_n726), .C1(new_n720), .C2(new_n722), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT45), .ZN(new_n1034));
  OR3_X1    g0834(.A1(new_n707), .A2(new_n1034), .A3(new_n998), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1034), .B1(new_n707), .B2(new_n998), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n707), .A2(new_n998), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT44), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n707), .A2(KEYINPUT44), .A3(new_n998), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n1035), .A2(new_n1036), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1031), .A2(new_n1033), .A3(new_n1041), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1044));
  OAI211_X1 g0844(.A(KEYINPUT114), .B(new_n1024), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n702), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n999), .B1(new_n726), .B2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n724), .B(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n771), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n730), .B(KEYINPUT41), .Z(new_n1051));
  OAI21_X1  g0851(.A(new_n776), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n1024), .B2(new_n998), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1030), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT115), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1030), .A2(new_n1052), .A3(KEYINPUT115), .A4(new_n1054), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n792), .B1(new_n227), .B2(new_n324), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n785), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1061), .A2(new_n245), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n780), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n801), .A2(new_n203), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n820), .A2(new_n274), .B1(new_n830), .B2(new_n218), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n287), .B1(new_n822), .B2(new_n201), .C1(new_n827), .C2(new_n834), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n826), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1065), .B(new_n1066), .C1(G58), .C2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n858), .B2(new_n815), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1064), .B(new_n1069), .C1(G143), .C2(new_n809), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n801), .A2(new_n207), .B1(new_n808), .B2(new_n823), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n826), .A2(new_n460), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n427), .B1(new_n1072), .B2(KEYINPUT46), .ZN(new_n1073));
  INV_X1    g0873(.A(G294), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1073), .B1(KEYINPUT46), .B2(new_n1072), .C1(new_n1074), .C2(new_n827), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G303), .A2(new_n855), .B1(new_n856), .B2(G283), .ZN(new_n1076));
  INV_X1    g0876(.A(G317), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1076), .B1(new_n515), .B2(new_n830), .C1(new_n815), .C2(new_n1077), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1071), .A2(new_n1075), .A3(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1070), .A2(new_n1079), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT47), .Z(new_n1081));
  AOI21_X1  g0881(.A(new_n1063), .B1(new_n1081), .B2(new_n791), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1017), .A2(new_n846), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1059), .A2(new_n1084), .ZN(G387));
  AND2_X1   g0885(.A1(new_n772), .A2(new_n1049), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1086), .A2(new_n731), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n772), .B2(new_n1049), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n726), .A2(new_n846), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G317), .A2(new_n855), .B1(new_n856), .B2(G303), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(new_n823), .B2(new_n827), .C1(new_n808), .C2(new_n821), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT48), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n802), .A2(G283), .B1(G294), .B2(new_n1067), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT49), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n405), .B1(new_n460), .B2(new_n830), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n816), .B2(G326), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1098), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G50), .A2(new_n855), .B1(new_n831), .B2(G97), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1103), .B1(new_n203), .B2(new_n822), .C1(new_n218), .C2(new_n826), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n827), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n405), .B(new_n1104), .C1(new_n322), .C2(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n474), .A2(new_n802), .B1(new_n809), .B2(G159), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(new_n274), .C2(new_n815), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n850), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n785), .B1(new_n242), .B2(new_n296), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n782), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1110), .B1(new_n732), .B2(new_n1111), .ZN(new_n1112));
  OR3_X1    g0912(.A1(new_n271), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1113));
  AOI21_X1  g0913(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1114));
  OAI21_X1  g0914(.A(KEYINPUT50), .B1(new_n271), .B2(G50), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1113), .A2(new_n732), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(G107), .B2(new_n227), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n781), .B(new_n1109), .C1(new_n792), .C2(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1049), .A2(new_n777), .B1(new_n1089), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1088), .A2(new_n1120), .ZN(G393));
  OR2_X1    g0921(.A1(new_n1086), .A2(new_n1046), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n731), .B1(new_n1086), .B2(new_n1046), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1046), .A2(new_n777), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n990), .A2(new_n846), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1061), .A2(new_n249), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n792), .B1(new_n227), .B2(new_n515), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n802), .A2(G116), .B1(G303), .B2(new_n1105), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1129), .A2(KEYINPUT116), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1129), .A2(KEYINPUT116), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n815), .A2(new_n821), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n287), .B1(new_n831), .B2(G107), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1133), .B1(new_n865), .B2(new_n826), .C1(new_n1074), .C2(new_n822), .ZN(new_n1134));
  NOR4_X1   g0934(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .A4(new_n1134), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n808), .A2(new_n1077), .B1(new_n823), .B2(new_n820), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT52), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n808), .A2(new_n274), .B1(new_n834), .B2(new_n820), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT51), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n802), .A2(G77), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n816), .A2(G143), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n271), .A2(new_n822), .B1(new_n830), .B2(new_n214), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G68), .B2(new_n1067), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n405), .B1(G50), .B2(new_n1105), .ZN(new_n1144));
  AND4_X1   g0944(.A1(new_n1140), .A2(new_n1141), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1135), .A2(new_n1137), .B1(new_n1139), .B2(new_n1145), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n780), .B1(new_n1127), .B2(new_n1128), .C1(new_n1146), .C2(new_n850), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1125), .B1(new_n1126), .B2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1124), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(G390));
  NOR2_X1   g0950(.A1(new_n880), .A2(new_n946), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n945), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n770), .B2(new_n874), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n954), .B1(new_n768), .B2(new_n961), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1154), .A2(new_n875), .A3(new_n945), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1151), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n954), .B1(new_n767), .B2(new_n768), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1158), .A2(new_n955), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n873), .A2(new_n331), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n742), .B2(new_n745), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n872), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1159), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n962), .A2(G330), .A3(new_n875), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT119), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1165), .A2(new_n1166), .A3(new_n1152), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1166), .B1(new_n1165), .B2(new_n1152), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1164), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1157), .A2(new_n1170), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n456), .A2(new_n1154), .A3(KEYINPUT118), .ZN(new_n1172));
  AOI21_X1  g0972(.A(KEYINPUT118), .B1(new_n456), .B2(new_n1154), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n688), .B(new_n951), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1171), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1155), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT117), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n937), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n378), .A2(KEYINPUT117), .A3(new_n700), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n967), .A2(new_n897), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n911), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT38), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n929), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1179), .B(new_n1180), .C1(new_n1183), .C2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n1163), .B2(new_n945), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n948), .A2(KEYINPUT39), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n935), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1187), .A2(new_n1188), .B1(new_n937), .B2(new_n947), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1177), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n947), .A2(new_n937), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n930), .B2(new_n936), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1159), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1152), .B1(new_n1162), .B2(new_n872), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1192), .B(new_n1193), .C1(new_n1194), .C2(new_n1185), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1190), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1176), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1174), .B1(new_n1157), .B2(new_n1170), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1198), .A2(new_n1195), .A3(new_n1190), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1197), .A2(new_n1199), .A3(new_n730), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1196), .A2(new_n776), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n789), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n930), .B2(new_n936), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n780), .B1(new_n852), .B2(new_n322), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1140), .B1(new_n808), .B2(new_n865), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n816), .A2(G294), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n287), .B(new_n837), .C1(G107), .C2(new_n1105), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n855), .A2(G116), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n515), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(G68), .A2(new_n831), .B1(new_n856), .B2(new_n1209), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .A4(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(KEYINPUT54), .B(G143), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n820), .A2(new_n862), .B1(new_n822), .B2(new_n1212), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n600), .B(new_n1213), .C1(G50), .C2(new_n831), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n826), .A2(new_n274), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT53), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n1215), .A2(new_n1216), .B1(new_n858), .B2(new_n827), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n1216), .B2(new_n1215), .ZN(new_n1218));
  INV_X1    g1018(.A(G125), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1214), .B(new_n1218), .C1(new_n1219), .C2(new_n815), .ZN(new_n1220));
  INV_X1    g1020(.A(G128), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n801), .A2(new_n834), .B1(new_n808), .B2(new_n1221), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n1205), .A2(new_n1211), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1204), .B1(new_n1223), .B2(new_n791), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1201), .B1(new_n1203), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1200), .A2(new_n1225), .ZN(G378));
  NOR2_X1   g1026(.A1(new_n427), .A2(G41), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n831), .A2(G58), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT120), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1228), .B(new_n1231), .C1(G283), .C2(new_n816), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(G77), .A2(new_n1067), .B1(new_n856), .B2(new_n474), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n206), .B2(new_n827), .C1(new_n207), .C2(new_n820), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n808), .A2(new_n460), .ZN(new_n1236));
  NOR4_X1   g1036(.A1(new_n1233), .A2(new_n1235), .A3(new_n1064), .A4(new_n1236), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1237), .A2(KEYINPUT58), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n1221), .A2(new_n820), .B1(new_n826), .B2(new_n1212), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G137), .B2(new_n856), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n862), .B2(new_n827), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(G150), .B2(new_n802), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n1219), .B2(new_n808), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1243), .A2(KEYINPUT59), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(KEYINPUT59), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n816), .A2(G124), .ZN(new_n1246));
  AOI211_X1 g1046(.A(G33), .B(G41), .C1(new_n831), .C2(G159), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1237), .A2(KEYINPUT58), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1228), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1238), .A2(new_n1248), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n791), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n852), .A2(G50), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1253), .A2(new_n730), .A3(new_n777), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n310), .A2(new_n314), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1255), .B(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n280), .A2(new_n919), .ZN(new_n1258));
  XOR2_X1   g1058(.A(new_n1258), .B(KEYINPUT121), .Z(new_n1259));
  XNOR2_X1  g1059(.A(new_n1257), .B(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1252), .B(new_n1254), .C1(new_n1261), .C2(new_n789), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n965), .A2(new_n970), .A3(G330), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT122), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n965), .A2(new_n970), .A3(KEYINPUT122), .A4(G330), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1266), .A2(new_n1267), .A3(new_n1261), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n971), .A2(new_n1260), .A3(KEYINPUT122), .A4(G330), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n950), .A3(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n950), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1263), .B1(new_n1273), .B2(new_n777), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1168), .A2(new_n1159), .A3(new_n1163), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1156), .B1(new_n1275), .B2(new_n1167), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1175), .B1(new_n1196), .B2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT57), .B1(new_n1273), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n950), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1281), .A2(KEYINPUT57), .A3(new_n1277), .A4(new_n1270), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n730), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1274), .B1(new_n1278), .B2(new_n1283), .ZN(G375));
  XOR2_X1   g1084(.A(new_n776), .B(KEYINPUT123), .Z(new_n1285));
  NAND2_X1  g1085(.A1(new_n1171), .A2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n780), .B1(new_n852), .B2(G68), .ZN(new_n1287));
  OAI22_X1  g1087(.A1(new_n826), .A2(new_n834), .B1(new_n822), .B2(new_n274), .ZN(new_n1288));
  NOR3_X1   g1088(.A1(new_n1231), .A2(new_n405), .A3(new_n1288), .ZN(new_n1289));
  OAI221_X1 g1089(.A(new_n1289), .B1(new_n201), .B2(new_n801), .C1(new_n1221), .C2(new_n815), .ZN(new_n1290));
  XOR2_X1   g1090(.A(new_n1290), .B(KEYINPUT124), .Z(new_n1291));
  OAI22_X1  g1091(.A1(new_n827), .A2(new_n1212), .B1(new_n820), .B2(new_n858), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1292), .B1(new_n809), .B2(G132), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1294));
  OAI22_X1  g1094(.A1(new_n820), .A2(new_n865), .B1(new_n822), .B2(new_n207), .ZN(new_n1295));
  OAI221_X1 g1095(.A(new_n600), .B1(new_n830), .B2(new_n218), .C1(new_n827), .C2(new_n460), .ZN(new_n1296));
  AOI211_X1 g1096(.A(new_n1295), .B(new_n1296), .C1(G97), .C2(new_n1067), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1297), .B1(new_n594), .B2(new_n815), .ZN(new_n1298));
  OAI22_X1  g1098(.A1(new_n801), .A2(new_n324), .B1(new_n808), .B2(new_n1074), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1294), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1287), .B1(new_n1300), .B2(new_n791), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(new_n789), .B2(new_n945), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1286), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1276), .A2(new_n1174), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1051), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1176), .A2(new_n1305), .A3(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1304), .A2(new_n1307), .ZN(G381));
  NOR2_X1   g1108(.A1(G393), .A2(G396), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1149), .A2(new_n1309), .A3(new_n886), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n1310), .A2(G378), .A3(G381), .ZN(new_n1311));
  AOI22_X1  g1111(.A1(new_n1057), .A2(new_n1058), .B1(new_n1083), .B2(new_n1082), .ZN(new_n1312));
  INV_X1    g1112(.A(G375), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1311), .A2(new_n1312), .A3(new_n1313), .ZN(G407));
  INV_X1    g1114(.A(G378), .ZN(new_n1315));
  INV_X1    g1115(.A(G213), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1316), .A2(G343), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1313), .A2(new_n1315), .A3(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(G407), .A2(G213), .A3(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT125), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(new_n1319), .B(new_n1320), .ZN(G409));
  INV_X1    g1121(.A(KEYINPUT126), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(G387), .A2(new_n1322), .A3(G390), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1149), .B1(new_n1312), .B2(KEYINPUT126), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n848), .B1(new_n1088), .B2(new_n1120), .ZN(new_n1326));
  AOI211_X1 g1126(.A(new_n1309), .B(new_n1326), .C1(new_n1312), .C2(KEYINPUT126), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1309), .A2(new_n1326), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT127), .B1(new_n1059), .B2(new_n1084), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1328), .B1(new_n1329), .B2(G390), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1149), .B1(new_n1312), .B2(KEYINPUT127), .ZN(new_n1331));
  AOI22_X1  g1131(.A1(new_n1325), .A2(new_n1327), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  OAI211_X1 g1132(.A(G378), .B(new_n1274), .C1(new_n1278), .C2(new_n1283), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1281), .A2(new_n1270), .A3(new_n1285), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1281), .A2(new_n1277), .A3(new_n1270), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1262), .B(new_n1334), .C1(new_n1335), .C2(new_n1051), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1315), .A2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1333), .A2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1317), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1317), .A2(G2897), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1341), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1157), .A2(new_n1170), .A3(KEYINPUT60), .A4(new_n1174), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(new_n730), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1176), .A2(KEYINPUT60), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1344), .B1(new_n1345), .B2(new_n1305), .ZN(new_n1346));
  NOR3_X1   g1146(.A1(new_n1346), .A2(new_n886), .A3(new_n1303), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT60), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1305), .B1(new_n1198), .B2(new_n1348), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1349), .A2(new_n730), .A3(new_n1343), .ZN(new_n1350));
  AOI21_X1  g1150(.A(G384), .B1(new_n1350), .B2(new_n1304), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1342), .B1(new_n1347), .B2(new_n1351), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n886), .B1(new_n1346), .B2(new_n1303), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1350), .A2(G384), .A3(new_n1304), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1353), .A2(new_n1354), .A3(new_n1341), .ZN(new_n1355));
  AND2_X1   g1155(.A1(new_n1352), .A2(new_n1355), .ZN(new_n1356));
  AOI21_X1  g1156(.A(KEYINPUT61), .B1(new_n1340), .B2(new_n1356), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1317), .B1(new_n1333), .B2(new_n1337), .ZN(new_n1358));
  NOR2_X1   g1158(.A1(new_n1347), .A2(new_n1351), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1358), .A2(KEYINPUT63), .A3(new_n1359), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1338), .A2(new_n1339), .A3(new_n1359), .ZN(new_n1361));
  INV_X1    g1161(.A(KEYINPUT63), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1357), .A2(new_n1360), .A3(new_n1363), .ZN(new_n1364));
  INV_X1    g1164(.A(KEYINPUT62), .ZN(new_n1365));
  AND3_X1   g1165(.A1(new_n1358), .A2(new_n1365), .A3(new_n1359), .ZN(new_n1366));
  AOI21_X1  g1166(.A(new_n1365), .B1(new_n1358), .B2(new_n1359), .ZN(new_n1367));
  NOR2_X1   g1167(.A1(new_n1366), .A2(new_n1367), .ZN(new_n1368));
  INV_X1    g1168(.A(KEYINPUT61), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1352), .A2(new_n1355), .ZN(new_n1370));
  OAI21_X1  g1170(.A(new_n1369), .B1(new_n1358), .B2(new_n1370), .ZN(new_n1371));
  NOR2_X1   g1171(.A1(new_n1332), .A2(new_n1371), .ZN(new_n1372));
  AOI22_X1  g1172(.A1(new_n1332), .A2(new_n1364), .B1(new_n1368), .B2(new_n1372), .ZN(G405));
  NAND2_X1  g1173(.A1(G375), .A2(new_n1315), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1374), .A2(new_n1333), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1375), .A2(new_n1359), .ZN(new_n1376));
  OAI211_X1 g1176(.A(new_n1374), .B(new_n1333), .C1(new_n1351), .C2(new_n1347), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1376), .A2(new_n1377), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1379), .A2(new_n1380), .ZN(new_n1381));
  XNOR2_X1  g1181(.A(new_n1378), .B(new_n1381), .ZN(G402));
endmodule


