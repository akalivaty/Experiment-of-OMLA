

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820;

  INV_X2 U379 ( .A(G119), .ZN(n698) );
  XNOR2_X1 U380 ( .A(KEYINPUT76), .B(KEYINPUT16), .ZN(n566) );
  XNOR2_X2 U381 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X2 U382 ( .A(n381), .B(n774), .ZN(n776) );
  NOR2_X2 U383 ( .A1(n441), .A2(n433), .ZN(n431) );
  OR2_X1 U384 ( .A1(n642), .A2(n710), .ZN(n643) );
  AND2_X1 U385 ( .A1(G227), .A2(n806), .ZN(n493) );
  NAND2_X1 U386 ( .A1(n490), .A2(n738), .ZN(n741) );
  XNOR2_X1 U387 ( .A(G134), .B(G122), .ZN(n562) );
  INV_X2 U388 ( .A(n653), .ZN(n490) );
  BUF_X1 U389 ( .A(G953), .Z(n812) );
  BUF_X1 U390 ( .A(G143), .Z(n819) );
  NOR2_X2 U391 ( .A1(n754), .A2(n756), .ZN(n614) );
  NAND2_X2 U392 ( .A1(n443), .A2(n447), .ZN(n427) );
  AND2_X2 U393 ( .A1(n599), .A2(KEYINPUT79), .ZN(n432) );
  XNOR2_X2 U394 ( .A(n384), .B(n536), .ZN(n599) );
  XNOR2_X1 U395 ( .A(n597), .B(KEYINPUT101), .ZN(n755) );
  NAND2_X1 U396 ( .A1(n686), .A2(n510), .ZN(n508) );
  INV_X4 U397 ( .A(G953), .ZN(n806) );
  NOR2_X1 U398 ( .A1(n772), .A2(n812), .ZN(n773) );
  NAND2_X1 U399 ( .A1(n409), .A2(n408), .ZN(n675) );
  AND2_X1 U400 ( .A1(n444), .A2(n445), .ZN(n443) );
  AND2_X1 U401 ( .A1(n375), .A2(n454), .ZN(n726) );
  OR2_X1 U402 ( .A1(n648), .A2(n635), .ZN(n637) );
  NOR2_X1 U403 ( .A1(n594), .A2(n379), .ZN(n615) );
  AND2_X1 U404 ( .A1(n484), .A2(n483), .ZN(n482) );
  OR2_X1 U405 ( .A1(n589), .A2(n590), .ZN(n368) );
  XOR2_X1 U406 ( .A(KEYINPUT10), .B(n575), .Z(n554) );
  XNOR2_X1 U407 ( .A(n425), .B(n424), .ZN(n558) );
  XNOR2_X1 U408 ( .A(n550), .B(G134), .ZN(n496) );
  XNOR2_X1 U409 ( .A(KEYINPUT74), .B(KEYINPUT14), .ZN(n420) );
  NOR2_X1 U410 ( .A1(G953), .A2(G237), .ZN(n543) );
  XNOR2_X2 U411 ( .A(KEYINPUT3), .B(G113), .ZN(n503) );
  INV_X2 U412 ( .A(G104), .ZN(n455) );
  XNOR2_X1 U413 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n574) );
  NAND2_X1 U414 ( .A1(n410), .A2(n412), .ZN(n403) );
  NAND2_X1 U415 ( .A1(n385), .A2(n727), .ZN(n356) );
  NAND2_X1 U416 ( .A1(n385), .A2(n727), .ZN(n805) );
  XNOR2_X2 U417 ( .A(n802), .B(G146), .ZN(n528) );
  NAND2_X1 U418 ( .A1(n577), .A2(n496), .ZN(n359) );
  NAND2_X1 U419 ( .A1(n357), .A2(n358), .ZN(n360) );
  NAND2_X1 U420 ( .A1(n360), .A2(n359), .ZN(n802) );
  INV_X1 U421 ( .A(n577), .ZN(n357) );
  INV_X1 U422 ( .A(n496), .ZN(n358) );
  XNOR2_X1 U423 ( .A(n805), .B(KEYINPUT77), .ZN(n402) );
  AND2_X2 U424 ( .A1(n488), .A2(n732), .ZN(n361) );
  BUF_X1 U425 ( .A(n528), .Z(n507) );
  XNOR2_X2 U426 ( .A(n438), .B(n440), .ZN(n385) );
  NAND2_X1 U427 ( .A1(n630), .A2(n476), .ZN(n475) );
  NAND2_X1 U428 ( .A1(n466), .A2(n659), .ZN(n465) );
  OR2_X1 U429 ( .A1(n608), .A2(n607), .ZN(n400) );
  INV_X1 U430 ( .A(G902), .ZN(n510) );
  INV_X1 U431 ( .A(n632), .ZN(n476) );
  INV_X1 U432 ( .A(KEYINPUT93), .ZN(n453) );
  XNOR2_X1 U433 ( .A(n399), .B(KEYINPUT84), .ZN(n398) );
  XOR2_X1 U434 ( .A(KEYINPUT5), .B(G119), .Z(n498) );
  XNOR2_X1 U435 ( .A(G116), .B(KEYINPUT98), .ZN(n500) );
  NOR2_X1 U436 ( .A1(n482), .A2(n475), .ZN(n474) );
  OR2_X1 U437 ( .A1(n666), .A2(n667), .ZN(n456) );
  NAND2_X1 U438 ( .A1(n463), .A2(n461), .ZN(n411) );
  INV_X1 U439 ( .A(KEYINPUT8), .ZN(n424) );
  NAND2_X1 U440 ( .A1(n806), .A2(G234), .ZN(n425) );
  INV_X1 U441 ( .A(G116), .ZN(n561) );
  XOR2_X1 U442 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n545) );
  INV_X1 U443 ( .A(n552), .ZN(n416) );
  XOR2_X1 U444 ( .A(KEYINPUT99), .B(G140), .Z(n547) );
  INV_X1 U445 ( .A(KEYINPUT90), .ZN(n440) );
  NAND2_X1 U446 ( .A1(n472), .A2(n468), .ZN(n648) );
  AND2_X1 U447 ( .A1(n470), .A2(n469), .ZN(n468) );
  AND2_X1 U448 ( .A1(n477), .A2(n473), .ZN(n472) );
  OR2_X1 U449 ( .A1(n630), .A2(n476), .ZN(n469) );
  XNOR2_X1 U450 ( .A(n614), .B(n423), .ZN(n749) );
  INV_X1 U451 ( .A(KEYINPUT41), .ZN(n423) );
  INV_X1 U452 ( .A(KEYINPUT78), .ZN(n434) );
  BUF_X1 U453 ( .A(n591), .Z(n653) );
  XNOR2_X1 U454 ( .A(n508), .B(n378), .ZN(n654) );
  XNOR2_X1 U455 ( .A(n601), .B(G472), .ZN(n378) );
  XNOR2_X1 U456 ( .A(n755), .B(n414), .ZN(n650) );
  INV_X1 U457 ( .A(KEYINPUT85), .ZN(n414) );
  INV_X1 U458 ( .A(KEYINPUT48), .ZN(n486) );
  INV_X1 U459 ( .A(KEYINPUT4), .ZN(n495) );
  XOR2_X1 U460 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n580) );
  INV_X1 U461 ( .A(KEYINPUT79), .ZN(n433) );
  AND2_X1 U462 ( .A1(n471), .A2(n480), .ZN(n467) );
  INV_X1 U463 ( .A(n475), .ZN(n471) );
  INV_X1 U464 ( .A(G137), .ZN(n499) );
  XNOR2_X1 U465 ( .A(G101), .B(G110), .ZN(n529) );
  XOR2_X1 U466 ( .A(KEYINPUT81), .B(G107), .Z(n530) );
  XNOR2_X1 U467 ( .A(G902), .B(KEYINPUT15), .ZN(n670) );
  XNOR2_X1 U468 ( .A(n420), .B(n537), .ZN(n538) );
  XNOR2_X1 U469 ( .A(n621), .B(KEYINPUT38), .ZN(n752) );
  INV_X1 U470 ( .A(G237), .ZN(n509) );
  NOR2_X1 U471 ( .A1(n595), .A2(KEYINPUT19), .ZN(n480) );
  INV_X1 U472 ( .A(KEYINPUT69), .ZN(n421) );
  INV_X1 U473 ( .A(n411), .ZN(n409) );
  XOR2_X1 U474 ( .A(KEYINPUT9), .B(KEYINPUT100), .Z(n560) );
  XNOR2_X1 U475 ( .A(n553), .B(n415), .ZN(n678) );
  XNOR2_X1 U476 ( .A(n554), .B(n416), .ZN(n415) );
  AND2_X1 U477 ( .A1(n446), .A2(n633), .ZN(n445) );
  NAND2_X1 U478 ( .A1(n418), .A2(KEYINPUT34), .ZN(n446) );
  NAND2_X1 U479 ( .A1(n595), .A2(KEYINPUT19), .ZN(n483) );
  XNOR2_X1 U480 ( .A(n517), .B(n516), .ZN(n519) );
  XNOR2_X1 U481 ( .A(n515), .B(n514), .ZN(n517) );
  NOR2_X1 U482 ( .A1(n618), .A2(n454), .ZN(n620) );
  NAND2_X1 U483 ( .A1(n749), .A2(n615), .ZN(n616) );
  XNOR2_X1 U484 ( .A(KEYINPUT109), .B(KEYINPUT40), .ZN(n611) );
  XNOR2_X1 U485 ( .A(n377), .B(n376), .ZN(n375) );
  INV_X1 U486 ( .A(KEYINPUT36), .ZN(n376) );
  NAND2_X1 U487 ( .A1(n657), .A2(n362), .ZN(n485) );
  XNOR2_X1 U488 ( .A(n389), .B(n388), .ZN(n818) );
  INV_X1 U489 ( .A(KEYINPUT108), .ZN(n388) );
  INV_X1 U490 ( .A(n741), .ZN(n487) );
  AND2_X1 U491 ( .A1(n450), .A2(n490), .ZN(n655) );
  AND2_X1 U492 ( .A1(n369), .A2(n654), .ZN(n362) );
  OR2_X1 U493 ( .A1(G902), .A2(n783), .ZN(n363) );
  XNOR2_X1 U494 ( .A(KEYINPUT83), .B(n672), .ZN(n364) );
  AND2_X1 U495 ( .A1(n604), .A2(n717), .ZN(n365) );
  AND2_X1 U496 ( .A1(n664), .A2(n459), .ZN(n366) );
  BUF_X1 U497 ( .A(n648), .Z(n418) );
  AND2_X1 U498 ( .A1(n442), .A2(n487), .ZN(n367) );
  BUF_X1 U499 ( .A(n742), .Z(n450) );
  INV_X1 U500 ( .A(n450), .ZN(n454) );
  NOR2_X1 U501 ( .A1(n450), .A2(n490), .ZN(n369) );
  XOR2_X1 U502 ( .A(KEYINPUT46), .B(KEYINPUT92), .Z(n370) );
  XNOR2_X1 U503 ( .A(KEYINPUT88), .B(KEYINPUT45), .ZN(n667) );
  XOR2_X1 U504 ( .A(n678), .B(n677), .Z(n371) );
  XOR2_X1 U505 ( .A(n694), .B(n693), .Z(n372) );
  NAND2_X1 U506 ( .A1(n604), .A2(n373), .ZN(n377) );
  NOR2_X1 U507 ( .A1(n374), .A2(n605), .ZN(n373) );
  INV_X1 U508 ( .A(n717), .ZN(n374) );
  XNOR2_X2 U509 ( .A(n507), .B(n506), .ZN(n686) );
  INV_X1 U510 ( .A(n442), .ZN(n379) );
  XNOR2_X1 U511 ( .A(n508), .B(G472), .ZN(n380) );
  BUF_X1 U512 ( .A(n775), .Z(n381) );
  BUF_X1 U513 ( .A(n692), .Z(n382) );
  INV_X1 U514 ( .A(n816), .ZN(n390) );
  BUF_X1 U515 ( .A(n557), .Z(n383) );
  XNOR2_X1 U516 ( .A(n511), .B(KEYINPUT30), .ZN(n542) );
  NOR2_X1 U517 ( .A1(n692), .A2(G902), .ZN(n384) );
  XNOR2_X1 U518 ( .A(n599), .B(KEYINPUT1), .ZN(n742) );
  BUF_X1 U519 ( .A(n361), .Z(n786) );
  AND2_X1 U520 ( .A1(n385), .A2(n364), .ZN(n674) );
  INV_X1 U521 ( .A(n370), .ZN(n394) );
  XNOR2_X1 U522 ( .A(n386), .B(n669), .ZN(n401) );
  NAND2_X1 U523 ( .A1(n402), .A2(n403), .ZN(n386) );
  NAND2_X1 U524 ( .A1(n387), .A2(n397), .ZN(n406) );
  NOR2_X1 U525 ( .A1(n391), .A2(n395), .ZN(n387) );
  NAND2_X1 U526 ( .A1(n419), .A2(n818), .ZN(n399) );
  AND2_X1 U527 ( .A1(n609), .A2(n588), .ZN(n389) );
  NAND2_X1 U528 ( .A1(n390), .A2(n370), .ZN(n396) );
  NAND2_X1 U529 ( .A1(n817), .A2(n394), .ZN(n393) );
  XNOR2_X2 U530 ( .A(n405), .B(n611), .ZN(n817) );
  NAND2_X1 U531 ( .A1(n393), .A2(n392), .ZN(n391) );
  NAND2_X1 U532 ( .A1(n816), .A2(n394), .ZN(n392) );
  NOR2_X1 U533 ( .A1(n817), .A2(n396), .ZN(n395) );
  NOR2_X1 U534 ( .A1(n400), .A2(n398), .ZN(n397) );
  NAND2_X1 U535 ( .A1(n401), .A2(n671), .ZN(n488) );
  AND2_X2 U536 ( .A1(n488), .A2(n732), .ZN(n782) );
  INV_X2 U537 ( .A(G146), .ZN(n518) );
  INV_X1 U538 ( .A(n404), .ZN(n644) );
  NOR2_X1 U539 ( .A1(n815), .A2(n643), .ZN(n404) );
  NAND2_X1 U540 ( .A1(n407), .A2(n717), .ZN(n405) );
  XNOR2_X1 U541 ( .A(n406), .B(n486), .ZN(n439) );
  XNOR2_X1 U542 ( .A(n603), .B(KEYINPUT106), .ZN(n604) );
  NAND2_X1 U543 ( .A1(n407), .A2(n719), .ZN(n727) );
  XNOR2_X2 U544 ( .A(n417), .B(n610), .ZN(n407) );
  NAND2_X1 U545 ( .A1(n458), .A2(n460), .ZN(n408) );
  NAND2_X1 U546 ( .A1(n411), .A2(n668), .ZN(n410) );
  NAND2_X1 U547 ( .A1(n413), .A2(n458), .ZN(n412) );
  AND2_X1 U548 ( .A1(n460), .A2(n668), .ZN(n413) );
  XNOR2_X2 U549 ( .A(n518), .B(G125), .ZN(n575) );
  XNOR2_X2 U550 ( .A(n617), .B(n616), .ZN(n816) );
  XNOR2_X1 U551 ( .A(n435), .B(n434), .ZN(n609) );
  NAND2_X1 U552 ( .A1(n437), .A2(n436), .ZN(n435) );
  NAND2_X1 U553 ( .A1(n609), .A2(n752), .ZN(n417) );
  NAND2_X1 U554 ( .A1(n598), .A2(KEYINPUT47), .ZN(n419) );
  XNOR2_X1 U555 ( .A(n422), .B(n421), .ZN(n592) );
  NOR2_X1 U556 ( .A1(n589), .A2(n590), .ZN(n422) );
  OR2_X2 U557 ( .A1(n775), .A2(n668), .ZN(n586) );
  XNOR2_X1 U558 ( .A(n726), .B(n453), .ZN(n608) );
  NOR2_X1 U559 ( .A1(n426), .A2(n654), .ZN(n625) );
  XNOR2_X1 U560 ( .A(n645), .B(KEYINPUT104), .ZN(n426) );
  XNOR2_X2 U561 ( .A(n427), .B(KEYINPUT35), .ZN(n815) );
  NAND2_X1 U562 ( .A1(n663), .A2(n366), .ZN(n457) );
  NAND2_X1 U563 ( .A1(n430), .A2(n428), .ZN(n437) );
  NAND2_X1 U564 ( .A1(n442), .A2(n429), .ZN(n428) );
  AND2_X1 U565 ( .A1(n441), .A2(n433), .ZN(n429) );
  NOR2_X1 U566 ( .A1(n432), .A2(n431), .ZN(n430) );
  INV_X1 U567 ( .A(n542), .ZN(n436) );
  NAND2_X1 U568 ( .A1(n439), .A2(n697), .ZN(n438) );
  NOR2_X1 U569 ( .A1(n591), .A2(n368), .ZN(n441) );
  INV_X1 U570 ( .A(n599), .ZN(n442) );
  OR2_X1 U571 ( .A1(n734), .A2(n448), .ZN(n447) );
  XNOR2_X1 U572 ( .A(n625), .B(n624), .ZN(n734) );
  NAND2_X1 U573 ( .A1(n734), .A2(KEYINPUT34), .ZN(n444) );
  NAND2_X1 U574 ( .A1(n706), .A2(n449), .ZN(n448) );
  INV_X1 U575 ( .A(KEYINPUT34), .ZN(n449) );
  NOR2_X1 U576 ( .A1(n742), .A2(n741), .ZN(n623) );
  AND2_X1 U577 ( .A1(n450), .A2(n491), .ZN(n639) );
  XNOR2_X1 U578 ( .A(n451), .B(KEYINPUT123), .ZN(G54) );
  NAND2_X1 U579 ( .A1(n452), .A2(n681), .ZN(n451) );
  XNOR2_X1 U580 ( .A(n695), .B(n372), .ZN(n452) );
  XNOR2_X2 U581 ( .A(n455), .B(G122), .ZN(n567) );
  NAND2_X1 U582 ( .A1(n663), .A2(n664), .ZN(n464) );
  NAND2_X1 U583 ( .A1(n457), .A2(n456), .ZN(n458) );
  INV_X1 U584 ( .A(n667), .ZN(n459) );
  INV_X1 U585 ( .A(n465), .ZN(n460) );
  NAND2_X1 U586 ( .A1(n464), .A2(n462), .ZN(n461) );
  AND2_X1 U587 ( .A1(n666), .A2(n667), .ZN(n462) );
  NAND2_X1 U588 ( .A1(n465), .A2(n667), .ZN(n463) );
  NAND2_X1 U589 ( .A1(n644), .A2(KEYINPUT44), .ZN(n466) );
  NAND2_X1 U590 ( .A1(n481), .A2(n480), .ZN(n479) );
  NAND2_X1 U591 ( .A1(n481), .A2(n467), .ZN(n470) );
  NAND2_X1 U592 ( .A1(n482), .A2(n479), .ZN(n631) );
  INV_X1 U593 ( .A(n474), .ZN(n473) );
  NAND2_X1 U594 ( .A1(n478), .A2(n482), .ZN(n477) );
  AND2_X1 U595 ( .A1(n479), .A2(n632), .ZN(n478) );
  NAND2_X1 U596 ( .A1(n481), .A2(n751), .ZN(n605) );
  INV_X1 U597 ( .A(n621), .ZN(n481) );
  NAND2_X1 U598 ( .A1(n621), .A2(KEYINPUT19), .ZN(n484) );
  XNOR2_X2 U599 ( .A(n485), .B(n638), .ZN(n700) );
  XNOR2_X2 U600 ( .A(n637), .B(n636), .ZN(n657) );
  XNOR2_X1 U601 ( .A(n528), .B(G104), .ZN(n489) );
  XNOR2_X1 U602 ( .A(n489), .B(n535), .ZN(n692) );
  INV_X1 U603 ( .A(n380), .ZN(n491) );
  XOR2_X1 U604 ( .A(n570), .B(n562), .Z(n492) );
  XNOR2_X1 U605 ( .A(n531), .B(n493), .ZN(n532) );
  XNOR2_X1 U606 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U607 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U608 ( .A(n502), .B(n501), .ZN(n505) );
  BUF_X1 U609 ( .A(n734), .Z(n761) );
  XNOR2_X1 U610 ( .A(n563), .B(n492), .ZN(n564) );
  XNOR2_X1 U611 ( .A(n524), .B(n523), .ZN(n591) );
  INV_X1 U612 ( .A(n791), .ZN(n681) );
  INV_X1 U613 ( .A(KEYINPUT63), .ZN(n690) );
  INV_X1 U614 ( .A(KEYINPUT60), .ZN(n683) );
  INV_X2 U615 ( .A(G143), .ZN(n494) );
  XNOR2_X2 U616 ( .A(n494), .B(G128), .ZN(n557) );
  XNOR2_X2 U617 ( .A(n557), .B(n495), .ZN(n577) );
  XNOR2_X2 U618 ( .A(KEYINPUT68), .B(G131), .ZN(n550) );
  NAND2_X1 U619 ( .A1(n543), .A2(G210), .ZN(n497) );
  XNOR2_X1 U620 ( .A(n498), .B(n497), .ZN(n502) );
  XNOR2_X1 U621 ( .A(n503), .B(G101), .ZN(n568) );
  INV_X1 U622 ( .A(n568), .ZN(n504) );
  XNOR2_X1 U623 ( .A(n505), .B(n504), .ZN(n506) );
  NAND2_X1 U624 ( .A1(n510), .A2(n509), .ZN(n584) );
  NAND2_X1 U625 ( .A1(n584), .A2(G214), .ZN(n751) );
  NAND2_X1 U626 ( .A1(n380), .A2(n751), .ZN(n511) );
  NAND2_X1 U627 ( .A1(n558), .A2(G221), .ZN(n515) );
  XOR2_X1 U628 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n513) );
  XNOR2_X1 U629 ( .A(G128), .B(KEYINPUT71), .ZN(n512) );
  XNOR2_X1 U630 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U631 ( .A(n698), .B(G110), .ZN(n571) );
  XOR2_X1 U632 ( .A(n571), .B(KEYINPUT97), .Z(n516) );
  XOR2_X1 U633 ( .A(G137), .B(G140), .Z(n531) );
  XNOR2_X1 U634 ( .A(n531), .B(n554), .ZN(n803) );
  XNOR2_X1 U635 ( .A(n519), .B(n803), .ZN(n787) );
  NOR2_X1 U636 ( .A1(n787), .A2(G902), .ZN(n524) );
  XOR2_X1 U637 ( .A(KEYINPUT25), .B(KEYINPUT80), .Z(n522) );
  NAND2_X1 U638 ( .A1(n670), .A2(G234), .ZN(n520) );
  XNOR2_X1 U639 ( .A(n520), .B(KEYINPUT20), .ZN(n525) );
  NAND2_X1 U640 ( .A1(G217), .A2(n525), .ZN(n521) );
  XNOR2_X1 U641 ( .A(n522), .B(n521), .ZN(n523) );
  AND2_X1 U642 ( .A1(n525), .A2(G221), .ZN(n527) );
  INV_X1 U643 ( .A(KEYINPUT21), .ZN(n526) );
  XNOR2_X1 U644 ( .A(n527), .B(n526), .ZN(n590) );
  INV_X1 U645 ( .A(n590), .ZN(n738) );
  XNOR2_X1 U646 ( .A(n530), .B(n529), .ZN(n533) );
  XOR2_X1 U647 ( .A(n534), .B(KEYINPUT76), .Z(n535) );
  XNOR2_X1 U648 ( .A(KEYINPUT70), .B(G469), .ZN(n536) );
  NAND2_X1 U649 ( .A1(G234), .A2(G237), .ZN(n537) );
  NAND2_X1 U650 ( .A1(G952), .A2(n538), .ZN(n768) );
  NOR2_X1 U651 ( .A1(n768), .A2(n812), .ZN(n626) );
  AND2_X1 U652 ( .A1(n538), .A2(n812), .ZN(n539) );
  NAND2_X1 U653 ( .A1(G902), .A2(n539), .ZN(n627) );
  XOR2_X1 U654 ( .A(KEYINPUT105), .B(n627), .Z(n540) );
  NOR2_X1 U655 ( .A1(G900), .A2(n540), .ZN(n541) );
  NOR2_X1 U656 ( .A1(n626), .A2(n541), .ZN(n589) );
  NAND2_X1 U657 ( .A1(G214), .A2(n543), .ZN(n544) );
  XNOR2_X1 U658 ( .A(n545), .B(n544), .ZN(n549) );
  XNOR2_X1 U659 ( .A(n819), .B(G113), .ZN(n546) );
  XNOR2_X1 U660 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U661 ( .A(n549), .B(n548), .Z(n553) );
  INV_X1 U662 ( .A(n550), .ZN(n551) );
  XNOR2_X1 U663 ( .A(n551), .B(n567), .ZN(n552) );
  NOR2_X1 U664 ( .A1(G902), .A2(n678), .ZN(n556) );
  XNOR2_X1 U665 ( .A(KEYINPUT13), .B(G475), .ZN(n555) );
  XNOR2_X1 U666 ( .A(n556), .B(n555), .ZN(n613) );
  XNOR2_X1 U667 ( .A(n383), .B(KEYINPUT7), .ZN(n565) );
  NAND2_X1 U668 ( .A1(G217), .A2(n558), .ZN(n559) );
  XNOR2_X1 U669 ( .A(n560), .B(n559), .ZN(n563) );
  XNOR2_X1 U670 ( .A(n561), .B(G107), .ZN(n570) );
  XNOR2_X1 U671 ( .A(n565), .B(n564), .ZN(n783) );
  XNOR2_X1 U672 ( .A(G478), .B(n363), .ZN(n612) );
  AND2_X1 U673 ( .A1(n613), .A2(n612), .ZN(n633) );
  INV_X1 U674 ( .A(n633), .ZN(n587) );
  XNOR2_X1 U675 ( .A(n567), .B(n566), .ZN(n569) );
  XNOR2_X1 U676 ( .A(n569), .B(n568), .ZN(n573) );
  XNOR2_X1 U677 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U678 ( .A(n573), .B(n572), .ZN(n796) );
  XNOR2_X1 U679 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U680 ( .A(n577), .B(n576), .ZN(n582) );
  NAND2_X1 U681 ( .A1(G224), .A2(n806), .ZN(n578) );
  XNOR2_X1 U682 ( .A(n578), .B(KEYINPUT82), .ZN(n579) );
  XNOR2_X1 U683 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U684 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U685 ( .A(n796), .B(n583), .ZN(n775) );
  INV_X1 U686 ( .A(n670), .ZN(n668) );
  NAND2_X1 U687 ( .A1(n584), .A2(G210), .ZN(n585) );
  XNOR2_X2 U688 ( .A(n586), .B(n585), .ZN(n621) );
  NOR2_X1 U689 ( .A1(n587), .A2(n621), .ZN(n588) );
  NAND2_X1 U690 ( .A1(n592), .A2(n591), .ZN(n602) );
  NOR2_X1 U691 ( .A1(n491), .A2(n602), .ZN(n593) );
  XOR2_X1 U692 ( .A(KEYINPUT28), .B(n593), .Z(n594) );
  INV_X1 U693 ( .A(n751), .ZN(n595) );
  AND2_X1 U694 ( .A1(n615), .A2(n631), .ZN(n714) );
  INV_X1 U695 ( .A(n612), .ZN(n596) );
  OR2_X1 U696 ( .A1(n613), .A2(n596), .ZN(n703) );
  INV_X2 U697 ( .A(n703), .ZN(n719) );
  AND2_X1 U698 ( .A1(n613), .A2(n596), .ZN(n717) );
  NOR2_X1 U699 ( .A1(n719), .A2(n717), .ZN(n597) );
  NAND2_X1 U700 ( .A1(n714), .A2(n755), .ZN(n598) );
  INV_X1 U701 ( .A(KEYINPUT103), .ZN(n600) );
  XNOR2_X1 U702 ( .A(n600), .B(KEYINPUT6), .ZN(n601) );
  NOR2_X1 U703 ( .A1(n654), .A2(n602), .ZN(n603) );
  NAND2_X1 U704 ( .A1(n714), .A2(n650), .ZN(n606) );
  NOR2_X1 U705 ( .A1(KEYINPUT47), .A2(n606), .ZN(n607) );
  XOR2_X1 U706 ( .A(KEYINPUT73), .B(KEYINPUT39), .Z(n610) );
  XOR2_X1 U707 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n617) );
  OR2_X1 U708 ( .A1(n613), .A2(n612), .ZN(n754) );
  NAND2_X1 U709 ( .A1(n752), .A2(n751), .ZN(n756) );
  NAND2_X1 U710 ( .A1(n365), .A2(n751), .ZN(n618) );
  XNOR2_X1 U711 ( .A(KEYINPUT43), .B(KEYINPUT107), .ZN(n619) );
  XNOR2_X1 U712 ( .A(n620), .B(n619), .ZN(n622) );
  NAND2_X1 U713 ( .A1(n622), .A2(n621), .ZN(n697) );
  XNOR2_X1 U714 ( .A(n623), .B(KEYINPUT75), .ZN(n645) );
  XNOR2_X1 U715 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n624) );
  INV_X1 U716 ( .A(n626), .ZN(n629) );
  OR2_X1 U717 ( .A1(n627), .A2(G898), .ZN(n628) );
  NAND2_X1 U718 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U719 ( .A(KEYINPUT66), .B(KEYINPUT0), .ZN(n632) );
  INV_X1 U720 ( .A(n754), .ZN(n634) );
  NAND2_X1 U721 ( .A1(n634), .A2(n738), .ZN(n635) );
  INV_X1 U722 ( .A(KEYINPUT22), .ZN(n636) );
  XNOR2_X1 U723 ( .A(KEYINPUT64), .B(KEYINPUT32), .ZN(n638) );
  INV_X1 U724 ( .A(KEYINPUT67), .ZN(n661) );
  NAND2_X1 U725 ( .A1(n700), .A2(n661), .ZN(n642) );
  NAND2_X1 U726 ( .A1(n657), .A2(n639), .ZN(n640) );
  XNOR2_X1 U727 ( .A(n640), .B(KEYINPUT65), .ZN(n641) );
  AND2_X1 U728 ( .A1(n641), .A2(n653), .ZN(n710) );
  NOR2_X1 U729 ( .A1(n491), .A2(n645), .ZN(n747) );
  INV_X1 U730 ( .A(n418), .ZN(n706) );
  AND2_X1 U731 ( .A1(n747), .A2(n706), .ZN(n647) );
  INV_X1 U732 ( .A(KEYINPUT31), .ZN(n646) );
  XNOR2_X1 U733 ( .A(n647), .B(n646), .ZN(n720) );
  NAND2_X1 U734 ( .A1(n367), .A2(n491), .ZN(n704) );
  NOR2_X1 U735 ( .A1(n418), .A2(n704), .ZN(n649) );
  OR2_X1 U736 ( .A1(n720), .A2(n649), .ZN(n651) );
  NAND2_X1 U737 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U738 ( .A(n652), .B(KEYINPUT102), .ZN(n658) );
  AND2_X1 U739 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U740 ( .A1(n657), .A2(n656), .ZN(n696) );
  AND2_X1 U741 ( .A1(n658), .A2(n696), .ZN(n659) );
  NAND2_X1 U742 ( .A1(n815), .A2(KEYINPUT67), .ZN(n664) );
  INV_X1 U743 ( .A(KEYINPUT44), .ZN(n660) );
  NAND2_X1 U744 ( .A1(n661), .A2(n660), .ZN(n662) );
  OR2_X1 U745 ( .A1(n815), .A2(n662), .ZN(n663) );
  INV_X1 U746 ( .A(n700), .ZN(n665) );
  NOR2_X1 U747 ( .A1(n710), .A2(n665), .ZN(n666) );
  INV_X1 U748 ( .A(KEYINPUT87), .ZN(n669) );
  INV_X1 U749 ( .A(KEYINPUT2), .ZN(n728) );
  OR2_X1 U750 ( .A1(n670), .A2(n728), .ZN(n671) );
  NAND2_X1 U751 ( .A1(KEYINPUT2), .A2(n727), .ZN(n672) );
  INV_X1 U752 ( .A(KEYINPUT89), .ZN(n673) );
  XNOR2_X1 U753 ( .A(n674), .B(n673), .ZN(n676) );
  NAND2_X1 U754 ( .A1(n676), .A2(n675), .ZN(n732) );
  NAND2_X1 U755 ( .A1(n361), .A2(G475), .ZN(n679) );
  XOR2_X1 U756 ( .A(KEYINPUT59), .B(KEYINPUT94), .Z(n677) );
  XNOR2_X1 U757 ( .A(n679), .B(n371), .ZN(n682) );
  INV_X1 U758 ( .A(G952), .ZN(n680) );
  AND2_X1 U759 ( .A1(n680), .A2(n812), .ZN(n791) );
  NAND2_X1 U760 ( .A1(n682), .A2(n681), .ZN(n684) );
  XNOR2_X1 U761 ( .A(n684), .B(n683), .ZN(G60) );
  NAND2_X1 U762 ( .A1(n782), .A2(G472), .ZN(n688) );
  XNOR2_X1 U763 ( .A(KEYINPUT111), .B(KEYINPUT62), .ZN(n685) );
  XNOR2_X1 U764 ( .A(n688), .B(n687), .ZN(n689) );
  NOR2_X2 U765 ( .A1(n689), .A2(n791), .ZN(n691) );
  XNOR2_X1 U766 ( .A(n691), .B(n690), .ZN(G57) );
  NAND2_X1 U767 ( .A1(n361), .A2(G469), .ZN(n695) );
  XOR2_X1 U768 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n694) );
  XNOR2_X1 U769 ( .A(n382), .B(KEYINPUT122), .ZN(n693) );
  XNOR2_X1 U770 ( .A(n696), .B(G101), .ZN(G3) );
  XNOR2_X1 U771 ( .A(n697), .B(G140), .ZN(G42) );
  XNOR2_X1 U772 ( .A(n698), .B(KEYINPUT127), .ZN(n699) );
  XNOR2_X1 U773 ( .A(n700), .B(n699), .ZN(G21) );
  NOR2_X1 U774 ( .A1(n704), .A2(n374), .ZN(n701) );
  NAND2_X1 U775 ( .A1(n706), .A2(n701), .ZN(n702) );
  XNOR2_X1 U776 ( .A(n702), .B(G104), .ZN(G6) );
  XOR2_X1 U777 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n708) );
  NOR2_X1 U778 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U779 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U780 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X1 U781 ( .A(G107), .B(n709), .ZN(G9) );
  XOR2_X1 U782 ( .A(G110), .B(n710), .Z(G12) );
  XOR2_X1 U783 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n712) );
  NAND2_X1 U784 ( .A1(n714), .A2(n719), .ZN(n711) );
  XNOR2_X1 U785 ( .A(n712), .B(n711), .ZN(n713) );
  XNOR2_X1 U786 ( .A(G128), .B(n713), .ZN(G30) );
  NAND2_X1 U787 ( .A1(n714), .A2(n717), .ZN(n715) );
  XNOR2_X1 U788 ( .A(n715), .B(KEYINPUT114), .ZN(n716) );
  XNOR2_X1 U789 ( .A(G146), .B(n716), .ZN(G48) );
  NAND2_X1 U790 ( .A1(n720), .A2(n717), .ZN(n718) );
  XNOR2_X1 U791 ( .A(n718), .B(G113), .ZN(G15) );
  XOR2_X1 U792 ( .A(G116), .B(KEYINPUT115), .Z(n722) );
  NAND2_X1 U793 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U794 ( .A(n722), .B(n721), .ZN(G18) );
  XOR2_X1 U795 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n724) );
  XNOR2_X1 U796 ( .A(G125), .B(KEYINPUT37), .ZN(n723) );
  XNOR2_X1 U797 ( .A(n724), .B(n723), .ZN(n725) );
  XNOR2_X1 U798 ( .A(n726), .B(n725), .ZN(G27) );
  XNOR2_X1 U799 ( .A(G134), .B(n727), .ZN(G36) );
  NAND2_X1 U800 ( .A1(n356), .A2(n728), .ZN(n729) );
  XNOR2_X1 U801 ( .A(n729), .B(KEYINPUT86), .ZN(n731) );
  OR2_X1 U802 ( .A1(n675), .A2(KEYINPUT2), .ZN(n730) );
  AND2_X1 U803 ( .A1(n731), .A2(n730), .ZN(n733) );
  AND2_X1 U804 ( .A1(n733), .A2(n732), .ZN(n737) );
  INV_X1 U805 ( .A(n749), .ZN(n735) );
  NOR2_X1 U806 ( .A1(n761), .A2(n735), .ZN(n736) );
  NOR2_X1 U807 ( .A1(n737), .A2(n736), .ZN(n771) );
  XNOR2_X1 U808 ( .A(KEYINPUT119), .B(KEYINPUT52), .ZN(n766) );
  NOR2_X1 U809 ( .A1(n490), .A2(n738), .ZN(n739) );
  XNOR2_X1 U810 ( .A(n739), .B(KEYINPUT49), .ZN(n740) );
  NAND2_X1 U811 ( .A1(n491), .A2(n740), .ZN(n745) );
  NAND2_X1 U812 ( .A1(n450), .A2(n741), .ZN(n743) );
  XOR2_X1 U813 ( .A(KEYINPUT50), .B(n743), .Z(n744) );
  NOR2_X1 U814 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U815 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U816 ( .A(KEYINPUT51), .B(n748), .ZN(n750) );
  NAND2_X1 U817 ( .A1(n750), .A2(n749), .ZN(n764) );
  NOR2_X1 U818 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U819 ( .A1(n754), .A2(n753), .ZN(n759) );
  INV_X1 U820 ( .A(n755), .ZN(n757) );
  NOR2_X1 U821 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U822 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U823 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U824 ( .A(KEYINPUT118), .B(n762), .Z(n763) );
  NAND2_X1 U825 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U826 ( .A(n766), .B(n765), .ZN(n767) );
  NOR2_X1 U827 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U828 ( .A(KEYINPUT120), .B(n769), .Z(n770) );
  NAND2_X1 U829 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U830 ( .A(n773), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U831 ( .A1(n782), .A2(G210), .ZN(n777) );
  XOR2_X1 U832 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n774) );
  XNOR2_X1 U833 ( .A(n777), .B(n776), .ZN(n778) );
  NOR2_X2 U834 ( .A1(n778), .A2(n791), .ZN(n781) );
  XNOR2_X1 U835 ( .A(KEYINPUT121), .B(KEYINPUT56), .ZN(n779) );
  XNOR2_X1 U836 ( .A(n779), .B(KEYINPUT91), .ZN(n780) );
  XNOR2_X1 U837 ( .A(n781), .B(n780), .ZN(G51) );
  NAND2_X1 U838 ( .A1(n786), .A2(G478), .ZN(n784) );
  XNOR2_X1 U839 ( .A(n784), .B(n783), .ZN(n785) );
  NOR2_X1 U840 ( .A1(n791), .A2(n785), .ZN(G63) );
  NAND2_X1 U841 ( .A1(n786), .A2(G217), .ZN(n789) );
  XNOR2_X1 U842 ( .A(n787), .B(KEYINPUT124), .ZN(n788) );
  XNOR2_X1 U843 ( .A(n789), .B(n788), .ZN(n790) );
  NOR2_X1 U844 ( .A1(n791), .A2(n790), .ZN(G66) );
  NAND2_X1 U845 ( .A1(n675), .A2(n806), .ZN(n795) );
  NAND2_X1 U846 ( .A1(n812), .A2(G224), .ZN(n792) );
  XNOR2_X1 U847 ( .A(KEYINPUT61), .B(n792), .ZN(n793) );
  NAND2_X1 U848 ( .A1(n793), .A2(G898), .ZN(n794) );
  NAND2_X1 U849 ( .A1(n795), .A2(n794), .ZN(n800) );
  INV_X1 U850 ( .A(n796), .ZN(n798) );
  NOR2_X1 U851 ( .A1(G898), .A2(n806), .ZN(n797) );
  NOR2_X1 U852 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U853 ( .A(n800), .B(n799), .ZN(n801) );
  XOR2_X1 U854 ( .A(KEYINPUT125), .B(n801), .Z(G69) );
  BUF_X1 U855 ( .A(n802), .Z(n804) );
  XNOR2_X1 U856 ( .A(n804), .B(n803), .ZN(n808) );
  XNOR2_X1 U857 ( .A(n356), .B(n808), .ZN(n807) );
  NAND2_X1 U858 ( .A1(n807), .A2(n806), .ZN(n814) );
  XNOR2_X1 U859 ( .A(G227), .B(n808), .ZN(n809) );
  NAND2_X1 U860 ( .A1(n809), .A2(G900), .ZN(n810) );
  XNOR2_X1 U861 ( .A(KEYINPUT126), .B(n810), .ZN(n811) );
  NAND2_X1 U862 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U863 ( .A1(n814), .A2(n813), .ZN(G72) );
  XOR2_X1 U864 ( .A(n815), .B(G122), .Z(G24) );
  XOR2_X1 U865 ( .A(G137), .B(n816), .Z(G39) );
  XOR2_X1 U866 ( .A(n817), .B(G131), .Z(G33) );
  XOR2_X1 U867 ( .A(n819), .B(n818), .Z(n820) );
  XNOR2_X1 U868 ( .A(KEYINPUT113), .B(n820), .ZN(G45) );
endmodule

