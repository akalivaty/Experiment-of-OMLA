//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 0 1 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT64), .B(G20), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n201), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n212), .B1(new_n216), .B2(new_n218), .C1(new_n227), .C2(KEYINPUT1), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n202), .A2(G68), .ZN(new_n242));
  INV_X1    g0042(.A(G68), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n241), .B(new_n247), .ZN(G351));
  NAND2_X1  g0048(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT64), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT3), .B(G33), .ZN(new_n253));
  OAI21_X1  g0053(.A(KEYINPUT7), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT7), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(new_n258), .A3(new_n207), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n254), .A2(G68), .A3(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(G58), .A2(G68), .ZN(new_n261));
  OAI21_X1  g0061(.A(G20), .B1(new_n261), .B2(new_n201), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G159), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT16), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n214), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  OR2_X1    g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(new_n207), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n243), .B1(new_n275), .B2(KEYINPUT7), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n257), .A2(new_n213), .A3(new_n258), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n265), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n272), .B1(new_n278), .B2(KEYINPUT16), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n269), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G200), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G1), .A3(G13), .ZN(new_n283));
  INV_X1    g0083(.A(G223), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G226), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G1698), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n286), .B(new_n288), .C1(new_n255), .C2(new_n256), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G87), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n283), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n283), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G274), .ZN(new_n296));
  INV_X1    g0096(.A(new_n214), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n296), .B1(new_n297), .B2(new_n282), .ZN(new_n298));
  INV_X1    g0098(.A(new_n293), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n295), .A2(G232), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n281), .B1(new_n292), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G232), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n283), .A2(G274), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n302), .A2(new_n294), .B1(new_n303), .B2(new_n293), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n304), .A2(new_n291), .A3(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g0107(.A(KEYINPUT8), .B(G58), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(new_n206), .B2(G20), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(new_n271), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n309), .A2(new_n312), .B1(new_n308), .B2(new_n311), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n280), .A2(new_n307), .A3(KEYINPUT76), .A4(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT17), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n313), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(new_n269), .B2(new_n279), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n318), .A2(KEYINPUT76), .A3(KEYINPUT17), .A4(new_n307), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G179), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n304), .A2(new_n291), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n292), .A2(new_n300), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(G169), .ZN(new_n324));
  OAI211_X1 g0124(.A(KEYINPUT75), .B(KEYINPUT18), .C1(new_n318), .C2(new_n324), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n255), .A2(new_n256), .A3(G20), .ZN(new_n326));
  OAI21_X1  g0126(.A(G68), .B1(new_n326), .B2(new_n258), .ZN(new_n327));
  NOR3_X1   g0127(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT7), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n266), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n271), .B1(new_n329), .B2(new_n268), .ZN(new_n330));
  AOI21_X1  g0130(.A(KEYINPUT16), .B1(new_n260), .B2(new_n266), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n313), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n323), .A2(G169), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n323), .B2(new_n321), .ZN(new_n334));
  XOR2_X1   g0134(.A(KEYINPUT75), .B(KEYINPUT18), .Z(new_n335));
  NAND3_X1  g0135(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n325), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n320), .A2(new_n337), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n263), .A2(G50), .B1(G20), .B2(new_n243), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n213), .A2(G33), .ZN(new_n340));
  INV_X1    g0140(.A(G77), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n271), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT11), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n343), .B(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n311), .A2(new_n243), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n346), .B(KEYINPUT12), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n206), .A2(G20), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n312), .A2(G68), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT74), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n347), .A2(KEYINPUT74), .A3(new_n349), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n345), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT14), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n302), .A2(G1698), .ZN(new_n357));
  OAI221_X1 g0157(.A(new_n357), .B1(G226), .B2(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G97), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT73), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n283), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n358), .A2(KEYINPUT73), .A3(new_n359), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT13), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n298), .A2(new_n299), .ZN(new_n367));
  INV_X1    g0167(.A(G238), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n367), .B1(new_n294), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n365), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n366), .B1(new_n365), .B2(new_n370), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n356), .B(G169), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n365), .A2(new_n370), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT13), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n365), .A2(new_n366), .A3(new_n370), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(G179), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n375), .A2(new_n376), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n356), .B1(new_n379), .B2(G169), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n355), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(G200), .B1(new_n371), .B2(new_n372), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n375), .A2(G190), .A3(new_n376), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n354), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n253), .A2(G232), .A3(new_n285), .ZN(new_n386));
  INV_X1    g0186(.A(G107), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n253), .A2(G1698), .ZN(new_n388));
  OAI221_X1 g0188(.A(new_n386), .B1(new_n387), .B2(new_n253), .C1(new_n388), .C2(new_n368), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n363), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n295), .A2(G244), .B1(new_n298), .B2(new_n299), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(G190), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT69), .ZN(new_n393));
  XNOR2_X1  g0193(.A(new_n392), .B(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT71), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n348), .A2(G77), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n312), .A2(new_n397), .B1(new_n341), .B2(new_n311), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT70), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n308), .B(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n263), .ZN(new_n401));
  INV_X1    g0201(.A(new_n340), .ZN(new_n402));
  XNOR2_X1  g0202(.A(KEYINPUT15), .B(G87), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n402), .A2(new_n404), .B1(G77), .B2(new_n252), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n395), .B(new_n398), .C1(new_n406), .C2(new_n272), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n272), .B1(new_n401), .B2(new_n405), .ZN(new_n408));
  INV_X1    g0208(.A(new_n398), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT71), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n390), .A2(new_n391), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G200), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n407), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n411), .A2(G179), .ZN(new_n414));
  INV_X1    g0214(.A(G169), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(new_n411), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n407), .A2(new_n410), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n394), .A2(new_n413), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n338), .A2(new_n381), .A3(new_n385), .A4(new_n418), .ZN(new_n419));
  OAI211_X1 g0219(.A(G222), .B(new_n285), .C1(new_n255), .C2(new_n256), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT67), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n420), .B(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n257), .A2(new_n285), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n423), .A2(G223), .B1(new_n257), .B2(G77), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n283), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n367), .B1(new_n294), .B2(new_n287), .ZN(new_n426));
  NOR3_X1   g0226(.A1(new_n425), .A2(KEYINPUT68), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT68), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n420), .B(KEYINPUT67), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n388), .A2(new_n284), .B1(new_n341), .B2(new_n253), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n363), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n426), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n428), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(G190), .B1(new_n427), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n308), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n402), .A2(new_n435), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n263), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n271), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n202), .B1(new_n206), .B2(G20), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n312), .A2(new_n440), .B1(new_n202), .B2(new_n311), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(KEYINPUT9), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT9), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n272), .B1(new_n436), .B2(new_n437), .ZN(new_n444));
  INV_X1    g0244(.A(new_n441), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT68), .B1(new_n425), .B2(new_n426), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n431), .A2(new_n428), .A3(new_n432), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n449), .A2(new_n450), .A3(G200), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n434), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT72), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n434), .A2(new_n448), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT10), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n452), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n449), .A2(new_n450), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n447), .B1(new_n457), .B2(G190), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n458), .B(new_n451), .C1(new_n453), .C2(KEYINPUT10), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n321), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n439), .A2(new_n441), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n460), .B(new_n461), .C1(G169), .C2(new_n457), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n456), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n419), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n253), .A2(G257), .A3(G1698), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G294), .ZN(new_n467));
  OAI211_X1 g0267(.A(G250), .B(new_n285), .C1(new_n255), .C2(new_n256), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n363), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n206), .A2(G45), .ZN(new_n471));
  OR2_X1    g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  NAND2_X1  g0272(.A1(KEYINPUT5), .A2(G41), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n298), .ZN(new_n475));
  XNOR2_X1  g0275(.A(KEYINPUT5), .B(G41), .ZN(new_n476));
  INV_X1    g0276(.A(new_n471), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n476), .A2(new_n477), .B1(new_n297), .B2(new_n282), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G264), .ZN(new_n479));
  AND4_X1   g0279(.A1(new_n321), .A2(new_n470), .A3(new_n475), .A4(new_n479), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n469), .A2(new_n363), .B1(G264), .B2(new_n478), .ZN(new_n481));
  AOI21_X1  g0281(.A(G169), .B1(new_n481), .B2(new_n475), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n213), .A2(new_n253), .A3(G87), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT22), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT22), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n213), .A2(new_n253), .A3(new_n486), .A4(G87), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(KEYINPUT23), .A2(G107), .ZN(new_n489));
  AOI21_X1  g0289(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(G20), .ZN(new_n491));
  NOR2_X1   g0291(.A1(KEYINPUT23), .A2(G107), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n491), .B1(new_n252), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT24), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT24), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n488), .A2(new_n496), .A3(new_n493), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n272), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n311), .A2(KEYINPUT25), .A3(new_n387), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT25), .B1(new_n311), .B2(new_n387), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n206), .A2(G33), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n310), .A2(new_n502), .A3(new_n214), .A4(new_n270), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n500), .A2(new_n501), .B1(new_n387), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n483), .B1(new_n498), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n497), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n496), .B1(new_n488), .B2(new_n493), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n271), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n481), .A2(G190), .A3(new_n475), .ZN(new_n509));
  INV_X1    g0309(.A(new_n504), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n481), .A2(new_n475), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G200), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n508), .A2(new_n509), .A3(new_n510), .A4(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(G238), .B(new_n285), .C1(new_n255), .C2(new_n256), .ZN(new_n514));
  OAI211_X1 g0314(.A(G244), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G116), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n363), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n471), .A2(G250), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n298), .A2(new_n477), .B1(new_n519), .B2(new_n283), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G190), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT82), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n522), .A2(KEYINPUT82), .A3(G190), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n521), .A2(G200), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n404), .A2(new_n310), .ZN(new_n528));
  INV_X1    g0328(.A(G87), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n503), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n249), .A2(new_n251), .A3(G33), .A4(G97), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT19), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n213), .A2(new_n253), .A3(G68), .ZN(new_n534));
  NAND3_X1  g0334(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n249), .A2(new_n251), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(G97), .A2(G107), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n529), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n533), .A2(new_n534), .A3(new_n539), .ZN(new_n540));
  AOI211_X1 g0340(.A(new_n528), .B(new_n530), .C1(new_n540), .C2(new_n271), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n525), .A2(new_n526), .A3(new_n527), .A4(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n521), .A2(new_n321), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n415), .B1(new_n518), .B2(new_n520), .ZN(new_n544));
  OAI21_X1  g0344(.A(KEYINPUT81), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n521), .A2(G169), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT81), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n546), .B(new_n547), .C1(new_n321), .C2(new_n521), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n540), .A2(new_n271), .ZN(new_n549));
  INV_X1    g0349(.A(new_n528), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n549), .B(new_n550), .C1(new_n403), .C2(new_n503), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n545), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  AND4_X1   g0352(.A1(new_n505), .A2(new_n513), .A3(new_n542), .A4(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT80), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n254), .A2(G107), .A3(new_n259), .ZN(new_n555));
  INV_X1    g0355(.A(new_n263), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(new_n341), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT6), .ZN(new_n558));
  AND2_X1   g0358(.A1(G97), .A2(G107), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(new_n559), .B2(new_n537), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n387), .A2(KEYINPUT6), .A3(G97), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n557), .B1(new_n562), .B2(new_n252), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n272), .B1(new_n555), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n310), .A2(G97), .ZN(new_n565));
  INV_X1    g0365(.A(new_n503), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n565), .B1(new_n566), .B2(G97), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n554), .B1(new_n564), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n258), .B1(new_n257), .B2(new_n213), .ZN(new_n570));
  NOR4_X1   g0370(.A1(new_n255), .A2(new_n256), .A3(KEYINPUT7), .A4(G20), .ZN(new_n571));
  NOR3_X1   g0371(.A1(new_n570), .A2(new_n571), .A3(new_n387), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n387), .A2(KEYINPUT6), .A3(G97), .ZN(new_n573));
  XNOR2_X1  g0373(.A(G97), .B(G107), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n573), .B1(new_n574), .B2(new_n558), .ZN(new_n575));
  OAI22_X1  g0375(.A1(new_n575), .A2(new_n213), .B1(new_n341), .B2(new_n556), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n271), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n577), .A2(KEYINPUT80), .A3(new_n567), .ZN(new_n578));
  OAI211_X1 g0378(.A(G244), .B(new_n285), .C1(new_n255), .C2(new_n256), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT4), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n253), .A2(KEYINPUT4), .A3(G244), .A4(new_n285), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n253), .A2(G250), .A3(G1698), .ZN(new_n583));
  NAND2_X1  g0383(.A1(G33), .A2(G283), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT78), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT78), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(G33), .A3(G283), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n581), .A2(new_n582), .A3(new_n583), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n363), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n476), .A2(new_n477), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n591), .A2(G257), .A3(new_n283), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n475), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G169), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n593), .B1(new_n363), .B2(new_n589), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G179), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n569), .A2(new_n578), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n577), .A2(KEYINPUT77), .A3(new_n567), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT77), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n564), .B2(new_n568), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n590), .A2(new_n594), .A3(new_n305), .ZN(new_n603));
  AOI21_X1  g0403(.A(G200), .B1(new_n590), .B2(new_n594), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n600), .B(new_n602), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT79), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n590), .A2(new_n594), .A3(new_n305), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(G200), .B2(new_n597), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT79), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n608), .A2(new_n609), .A3(new_n602), .A4(new_n600), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n599), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n310), .A2(G116), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n566), .B2(G116), .ZN(new_n613));
  INV_X1    g0413(.A(G116), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n270), .A2(new_n214), .B1(G20), .B2(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n585), .A2(new_n587), .ZN(new_n616));
  INV_X1    g0416(.A(G33), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G97), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n249), .A2(new_n251), .A3(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(KEYINPUT20), .B(new_n615), .C1(new_n616), .C2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n588), .A2(new_n213), .A3(new_n618), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT20), .B1(new_n622), .B2(new_n615), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n613), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n478), .A2(G270), .B1(new_n298), .B2(new_n474), .ZN(new_n625));
  OAI211_X1 g0425(.A(G264), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n626));
  OAI211_X1 g0426(.A(G257), .B(new_n285), .C1(new_n255), .C2(new_n256), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n273), .A2(G303), .A3(new_n274), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n363), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n624), .A2(new_n631), .A3(G179), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n415), .B1(new_n625), .B2(new_n630), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n624), .A2(new_n633), .A3(KEYINPUT21), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT21), .B1(new_n624), .B2(new_n633), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n625), .A2(new_n630), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n624), .B1(G200), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n305), .B2(new_n638), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n553), .A2(new_n611), .A3(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n465), .A2(new_n643), .ZN(G372));
  AND2_X1   g0444(.A1(new_n416), .A2(new_n417), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n385), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n320), .B1(new_n646), .B2(new_n381), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT85), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n332), .A2(new_n648), .A3(new_n334), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT85), .B1(new_n318), .B2(new_n324), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT18), .ZN(new_n651));
  AOI21_X1  g0451(.A(KEYINPUT18), .B1(new_n649), .B2(new_n650), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n459), .B(new_n456), .C1(new_n647), .C2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n462), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n546), .B1(new_n321), .B2(new_n521), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n551), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n498), .A2(new_n504), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n512), .A2(new_n509), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n637), .A2(new_n505), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n611), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT83), .ZN(new_n663));
  INV_X1    g0463(.A(new_n530), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n549), .A2(new_n550), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n281), .B1(new_n518), .B2(new_n520), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n541), .A2(new_n527), .A3(KEYINPUT83), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(new_n668), .A3(new_n523), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT84), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n669), .A2(new_n670), .A3(new_n658), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n670), .B1(new_n669), .B2(new_n658), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n658), .B1(new_n662), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n542), .A2(new_n599), .A3(new_n552), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n602), .A2(new_n600), .B1(new_n596), .B2(new_n598), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n671), .B2(new_n672), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n677), .B1(new_n679), .B2(new_n676), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n464), .B1(new_n674), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n656), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT86), .ZN(G369));
  INV_X1    g0483(.A(new_n637), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n213), .A2(new_n206), .A3(G13), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G213), .A3(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G343), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n691), .A2(new_n624), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n684), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT87), .ZN(new_n694));
  OAI211_X1 g0494(.A(new_n693), .B(new_n694), .C1(new_n641), .C2(new_n692), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n684), .A2(KEYINPUT87), .A3(new_n692), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n505), .A2(new_n513), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n659), .B2(new_n690), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n505), .B2(new_n690), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n505), .A2(new_n691), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n637), .A2(new_n691), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(G399));
  INV_X1    g0506(.A(new_n210), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n538), .A2(G116), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G1), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n218), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n631), .A2(new_n522), .A3(G179), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(new_n595), .A3(new_n511), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n597), .A2(new_n522), .A3(new_n481), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n638), .A2(new_n321), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n716), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n522), .A2(new_n481), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n721), .A2(KEYINPUT30), .A3(new_n597), .A4(new_n718), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n715), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT88), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n723), .A2(new_n691), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT31), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n724), .A2(new_n725), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n726), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n553), .A2(new_n611), .A3(new_n642), .A4(new_n690), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G330), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n690), .B1(new_n674), .B2(new_n680), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT89), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI211_X1 g0539(.A(KEYINPUT89), .B(new_n690), .C1(new_n674), .C2(new_n680), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT29), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI221_X1 g0543(.A(new_n658), .B1(new_n675), .B2(KEYINPUT26), .C1(new_n662), .C2(new_n673), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n679), .A2(KEYINPUT26), .ZN(new_n745));
  OAI211_X1 g0545(.A(KEYINPUT29), .B(new_n690), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n736), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n713), .B1(new_n747), .B2(G1), .ZN(G364));
  NOR2_X1   g0548(.A1(new_n697), .A2(G330), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n213), .A2(G13), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G45), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n709), .A2(G1), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT90), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n698), .A2(new_n749), .A3(new_n753), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT91), .Z(new_n755));
  NOR2_X1   g0555(.A1(new_n707), .A2(new_n257), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n756), .A2(G355), .B1(new_n614), .B2(new_n707), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n707), .A2(new_n253), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(G45), .B2(new_n218), .ZN(new_n759));
  INV_X1    g0559(.A(G45), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n247), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n757), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT92), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n214), .B1(G20), .B2(new_n415), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(new_n762), .B2(new_n763), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n213), .A2(new_n321), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n281), .A2(G190), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G68), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n281), .A2(G179), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n252), .A2(new_n305), .A3(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n387), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n305), .A2(G179), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n213), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G97), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n776), .A2(G20), .A3(G190), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n529), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n257), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n775), .A2(new_n779), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  NOR4_X1   g0587(.A1(new_n213), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G159), .ZN(new_n790));
  OR3_X1    g0590(.A1(new_n789), .A2(KEYINPUT32), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(KEYINPUT32), .B1(new_n789), .B2(new_n790), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n771), .A2(G190), .A3(G200), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n791), .B(new_n792), .C1(new_n202), .C2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G190), .A2(G200), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n771), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(KEYINPUT94), .ZN(new_n798));
  AND3_X1   g0598(.A1(new_n771), .A2(KEYINPUT94), .A3(new_n795), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n787), .B(new_n794), .C1(G77), .C2(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n771), .A2(G190), .A3(new_n281), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT93), .Z(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G58), .ZN(new_n806));
  XOR2_X1   g0606(.A(KEYINPUT33), .B(G317), .Z(new_n807));
  INV_X1    g0607(.A(G283), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n773), .A2(new_n807), .B1(new_n808), .B2(new_n777), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(G329), .B2(new_n788), .ZN(new_n810));
  INV_X1    g0610(.A(new_n793), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G326), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n797), .A2(G311), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n782), .A2(G294), .ZN(new_n814));
  INV_X1    g0614(.A(new_n784), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n253), .B1(new_n815), .B2(G303), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n812), .A2(new_n813), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n803), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(G322), .B2(new_n818), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n802), .A2(new_n806), .B1(new_n810), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n768), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n753), .B1(new_n764), .B2(new_n770), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT95), .ZN(new_n823));
  INV_X1    g0623(.A(new_n767), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n697), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n755), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G396));
  INV_X1    g0627(.A(new_n753), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n811), .A2(G137), .B1(new_n774), .B2(G150), .ZN(new_n829));
  INV_X1    g0629(.A(G143), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n829), .B1(new_n800), .B2(new_n790), .C1(new_n804), .C2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT34), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT96), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n777), .A2(new_n243), .ZN(new_n836));
  INV_X1    g0636(.A(G58), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n253), .B1(new_n202), .B2(new_n784), .C1(new_n781), .C2(new_n837), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n836), .B(new_n838), .C1(G132), .C2(new_n788), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n834), .A2(new_n835), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n801), .A2(G116), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n783), .B(new_n257), .C1(new_n387), .C2(new_n784), .ZN(new_n842));
  INV_X1    g0642(.A(new_n777), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n842), .B1(G87), .B2(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n774), .A2(G283), .B1(G311), .B2(new_n788), .ZN(new_n845));
  AOI22_X1  g0645(.A1(G294), .A2(new_n818), .B1(new_n811), .B2(G303), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n841), .A2(new_n844), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n821), .B1(new_n840), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n768), .A2(new_n765), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n828), .B(new_n848), .C1(new_n341), .C2(new_n849), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n850), .A2(KEYINPUT97), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n850), .A2(KEYINPUT97), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n416), .A2(new_n417), .A3(new_n690), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n690), .B1(new_n407), .B2(new_n410), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n413), .B2(new_n394), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n853), .B1(new_n855), .B2(new_n645), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n857), .A2(new_n766), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n851), .A2(new_n852), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n856), .B(KEYINPUT98), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n741), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n418), .A2(new_n690), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n674), .B2(new_n680), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n753), .B1(new_n866), .B2(new_n735), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n862), .A2(new_n736), .A3(new_n865), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n859), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(G384));
  OR2_X1    g0671(.A1(new_n562), .A2(KEYINPUT35), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n562), .A2(KEYINPUT35), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n872), .A2(new_n873), .A3(G116), .A4(new_n215), .ZN(new_n874));
  XOR2_X1   g0674(.A(new_n874), .B(KEYINPUT36), .Z(new_n875));
  OR3_X1    g0675(.A1(new_n218), .A2(new_n341), .A3(new_n261), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n206), .B(G13), .C1(new_n876), .C2(new_n242), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n329), .A2(new_n268), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n317), .B1(new_n279), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n880), .A2(new_n688), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n320), .B2(new_n337), .ZN(new_n882));
  INV_X1    g0682(.A(new_n307), .ZN(new_n883));
  OAI22_X1  g0683(.A1(new_n332), .A2(new_n883), .B1(new_n880), .B2(new_n688), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n880), .A2(new_n324), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT37), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT37), .B1(new_n332), .B2(new_n334), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n318), .A2(new_n307), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n332), .A2(new_n689), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n882), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT38), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n882), .A2(new_n891), .A3(KEYINPUT38), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(KEYINPUT100), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  AOI211_X1 g0697(.A(KEYINPUT100), .B(KEYINPUT38), .C1(new_n882), .C2(new_n891), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n355), .A2(new_n691), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n381), .A2(new_n385), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(G169), .B1(new_n371), .B2(new_n372), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT14), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(new_n377), .A3(new_n373), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n355), .B(new_n691), .C1(new_n904), .C2(new_n384), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT99), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n865), .A2(new_n907), .A3(new_n853), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n907), .B1(new_n865), .B2(new_n853), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n899), .B(new_n906), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n904), .A2(new_n355), .A3(new_n690), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n898), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n896), .A2(new_n913), .A3(KEYINPUT101), .A4(KEYINPUT39), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n896), .A2(new_n913), .A3(KEYINPUT39), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n316), .A2(new_n319), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n651), .B2(new_n652), .ZN(new_n918));
  INV_X1    g0718(.A(new_n889), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n649), .A2(new_n650), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n889), .A2(new_n888), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT37), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n918), .A2(new_n919), .B1(new_n922), .B2(new_n890), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n916), .B(new_n895), .C1(new_n923), .C2(KEYINPUT38), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT101), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n912), .B(new_n914), .C1(new_n915), .C2(new_n926), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n651), .A2(new_n652), .A3(new_n689), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n910), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n746), .A2(new_n464), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n655), .B1(new_n743), .B2(new_n932), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n930), .B(new_n933), .Z(new_n934));
  AOI21_X1  g0734(.A(new_n856), .B1(new_n901), .B2(new_n905), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n732), .A2(new_n724), .A3(new_n729), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT40), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n937), .A2(new_n938), .A3(new_n913), .A4(new_n896), .ZN(new_n939));
  INV_X1    g0739(.A(new_n895), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n918), .A2(new_n919), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n922), .A2(new_n890), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n940), .B1(new_n943), .B2(new_n893), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n935), .A2(new_n936), .ZN(new_n945));
  OAI21_X1  g0745(.A(KEYINPUT40), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n939), .A2(new_n946), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n464), .A2(new_n936), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n949), .A2(G330), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n934), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n206), .B2(new_n750), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n934), .A2(new_n951), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n878), .B1(new_n953), .B2(new_n954), .ZN(G367));
  NAND2_X1  g0755(.A1(new_n600), .A2(new_n602), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n691), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n611), .A2(new_n957), .B1(new_n678), .B2(new_n691), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(new_n705), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT42), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n958), .A2(new_n505), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n690), .B1(new_n961), .B2(new_n599), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n690), .A2(new_n541), .ZN(new_n964));
  MUX2_X1   g0764(.A(new_n673), .B(new_n658), .S(new_n964), .Z(new_n965));
  XNOR2_X1  g0765(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  MUX2_X1   g0767(.A(KEYINPUT43), .B(new_n966), .S(new_n965), .Z(new_n968));
  OAI21_X1  g0768(.A(new_n967), .B1(new_n963), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT103), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n702), .A2(new_n958), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n967), .B(KEYINPUT103), .C1(new_n963), .C2(new_n968), .ZN(new_n973));
  AND3_X1   g0773(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n972), .B1(new_n971), .B2(new_n973), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n751), .A2(G1), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(KEYINPUT29), .B1(new_n739), .B2(new_n740), .ZN(new_n979));
  INV_X1    g0779(.A(new_n746), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n735), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n705), .A2(new_n703), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT104), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n982), .B(new_n958), .C1(new_n983), .C2(KEYINPUT44), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(KEYINPUT44), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n984), .B(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n982), .A2(new_n958), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT45), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n989), .A2(new_n698), .A3(new_n701), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(new_n702), .A3(new_n988), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT105), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n698), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n705), .B1(new_n701), .B2(new_n704), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n697), .A2(G330), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n996), .B1(new_n997), .B2(KEYINPUT105), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n995), .B(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n981), .B1(new_n993), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n708), .B(KEYINPUT41), .Z(new_n1001));
  OAI21_X1  g0801(.A(new_n978), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n976), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n758), .A2(new_n237), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1004), .B(new_n769), .C1(new_n210), .C2(new_n403), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1005), .A2(KEYINPUT106), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(KEYINPUT106), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1007), .A2(new_n753), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(G150), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n830), .A2(new_n793), .B1(new_n803), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n782), .A2(G68), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n837), .B2(new_n784), .C1(new_n790), .C2(new_n773), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1011), .B(new_n1013), .C1(G137), .C2(new_n788), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n257), .B1(new_n843), .B2(G77), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1015), .A2(KEYINPUT107), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n801), .A2(G50), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(KEYINPUT107), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n805), .A2(G303), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n257), .B1(new_n781), .B2(new_n387), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n784), .A2(new_n614), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT46), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1021), .B(new_n1023), .C1(G311), .C2(new_n811), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n801), .A2(G283), .ZN(new_n1025));
  INV_X1    g0825(.A(G97), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n777), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(G317), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1028), .B1(new_n1029), .B2(new_n789), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G294), .B2(new_n774), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1020), .A2(new_n1024), .A3(new_n1025), .A4(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1019), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT47), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1034), .A2(new_n768), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n1009), .B(new_n1035), .C1(new_n767), .C2(new_n965), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1003), .A2(new_n1037), .ZN(G387));
  XOR2_X1   g0838(.A(new_n995), .B(new_n998), .Z(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n981), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n747), .A2(new_n999), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1040), .A2(new_n1041), .A3(new_n708), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n710), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n756), .A2(new_n1043), .B1(new_n387), .B2(new_n707), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n400), .A2(new_n202), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT50), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n760), .B1(new_n243), .B2(new_n341), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n1046), .A2(new_n1043), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n758), .B1(new_n234), .B2(new_n760), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1044), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n828), .B1(new_n1050), .B2(new_n769), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n701), .B2(new_n824), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(KEYINPUT108), .B(G150), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n789), .A2(new_n1053), .B1(new_n308), .B2(new_n773), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G68), .B2(new_n797), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n782), .A2(new_n404), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n257), .B1(new_n815), .B2(G77), .ZN(new_n1057));
  AND3_X1   g0857(.A1(new_n1028), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n811), .A2(G159), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n818), .A2(G50), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1055), .A2(new_n1058), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(G294), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n781), .A2(new_n808), .B1(new_n1062), .B2(new_n784), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT109), .Z(new_n1064));
  INV_X1    g0864(.A(G322), .ZN(new_n1065));
  INV_X1    g0865(.A(G311), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n793), .A2(new_n1065), .B1(new_n773), .B2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n801), .A2(G303), .B1(KEYINPUT110), .B2(new_n1067), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(KEYINPUT110), .B2(new_n1067), .C1(new_n1029), .C2(new_n804), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT48), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1064), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n1070), .B2(new_n1069), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT49), .Z(new_n1073));
  AOI21_X1  g0873(.A(new_n253), .B1(new_n788), .B2(G326), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n614), .B2(new_n777), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1061), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1052), .B1(new_n1076), .B2(new_n768), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n977), .B2(new_n999), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1042), .A2(new_n1078), .ZN(G393));
  NAND3_X1  g0879(.A1(new_n990), .A2(new_n977), .A3(new_n991), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n958), .A2(new_n767), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n1066), .A2(new_n803), .B1(new_n793), .B2(new_n1029), .ZN(new_n1082));
  XOR2_X1   g0882(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n1083));
  XNOR2_X1  g0883(.A(new_n1082), .B(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n257), .B1(new_n784), .B2(new_n808), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1085), .B(new_n778), .C1(G116), .C2(new_n782), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n789), .A2(new_n1065), .B1(new_n1062), .B2(new_n796), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G303), .B2(new_n774), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1084), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n801), .A2(new_n400), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n253), .B1(new_n243), .B2(new_n784), .C1(new_n781), .C2(new_n341), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G87), .B2(new_n843), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n774), .A2(G50), .B1(G143), .B2(new_n788), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1090), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n1010), .A2(new_n793), .B1(new_n803), .B2(new_n790), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT51), .Z(new_n1096));
  OAI21_X1  g0896(.A(new_n1089), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n768), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n758), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n769), .B1(new_n1026), .B2(new_n210), .C1(new_n1099), .C2(new_n241), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1081), .A2(new_n753), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1041), .A2(new_n992), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n708), .B1(new_n1041), .B2(new_n992), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1080), .B(new_n1101), .C1(new_n1103), .C2(new_n1104), .ZN(G390));
  NAND3_X1  g0905(.A1(new_n896), .A2(new_n913), .A3(KEYINPUT39), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1106), .A2(new_n925), .A3(new_n924), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n914), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n765), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n849), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n753), .B1(new_n435), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n784), .A2(new_n1053), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT53), .Z(new_n1113));
  AOI211_X1 g0913(.A(new_n257), .B(new_n1113), .C1(G159), .C2(new_n782), .ZN(new_n1114));
  INV_X1    g0914(.A(G128), .ZN(new_n1115));
  INV_X1    g0915(.A(G132), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1114), .B1(new_n1115), .B2(new_n793), .C1(new_n1116), .C2(new_n803), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n774), .A2(G137), .B1(G125), .B2(new_n788), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT54), .B(G143), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n1118), .B1(new_n202), .B2(new_n777), .C1(new_n800), .C2(new_n1119), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n789), .A2(new_n1062), .B1(new_n387), .B2(new_n773), .ZN(new_n1121));
  NOR4_X1   g0921(.A1(new_n1121), .A2(new_n253), .A3(new_n785), .A4(new_n836), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1122), .B1(new_n808), .B2(new_n793), .C1(new_n1026), .C2(new_n800), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n803), .A2(new_n614), .B1(new_n341), .B2(new_n781), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT113), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n1117), .A2(new_n1120), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1111), .B1(new_n1126), .B2(new_n768), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1109), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n906), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n658), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n611), .A2(new_n661), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n673), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n679), .A2(new_n676), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n677), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n863), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n853), .ZN(new_n1138));
  OAI21_X1  g0938(.A(KEYINPUT99), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n865), .A2(new_n907), .A3(new_n853), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1129), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1108), .B1(new_n1141), .B2(new_n912), .ZN(new_n1142));
  OR2_X1    g0942(.A1(new_n855), .A2(new_n645), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n690), .B(new_n1143), .C1(new_n744), .C2(new_n745), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n853), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n906), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n895), .B1(new_n923), .B2(KEYINPUT38), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1146), .A2(new_n911), .A3(new_n1147), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n857), .B(G330), .C1(new_n731), .C2(new_n733), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1149), .A2(new_n1129), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1142), .A2(new_n1148), .A3(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n912), .B(new_n944), .C1(new_n1145), .C2(new_n906), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n911), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1153), .B1(new_n1155), .B2(new_n1108), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n936), .A2(G330), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n935), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1152), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1128), .B1(new_n1159), .B2(new_n978), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1157), .A2(new_n464), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n656), .B(new_n1162), .C1(new_n979), .C2(new_n931), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT112), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1154), .A2(new_n911), .B1(new_n1107), .B2(new_n914), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n935), .B(new_n1157), .C1(new_n1168), .C2(new_n1153), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n906), .B1(new_n1157), .B2(new_n860), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1170), .A2(new_n1145), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n1151), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1149), .A2(new_n1129), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n1158), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n908), .B2(new_n909), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1167), .A2(new_n1152), .A3(new_n1169), .A4(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n933), .A2(KEYINPUT112), .A3(new_n1162), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1178), .A2(new_n1179), .A3(new_n1176), .ZN(new_n1180));
  NOR3_X1   g0980(.A1(new_n1168), .A2(new_n1153), .A3(new_n1150), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1158), .B1(new_n1142), .B2(new_n1148), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1180), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1177), .A2(new_n1183), .A3(new_n708), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1161), .A2(new_n1184), .ZN(G378));
  AND2_X1   g0985(.A1(new_n927), .A2(new_n929), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n897), .A2(new_n1187), .A3(new_n898), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n938), .B1(new_n937), .B2(new_n1147), .ZN(new_n1189));
  OAI21_X1  g0989(.A(G330), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  XOR2_X1   g0990(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n461), .A2(new_n689), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n463), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT116), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n456), .A2(new_n459), .A3(new_n462), .A4(new_n1193), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1196), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1192), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(KEYINPUT116), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1203), .A2(new_n1191), .A3(new_n1198), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1201), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1190), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n947), .A2(new_n1205), .A3(G330), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1186), .A2(new_n1207), .A3(new_n910), .A4(new_n1208), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n947), .A2(G330), .A3(new_n1205), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1205), .B1(new_n947), .B2(G330), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n930), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1209), .A2(new_n1212), .A3(new_n977), .ZN(new_n1213));
  INV_X1    g1013(.A(G137), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n796), .A2(new_n1214), .B1(new_n773), .B2(new_n1116), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT115), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1119), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n782), .A2(G150), .B1(new_n815), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(G125), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1218), .B1(new_n1219), .B2(new_n793), .C1(new_n1115), .C2(new_n803), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1216), .A2(new_n1220), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1223));
  INV_X1    g1023(.A(G41), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n617), .B(new_n1224), .C1(new_n777), .C2(new_n790), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G124), .B2(new_n788), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1222), .A2(new_n1223), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n843), .A2(G58), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n257), .A2(new_n1224), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n815), .B2(G77), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1228), .B(new_n1230), .C1(new_n789), .C2(new_n808), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT114), .Z(new_n1232));
  OAI221_X1 g1032(.A(new_n1012), .B1(new_n773), .B2(new_n1026), .C1(new_n403), .C2(new_n796), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n387), .A2(new_n803), .B1(new_n793), .B2(new_n614), .ZN(new_n1234));
  OR3_X1    g1034(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT58), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1229), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1239));
  AND4_X1   g1039(.A1(new_n1227), .A2(new_n1237), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n753), .B1(G50), .B2(new_n1110), .C1(new_n1240), .C2(new_n821), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1205), .B2(new_n765), .ZN(new_n1242));
  XOR2_X1   g1042(.A(new_n1242), .B(KEYINPUT117), .Z(new_n1243));
  NAND2_X1  g1043(.A1(new_n1213), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(KEYINPUT118), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT118), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1213), .A2(new_n1246), .A3(new_n1243), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1249), .B1(new_n1250), .B2(new_n1176), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1209), .A2(new_n1212), .A3(KEYINPUT57), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n708), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1167), .B1(new_n1159), .B2(new_n1180), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1209), .A2(new_n1212), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT57), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1248), .B1(new_n1253), .B2(new_n1256), .ZN(G375));
  NOR2_X1   g1057(.A1(new_n906), .A2(new_n766), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT119), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n843), .A2(G77), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n774), .A2(G116), .B1(G303), .B2(new_n788), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n253), .B1(new_n815), .B2(G97), .ZN(new_n1262));
  AND4_X1   g1062(.A1(new_n1260), .A2(new_n1261), .A3(new_n1056), .A4(new_n1262), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(G283), .A2(new_n818), .B1(new_n811), .B2(G294), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1263), .B(new_n1264), .C1(new_n387), .C2(new_n800), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(KEYINPUT120), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n797), .A2(G150), .B1(G50), .B2(new_n782), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT122), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n257), .B1(new_n815), .B2(G159), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1228), .B(new_n1271), .C1(new_n789), .C2(new_n1115), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n811), .A2(G132), .B1(new_n774), .B2(new_n1217), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(new_n804), .B2(new_n1214), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1269), .B(new_n1273), .C1(new_n1275), .C2(KEYINPUT121), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(KEYINPUT121), .B2(new_n1275), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n768), .B1(new_n1266), .B2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1278), .B(new_n753), .C1(G68), .C2(new_n1110), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1259), .A2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n1176), .B2(new_n977), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1001), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1180), .A2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1176), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1281), .B1(new_n1283), .B2(new_n1284), .ZN(G381));
  NAND2_X1  g1085(.A1(new_n1080), .A2(new_n1101), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1104), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1286), .B1(new_n1287), .B2(new_n1102), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1042), .A2(new_n826), .A3(new_n1078), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1288), .A2(new_n1290), .A3(new_n870), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(G387), .A2(G381), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(G375), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n709), .B1(new_n1159), .B2(new_n1180), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1160), .B1(new_n1177), .B2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1292), .A2(new_n1293), .A3(new_n1295), .ZN(G407));
  INV_X1    g1096(.A(G213), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1297), .A2(G343), .ZN(new_n1298));
  XOR2_X1   g1098(.A(new_n1298), .B(KEYINPUT123), .Z(new_n1299));
  NAND3_X1  g1099(.A1(new_n1293), .A2(new_n1295), .A3(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(G407), .A2(new_n1300), .A3(G213), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(KEYINPUT124), .ZN(G409));
  AOI21_X1  g1102(.A(new_n826), .B1(new_n1042), .B2(new_n1078), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1288), .B1(new_n1290), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(G393), .A2(G396), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1305), .A2(G390), .A3(new_n1289), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(G387), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1304), .A2(new_n1003), .A3(new_n1306), .A4(new_n1037), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1308), .A2(KEYINPUT126), .A3(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT126), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  OAI211_X1 g1113(.A(G378), .B(new_n1248), .C1(new_n1253), .C2(new_n1256), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1254), .A2(new_n1282), .A3(new_n1255), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1295), .B1(new_n1315), .B2(new_n1244), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1298), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1284), .B1(KEYINPUT60), .B2(new_n1180), .ZN(new_n1319));
  AND2_X1   g1119(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1320), .B(KEYINPUT60), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n708), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1281), .B1(new_n1319), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n870), .ZN(new_n1324));
  OAI211_X1 g1124(.A(G384), .B(new_n1281), .C1(new_n1319), .C2(new_n1322), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1317), .A2(new_n1318), .A3(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT62), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1299), .B1(new_n1314), .B2(new_n1316), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1326), .A2(new_n1329), .ZN(new_n1331));
  AOI22_X1  g1131(.A1(new_n1328), .A2(new_n1329), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT61), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1299), .A2(G2897), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1326), .A2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1298), .A2(G2897), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1324), .A2(new_n1325), .A3(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1336), .A2(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1333), .B1(new_n1339), .B2(new_n1330), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1313), .B1(new_n1332), .B2(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1298), .B1(new_n1314), .B2(new_n1316), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT125), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1343), .A2(new_n1344), .A3(new_n1338), .A4(new_n1336), .ZN(new_n1345));
  OAI21_X1  g1145(.A(KEYINPUT125), .B1(new_n1339), .B2(new_n1342), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT63), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1328), .A2(new_n1347), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1308), .A2(new_n1333), .A3(new_n1309), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1326), .A2(new_n1347), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1349), .B1(new_n1330), .B2(new_n1350), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1345), .A2(new_n1346), .A3(new_n1348), .A4(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1341), .A2(new_n1352), .ZN(G405));
  NAND2_X1  g1153(.A1(G375), .A2(new_n1295), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1354), .A2(new_n1314), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT127), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1355), .A2(new_n1356), .A3(new_n1326), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1326), .A2(new_n1356), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1324), .A2(KEYINPUT127), .A3(new_n1325), .ZN(new_n1359));
  NAND4_X1  g1159(.A1(new_n1358), .A2(new_n1354), .A3(new_n1314), .A4(new_n1359), .ZN(new_n1360));
  AND3_X1   g1160(.A1(new_n1312), .A2(new_n1357), .A3(new_n1360), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1312), .B1(new_n1357), .B2(new_n1360), .ZN(new_n1362));
  NOR2_X1   g1162(.A1(new_n1361), .A2(new_n1362), .ZN(G402));
endmodule


