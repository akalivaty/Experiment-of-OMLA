//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT73), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G140), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT74), .B1(new_n191), .B2(G125), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT74), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(new_n189), .A3(G140), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(KEYINPUT73), .A3(G125), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n190), .A2(new_n192), .A3(new_n194), .A4(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT16), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT16), .B1(new_n191), .B2(G125), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n187), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  AOI211_X1 g014(.A(G146), .B(new_n198), .C1(new_n196), .C2(KEYINPUT16), .ZN(new_n201));
  OR2_X1    g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G119), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT71), .B1(new_n203), .B2(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT23), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G119), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(KEYINPUT71), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n203), .A2(G128), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n205), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G110), .ZN(new_n212));
  XNOR2_X1  g026(.A(new_n212), .B(KEYINPUT72), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n207), .A2(new_n210), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT24), .B(G110), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n202), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  OR3_X1    g030(.A1(new_n211), .A2(KEYINPUT75), .A3(G110), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT75), .B1(new_n211), .B2(G110), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n214), .A2(new_n215), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n200), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n191), .A2(G125), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n189), .A2(G140), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n223), .A3(new_n187), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n220), .A2(new_n221), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n216), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT22), .B(G137), .ZN(new_n227));
  INV_X1    g041(.A(G953), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n228), .A2(G221), .A3(G234), .ZN(new_n229));
  XOR2_X1   g043(.A(new_n227), .B(new_n229), .Z(new_n230));
  NAND2_X1  g044(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n230), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n216), .A2(new_n225), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G217), .ZN(new_n235));
  INV_X1    g049(.A(G902), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n235), .B1(G234), .B2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(G902), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n237), .ZN(new_n240));
  AOI21_X1  g054(.A(G902), .B1(new_n231), .B2(new_n233), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT25), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n241), .A2(new_n242), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n239), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n187), .A2(G143), .ZN(new_n247));
  INV_X1    g061(.A(G143), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G146), .ZN(new_n249));
  AND2_X1   g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n247), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT65), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(G143), .B(G146), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(KEYINPUT65), .A3(new_n250), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT0), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(new_n206), .A3(KEYINPUT64), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT64), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n258), .B1(KEYINPUT0), .B2(G128), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n250), .B1(new_n247), .B2(new_n249), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n253), .A2(new_n255), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n263));
  INV_X1    g077(.A(G137), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(G134), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT11), .ZN(new_n266));
  INV_X1    g080(.A(G134), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n266), .B1(new_n267), .B2(G137), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(KEYINPUT67), .A3(G137), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n264), .A2(KEYINPUT11), .A3(G134), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n265), .A2(new_n268), .A3(new_n269), .A4(new_n270), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n271), .A2(G131), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(G131), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n262), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n247), .A2(new_n249), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n247), .A2(KEYINPUT1), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n276), .A3(G128), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n247), .B(new_n249), .C1(KEYINPUT1), .C2(new_n206), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OR2_X1    g093(.A1(new_n271), .A2(G131), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT68), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n281), .B1(G134), .B2(new_n264), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n267), .A2(KEYINPUT68), .A3(G137), .ZN(new_n283));
  OAI22_X1  g097(.A1(new_n282), .A2(new_n283), .B1(G134), .B2(new_n264), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G131), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n279), .A2(new_n280), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n203), .A2(G116), .ZN(new_n287));
  INV_X1    g101(.A(G116), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G119), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT2), .B(G113), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n290), .B(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n274), .A2(new_n286), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(G237), .A2(G953), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G210), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n296), .B(KEYINPUT27), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT26), .B(G101), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n297), .B(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT69), .B1(new_n294), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n274), .A2(new_n286), .A3(new_n293), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT69), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n303), .A3(new_n299), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G131), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n271), .B(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n261), .A2(new_n260), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT65), .B1(new_n254), .B2(new_n250), .ZN(new_n310));
  AND4_X1   g124(.A1(KEYINPUT65), .A2(new_n247), .A3(new_n249), .A4(new_n250), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n312), .A2(KEYINPUT66), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT66), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n253), .A2(new_n255), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(new_n309), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n308), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT30), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(new_n286), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n274), .A2(new_n286), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT30), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n293), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT31), .B1(new_n305), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n262), .A2(new_n314), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n312), .A2(KEYINPUT66), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n307), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n286), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n326), .A2(KEYINPUT30), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n321), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n292), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n302), .A2(new_n303), .A3(new_n299), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n303), .B1(new_n302), .B2(new_n299), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT31), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n330), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT28), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n292), .B1(new_n326), .B2(new_n327), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n336), .B1(new_n337), .B2(new_n302), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n294), .A2(KEYINPUT28), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n300), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n323), .A2(new_n335), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G472), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n342), .A3(new_n236), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT32), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT32), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n341), .A2(new_n345), .A3(new_n342), .A4(new_n236), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n300), .B1(new_n322), .B2(new_n294), .ZN(new_n348));
  INV_X1    g162(.A(new_n339), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n317), .A2(new_n286), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n294), .B1(new_n350), .B2(new_n292), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n299), .B(new_n349), .C1(new_n351), .C2(new_n336), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n348), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT70), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT70), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n348), .A2(new_n352), .A3(new_n356), .A4(new_n353), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n320), .A2(new_n292), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n336), .B1(new_n358), .B2(new_n302), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(new_n339), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n300), .A2(new_n353), .ZN(new_n361));
  AOI21_X1  g175(.A(G902), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n355), .A2(new_n357), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G472), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n246), .B1(new_n347), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT78), .ZN(new_n366));
  INV_X1    g180(.A(G107), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(G104), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT3), .ZN(new_n369));
  INV_X1    g183(.A(G104), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n369), .B1(new_n370), .B2(G107), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n367), .A2(KEYINPUT3), .A3(G104), .ZN(new_n372));
  AOI211_X1 g186(.A(G101), .B(new_n368), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G101), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n367), .B2(G104), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n370), .A2(KEYINPUT77), .A3(G107), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n367), .A2(G104), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n374), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n366), .B1(new_n373), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n370), .A2(G107), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n367), .A2(KEYINPUT3), .A3(G104), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT3), .B1(new_n367), .B2(G104), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n374), .B(new_n382), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n376), .A2(new_n377), .B1(G104), .B2(new_n367), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n385), .B(KEYINPUT78), .C1(new_n374), .C2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n381), .A2(new_n279), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT10), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n385), .B1(new_n374), .B2(new_n386), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n277), .A2(new_n278), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT10), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G101), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n396), .A2(KEYINPUT76), .A3(KEYINPUT4), .A4(new_n385), .ZN(new_n397));
  NAND2_X1  g211(.A1(KEYINPUT76), .A2(KEYINPUT4), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n395), .A2(G101), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n397), .A2(new_n262), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n394), .A2(new_n307), .A3(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G110), .B(G140), .ZN(new_n402));
  INV_X1    g216(.A(G227), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(G953), .ZN(new_n404));
  XOR2_X1   g218(.A(new_n402), .B(new_n404), .Z(new_n405));
  INV_X1    g219(.A(KEYINPUT12), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT79), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n406), .B1(new_n307), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n387), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n370), .A2(KEYINPUT77), .A3(G107), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT77), .B1(new_n370), .B2(G107), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n379), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G101), .ZN(new_n413));
  AOI21_X1  g227(.A(KEYINPUT78), .B1(new_n413), .B2(new_n385), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n391), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n390), .A2(new_n391), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n408), .B1(new_n418), .B2(new_n308), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n279), .B1(new_n381), .B2(new_n387), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n308), .B(new_n408), .C1(new_n420), .C2(new_n416), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n401), .B(new_n405), .C1(new_n419), .C2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n392), .B1(new_n388), .B2(KEYINPUT10), .ZN(new_n424));
  INV_X1    g238(.A(new_n400), .ZN(new_n425));
  NOR3_X1   g239(.A1(new_n424), .A2(new_n308), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n308), .B1(new_n424), .B2(new_n425), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT80), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT80), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n429), .B(new_n308), .C1(new_n424), .C2(new_n425), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n426), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n423), .B1(new_n431), .B2(new_n405), .ZN(new_n432));
  XOR2_X1   g246(.A(KEYINPUT81), .B(G469), .Z(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n236), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n428), .A2(new_n430), .ZN(new_n435));
  INV_X1    g249(.A(new_n405), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n426), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n401), .B1(new_n419), .B2(new_n422), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n435), .A2(new_n437), .B1(new_n438), .B2(new_n436), .ZN(new_n439));
  OAI21_X1  g253(.A(G469), .B1(new_n439), .B2(G902), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n434), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT9), .B(G234), .ZN(new_n442));
  OAI21_X1  g256(.A(G221), .B1(new_n442), .B2(G902), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT82), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n443), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n434), .B2(new_n440), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT82), .ZN(new_n449));
  INV_X1    g263(.A(G237), .ZN(new_n450));
  AND4_X1   g264(.A1(G143), .A2(new_n450), .A3(new_n228), .A4(G214), .ZN(new_n451));
  AOI21_X1  g265(.A(G143), .B1(new_n295), .B2(G214), .ZN(new_n452));
  OAI21_X1  g266(.A(G131), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT18), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n224), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n456), .B1(new_n196), .B2(G146), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n450), .A2(new_n228), .A3(G214), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n248), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n295), .A2(G143), .A3(G214), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n454), .A2(new_n306), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OR3_X1    g277(.A1(new_n455), .A2(new_n457), .A3(new_n463), .ZN(new_n464));
  XOR2_X1   g278(.A(G113), .B(G122), .Z(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT88), .B(G104), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT17), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT89), .B1(new_n453), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT89), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n461), .A2(new_n470), .A3(KEYINPUT17), .A4(G131), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n459), .A2(new_n306), .A3(new_n460), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n453), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n469), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n464), .B(new_n467), .C1(new_n202), .C2(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n475), .A2(KEYINPUT90), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT90), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n455), .A2(new_n457), .A3(new_n463), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n469), .A2(new_n471), .A3(new_n473), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n200), .A2(new_n201), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n477), .B1(new_n481), .B2(new_n467), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n453), .A2(new_n472), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n196), .A2(KEYINPUT19), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n196), .A2(KEYINPUT87), .A3(KEYINPUT19), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT19), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n222), .A2(new_n223), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n221), .B(new_n483), .C1(new_n490), .C2(G146), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n491), .A2(new_n464), .ZN(new_n492));
  OAI22_X1  g306(.A1(new_n476), .A2(new_n482), .B1(new_n492), .B2(new_n467), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT20), .ZN(new_n494));
  NOR2_X1   g308(.A1(G475), .A2(G902), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  XOR2_X1   g310(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n467), .B1(new_n491), .B2(new_n464), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n475), .A2(KEYINPUT90), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n481), .A2(new_n477), .A3(new_n467), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n495), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n498), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OR2_X1    g318(.A1(new_n481), .A2(new_n467), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(new_n476), .B2(new_n482), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n236), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n496), .A2(new_n504), .B1(new_n507), .B2(G475), .ZN(new_n508));
  NAND2_X1  g322(.A1(G234), .A2(G237), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n509), .A2(G952), .A3(new_n228), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(G902), .A3(G953), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(KEYINPUT94), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT21), .B(G898), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n288), .A2(G122), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT14), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  AND2_X1   g331(.A1(KEYINPUT91), .A2(G122), .ZN(new_n518));
  NOR2_X1   g332(.A1(KEYINPUT91), .A2(G122), .ZN(new_n519));
  OAI21_X1  g333(.A(G116), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n367), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n248), .A2(G128), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n206), .A2(G143), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(new_n267), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n520), .A2(new_n367), .A3(new_n515), .ZN(new_n526));
  OR3_X1    g340(.A1(new_n521), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n442), .A2(new_n235), .A3(G953), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT92), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT13), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n267), .B1(new_n523), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n531), .A2(new_n524), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n524), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n367), .B1(new_n520), .B2(new_n515), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n532), .B(new_n533), .C1(new_n526), .C2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n527), .A2(new_n529), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n529), .B1(new_n527), .B2(new_n535), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n236), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT93), .ZN(new_n540));
  INV_X1    g354(.A(new_n538), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n536), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT93), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n543), .A3(new_n236), .ZN(new_n544));
  INV_X1    g358(.A(G478), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(KEYINPUT15), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n540), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n542), .A2(new_n543), .A3(new_n236), .A4(new_n546), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n514), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n508), .A2(new_n550), .ZN(new_n551));
  OR2_X1    g365(.A1(new_n290), .A2(new_n291), .ZN(new_n552));
  INV_X1    g366(.A(new_n290), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT5), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n287), .A2(KEYINPUT5), .ZN(new_n555));
  INV_X1    g369(.A(G113), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n381), .A2(new_n552), .A3(new_n387), .A4(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n397), .A2(new_n292), .A3(new_n399), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(G110), .B(G122), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(KEYINPUT6), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT6), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n561), .A2(new_n567), .A3(new_n563), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n309), .B(G125), .C1(new_n310), .C2(new_n311), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n277), .A2(new_n189), .A3(new_n278), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n228), .A2(G224), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n571), .B(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n566), .A2(new_n568), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(KEYINPUT7), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n569), .A2(new_n570), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n575), .B1(new_n569), .B2(new_n570), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n565), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n558), .A2(new_n552), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n390), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT84), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n557), .B1(new_n554), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(KEYINPUT84), .B1(new_n553), .B2(KEYINPUT5), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n552), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n381), .A2(new_n387), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n581), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n562), .B(KEYINPUT8), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(G902), .B1(new_n579), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n574), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(G210), .B1(G237), .B2(G902), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n574), .A2(new_n590), .A3(new_n592), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(KEYINPUT85), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT85), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n574), .A2(new_n590), .A3(new_n597), .A4(new_n592), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(G214), .B1(G237), .B2(G902), .ZN(new_n600));
  XOR2_X1   g414(.A(new_n600), .B(KEYINPUT83), .Z(new_n601));
  NOR3_X1   g415(.A1(new_n551), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n365), .A2(new_n446), .A3(new_n449), .A4(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  NAND2_X1  g418(.A1(new_n341), .A2(new_n236), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(G472), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT95), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n607), .A3(new_n343), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n605), .A2(KEYINPUT95), .A3(G472), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n246), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(new_n446), .A3(new_n449), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT96), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n496), .A2(new_n504), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n507), .A2(G475), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n542), .A2(new_n545), .A3(new_n236), .ZN(new_n617));
  OAI21_X1  g431(.A(KEYINPUT33), .B1(new_n537), .B2(new_n538), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n541), .A2(new_n619), .A3(new_n536), .ZN(new_n620));
  AOI21_X1  g434(.A(G902), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n617), .B1(new_n621), .B2(new_n545), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n616), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n601), .B1(new_n594), .B2(new_n595), .ZN(new_n625));
  INV_X1    g439(.A(new_n514), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n613), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n622), .B1(new_n614), .B2(new_n615), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n629), .A2(KEYINPUT96), .A3(new_n626), .A4(new_n625), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n612), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n632), .B(KEYINPUT97), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT34), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G104), .ZN(G6));
  AND2_X1   g449(.A1(new_n548), .A2(new_n549), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n493), .A2(new_n495), .A3(new_n497), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n504), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n638), .A2(new_n615), .ZN(new_n639));
  AND4_X1   g453(.A1(new_n636), .A2(new_n639), .A3(new_n626), .A4(new_n625), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n612), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT98), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT35), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G107), .ZN(G9));
  NAND3_X1  g458(.A1(new_n446), .A2(new_n449), .A3(new_n602), .ZN(new_n645));
  INV_X1    g459(.A(new_n245), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n232), .A2(KEYINPUT36), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n226), .B(new_n647), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n646), .A2(new_n243), .B1(new_n238), .B2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n343), .A2(new_n607), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n342), .B1(new_n341), .B2(new_n236), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n609), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(KEYINPUT99), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n608), .A2(new_n609), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT99), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n657), .A2(new_n658), .A3(new_n650), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n645), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT37), .B(G110), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  NAND2_X1  g476(.A1(new_n347), .A2(new_n364), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n650), .ZN(new_n664));
  INV_X1    g478(.A(new_n510), .ZN(new_n665));
  INV_X1    g479(.A(G900), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n512), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n665), .B1(new_n667), .B2(KEYINPUT100), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(KEYINPUT100), .B2(new_n667), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n636), .A2(new_n638), .A3(new_n615), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT101), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n664), .A2(new_n672), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n446), .A2(new_n449), .A3(new_n625), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G128), .ZN(G30));
  NAND2_X1  g490(.A1(new_n446), .A2(new_n449), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n669), .B(KEYINPUT39), .Z(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n305), .A2(new_n322), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n299), .B1(new_n358), .B2(new_n302), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n236), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G472), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n347), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n599), .B(KEYINPUT38), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n616), .A2(new_n636), .ZN(new_n690));
  INV_X1    g504(.A(new_n601), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n649), .A2(new_n691), .ZN(new_n692));
  NOR4_X1   g506(.A1(new_n688), .A2(new_n689), .A3(new_n690), .A4(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n681), .A2(new_n682), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G143), .ZN(G45));
  AOI22_X1  g509(.A1(new_n344), .A2(new_n346), .B1(new_n363), .B2(G472), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n629), .A2(new_n670), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n696), .A2(new_n649), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n674), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G146), .ZN(G48));
  INV_X1    g514(.A(new_n434), .ZN(new_n701));
  INV_X1    g515(.A(G469), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n432), .B2(new_n236), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n701), .A2(new_n703), .A3(new_n447), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n631), .A2(new_n365), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT41), .B(G113), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G15));
  NAND3_X1  g521(.A1(new_n365), .A2(new_n704), .A3(new_n640), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G116), .ZN(G18));
  NAND2_X1  g523(.A1(new_n704), .A2(new_n625), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n696), .A2(new_n649), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT102), .ZN(new_n713));
  INV_X1    g527(.A(new_n551), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n711), .A2(new_n712), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n663), .A2(new_n714), .A3(new_n650), .ZN(new_n716));
  OAI21_X1  g530(.A(KEYINPUT102), .B1(new_n716), .B2(new_n710), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  INV_X1    g533(.A(KEYINPUT103), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n300), .B1(new_n359), .B2(new_n339), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n323), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n335), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n720), .B1(new_n323), .B2(new_n721), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n342), .B(new_n236), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n606), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n246), .ZN(new_n727));
  INV_X1    g541(.A(new_n625), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n690), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n727), .A2(new_n626), .A3(new_n704), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  NOR2_X1   g545(.A1(new_n726), .A2(new_n649), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT104), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n629), .B2(new_n670), .ZN(new_n734));
  NOR4_X1   g548(.A1(new_n508), .A2(KEYINPUT104), .A3(new_n622), .A4(new_n669), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n711), .A2(new_n732), .A3(new_n736), .ZN(new_n737));
  XOR2_X1   g551(.A(KEYINPUT105), .B(G125), .Z(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G27));
  AOI21_X1  g553(.A(KEYINPUT106), .B1(new_n599), .B2(new_n691), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT106), .ZN(new_n741));
  AOI211_X1 g555(.A(new_n741), .B(new_n601), .C1(new_n596), .C2(new_n598), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(new_n736), .A3(new_n365), .A4(new_n448), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n740), .A2(new_n742), .A3(new_n444), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n747), .A2(KEYINPUT42), .A3(new_n365), .A4(new_n736), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G131), .ZN(G33));
  XOR2_X1   g564(.A(new_n671), .B(KEYINPUT101), .Z(new_n751));
  NAND3_X1  g565(.A1(new_n747), .A2(new_n751), .A3(new_n365), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT107), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  NOR2_X1   g569(.A1(new_n439), .A2(KEYINPUT45), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n702), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n757), .A2(KEYINPUT108), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(KEYINPUT108), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n439), .A2(KEYINPUT45), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(G469), .A2(G902), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(KEYINPUT46), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n434), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT46), .B1(new_n761), .B2(new_n762), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n443), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n767));
  INV_X1    g581(.A(new_n679), .ZN(new_n768));
  OR3_X1    g582(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n508), .A2(new_n623), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(KEYINPUT43), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n771), .A2(new_n657), .A3(new_n649), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT44), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n743), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n772), .A2(KEYINPUT44), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n775), .A2(KEYINPUT110), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(KEYINPUT110), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n767), .B1(new_n766), .B2(new_n768), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n769), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(KEYINPUT111), .B(G137), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G39));
  XOR2_X1   g596(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n783));
  NAND2_X1  g597(.A1(new_n766), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n783), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n443), .B(new_n785), .C1(new_n764), .C2(new_n765), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n740), .A2(new_n742), .ZN(new_n787));
  INV_X1    g601(.A(new_n246), .ZN(new_n788));
  NOR4_X1   g602(.A1(new_n787), .A2(new_n663), .A3(new_n788), .A4(new_n697), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n784), .A2(new_n786), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  NAND4_X1  g605(.A1(new_n596), .A2(new_n691), .A3(new_n598), .A4(new_n626), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n508), .A2(new_n636), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n610), .A2(new_n446), .A3(new_n449), .A4(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT115), .B1(new_n660), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n658), .B1(new_n657), .B2(new_n650), .ZN(new_n799));
  AOI211_X1 g613(.A(KEYINPUT99), .B(new_n649), .C1(new_n608), .C2(new_n609), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n798), .B(new_n795), .C1(new_n801), .C2(new_n645), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n803));
  OR3_X1    g617(.A1(new_n792), .A2(new_n624), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n803), .B1(new_n792), .B2(new_n624), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n603), .B1(new_n806), .B2(new_n611), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n797), .A2(new_n802), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT116), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n795), .B1(new_n801), .B2(new_n645), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n807), .B1(new_n811), .B2(KEYINPUT115), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n812), .A2(new_n813), .A3(new_n802), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n636), .A2(new_n669), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n639), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n787), .A2(new_n664), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(KEYINPUT117), .A3(new_n678), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n712), .A2(new_n743), .A3(new_n639), .A4(new_n816), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n820), .B1(new_n821), .B2(new_n677), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n726), .A2(new_n734), .A3(new_n735), .A4(new_n649), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n747), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n754), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n705), .A2(new_n730), .A3(new_n708), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n749), .A2(new_n718), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n650), .A2(new_n669), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n687), .A3(new_n448), .A4(new_n729), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n675), .A2(new_n699), .A3(new_n737), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n673), .A2(new_n674), .B1(new_n824), .B2(new_n711), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(KEYINPUT52), .A3(new_n699), .A4(new_n832), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n830), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  AND4_X1   g652(.A1(new_n815), .A2(new_n826), .A3(new_n829), .A4(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n754), .A2(new_n823), .A3(new_n825), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n810), .B2(new_n814), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n828), .B1(new_n835), .B2(new_n837), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT53), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT54), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n813), .B1(new_n812), .B2(new_n802), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n813), .A2(new_n797), .A3(new_n802), .A4(new_n808), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n826), .B(new_n842), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n830), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n827), .A2(new_n718), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n827), .A2(new_n718), .A3(KEYINPUT118), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n852), .A2(new_n853), .B1(new_n746), .B2(new_n748), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n815), .A2(new_n826), .A3(new_n838), .A4(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n848), .A2(new_n849), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n844), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n771), .A2(new_n665), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n858), .A2(new_n727), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n689), .A2(new_n601), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n859), .A2(new_n704), .A3(new_n860), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT50), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n688), .A2(new_n788), .A3(new_n510), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n743), .A2(new_n704), .ZN(new_n864));
  OR3_X1    g678(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT119), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT119), .B1(new_n863), .B2(new_n864), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n508), .A2(new_n865), .A3(new_n622), .A4(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n864), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n868), .A2(new_n732), .A3(new_n858), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n862), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n701), .A2(new_n703), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n784), .A2(new_n786), .B1(new_n447), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n859), .A2(new_n743), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n870), .B(KEYINPUT51), .C1(new_n872), .C2(new_n873), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n868), .A2(new_n365), .A3(new_n858), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT48), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n865), .A2(new_n629), .A3(new_n866), .ZN(new_n880));
  INV_X1    g694(.A(G952), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n881), .B(G953), .C1(new_n859), .C2(new_n711), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT120), .Z(new_n884));
  NAND3_X1  g698(.A1(new_n876), .A2(new_n877), .A3(new_n884), .ZN(new_n885));
  OAI22_X1  g699(.A1(new_n857), .A2(new_n885), .B1(G952), .B2(G953), .ZN(new_n886));
  NOR4_X1   g700(.A1(new_n246), .A2(new_n770), .A3(new_n447), .A4(new_n601), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT113), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n871), .B(KEYINPUT49), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n888), .A2(new_n689), .A3(new_n688), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n886), .A2(new_n890), .ZN(G75));
  NOR2_X1   g705(.A1(new_n228), .A2(G952), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT122), .Z(new_n893));
  AOI21_X1  g707(.A(new_n236), .B1(new_n848), .B2(new_n855), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n894), .A2(G210), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n566), .A2(new_n568), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(new_n573), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT55), .ZN(new_n898));
  XOR2_X1   g712(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n893), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n894), .A2(G210), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT56), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n898), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n901), .A2(new_n904), .ZN(G51));
  XOR2_X1   g719(.A(new_n762), .B(KEYINPUT57), .Z(new_n906));
  AND3_X1   g720(.A1(new_n848), .A2(new_n849), .A3(new_n855), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n849), .B1(new_n848), .B2(new_n855), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n432), .ZN(new_n910));
  INV_X1    g724(.A(new_n761), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n894), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n892), .B1(new_n910), .B2(new_n912), .ZN(G54));
  AND2_X1   g727(.A1(KEYINPUT58), .A2(G475), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n894), .A2(new_n493), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n493), .B1(new_n894), .B2(new_n914), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n915), .A2(new_n916), .A3(new_n892), .ZN(G60));
  NAND2_X1  g731(.A1(G478), .A2(G902), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT59), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n618), .A2(new_n620), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT123), .Z(new_n921));
  OAI211_X1 g735(.A(new_n919), .B(new_n921), .C1(new_n907), .C2(new_n908), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n893), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n921), .B1(new_n857), .B2(new_n919), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(G63));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n848), .A2(new_n855), .ZN(new_n927));
  NAND2_X1  g741(.A1(G217), .A2(G902), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT124), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT60), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n648), .B(KEYINPUT125), .Z(new_n931));
  NAND3_X1  g745(.A1(new_n927), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n893), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n234), .B1(new_n927), .B2(new_n930), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n926), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n927), .A2(new_n930), .ZN(new_n936));
  INV_X1    g750(.A(new_n234), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n938), .A2(KEYINPUT61), .A3(new_n893), .A4(new_n932), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n935), .A2(new_n939), .ZN(G66));
  AOI21_X1  g754(.A(new_n850), .B1(new_n810), .B2(new_n814), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n941), .A2(G953), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n942), .A2(KEYINPUT126), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(KEYINPUT126), .ZN(new_n944));
  INV_X1    g758(.A(G224), .ZN(new_n945));
  OAI21_X1  g759(.A(G953), .B1(new_n513), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n896), .B1(G898), .B2(new_n228), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(G69));
  AND2_X1   g763(.A1(new_n836), .A2(new_n699), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n790), .A2(new_n749), .A3(new_n754), .A4(new_n950), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n769), .A2(new_n779), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n365), .A2(new_n729), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n778), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n951), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n228), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n328), .A2(new_n329), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(new_n490), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(new_n666), .B2(new_n228), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n694), .A2(new_n950), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT62), .Z(new_n963));
  NOR2_X1   g777(.A1(new_n677), .A2(new_n768), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n624), .A2(new_n793), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n964), .A2(new_n365), .A3(new_n743), .A4(new_n965), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n780), .A2(new_n790), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(G953), .B1(new_n963), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n961), .B1(new_n968), .B2(new_n958), .ZN(new_n969));
  INV_X1    g783(.A(new_n958), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n970), .A2(KEYINPUT127), .ZN(new_n971));
  OAI21_X1  g785(.A(G953), .B1(new_n403), .B2(new_n666), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  OAI221_X1 g788(.A(new_n961), .B1(new_n971), .B2(new_n972), .C1(new_n968), .C2(new_n958), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(G72));
  OAI21_X1  g790(.A(new_n299), .B1(new_n322), .B2(new_n294), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n963), .A2(new_n967), .A3(new_n941), .ZN(new_n978));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT63), .Z(new_n980));
  AOI21_X1  g794(.A(new_n977), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n330), .A2(new_n300), .A3(new_n302), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n955), .A2(new_n941), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n982), .B1(new_n983), .B2(new_n980), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n839), .A2(new_n843), .ZN(new_n985));
  INV_X1    g799(.A(new_n348), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n980), .B1(new_n986), .B2(new_n683), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NOR4_X1   g802(.A1(new_n981), .A2(new_n984), .A3(new_n988), .A4(new_n892), .ZN(G57));
endmodule


