//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT72), .A2(G953), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT72), .A2(G953), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G227), .ZN(new_n192));
  XOR2_X1   g006(.A(G110), .B(G140), .Z(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT86), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n197));
  XNOR2_X1  g011(.A(G143), .B(G146), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G128), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT68), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT68), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n200), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT64), .B1(new_n209), .B2(G146), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(new_n206), .A3(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(G146), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n199), .B1(new_n208), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT71), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n207), .ZN(new_n218));
  OAI21_X1  g032(.A(G128), .B1(new_n197), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(KEYINPUT71), .A3(new_n199), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT82), .ZN(new_n223));
  XNOR2_X1  g037(.A(G104), .B(G107), .ZN(new_n224));
  INV_X1    g038(.A(G101), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G104), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT3), .B1(new_n227), .B2(G107), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n229));
  INV_X1    g043(.A(G107), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(G104), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n227), .A2(G107), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n228), .A2(new_n231), .A3(new_n225), .A4(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n227), .A2(G107), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n230), .A2(G104), .ZN(new_n235));
  OAI211_X1 g049(.A(KEYINPUT82), .B(G101), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n226), .A2(new_n233), .A3(new_n236), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n217), .A2(KEYINPUT10), .A3(new_n222), .A4(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n228), .A2(new_n231), .A3(new_n232), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G101), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(KEYINPUT4), .A3(new_n233), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT81), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n241), .B(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n220), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT65), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n220), .A2(KEYINPUT65), .A3(new_n246), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n249), .A2(new_n250), .B1(new_n198), .B2(new_n244), .ZN(new_n251));
  OR2_X1    g065(.A1(new_n240), .A2(KEYINPUT4), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n238), .B1(new_n243), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(G128), .B1(new_n207), .B2(new_n213), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n209), .A2(KEYINPUT1), .A3(G146), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT83), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT83), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n259), .B(new_n256), .C1(new_n198), .C2(G128), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n258), .A2(new_n199), .A3(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n226), .A2(new_n233), .A3(new_n236), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT84), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n258), .A2(new_n199), .A3(new_n260), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT84), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(new_n237), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT10), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n196), .B1(new_n254), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT11), .ZN(new_n269));
  INV_X1    g083(.A(G134), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n269), .B1(new_n270), .B2(G137), .ZN(new_n271));
  INV_X1    g085(.A(G137), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(KEYINPUT11), .A3(G134), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n270), .A2(G137), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n271), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G131), .ZN(new_n276));
  INV_X1    g090(.A(G131), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n271), .A2(new_n273), .A3(new_n277), .A4(new_n274), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT10), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n264), .A2(new_n237), .A3(new_n265), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n265), .B1(new_n264), .B2(new_n237), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n241), .A2(KEYINPUT81), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n241), .A2(KEYINPUT81), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n251), .B(new_n252), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n283), .A2(new_n286), .A3(KEYINPUT86), .A4(new_n238), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n268), .A2(new_n279), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT87), .ZN(new_n289));
  INV_X1    g103(.A(new_n279), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n283), .A2(new_n286), .A3(new_n238), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n290), .B1(new_n291), .B2(new_n196), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT87), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n293), .A3(new_n287), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  XOR2_X1   g109(.A(new_n279), .B(KEYINPUT85), .Z(new_n296));
  OR2_X1    g110(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n195), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  OAI22_X1  g112(.A1(new_n281), .A2(new_n282), .B1(new_n215), .B2(new_n237), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n279), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT12), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n300), .B(new_n301), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n302), .A2(new_n297), .A3(new_n195), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n187), .B(new_n188), .C1(new_n298), .C2(new_n303), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n297), .A2(new_n195), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(new_n297), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n295), .A2(new_n305), .B1(new_n306), .B2(new_n194), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G469), .ZN(new_n308));
  NAND2_X1  g122(.A1(G469), .A2(G902), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n304), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G214), .B1(G237), .B2(G902), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(G210), .B1(G237), .B2(G902), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G119), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G116), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT69), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT69), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(new_n315), .A3(G116), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT70), .B1(new_n315), .B2(G116), .ZN(new_n321));
  OR3_X1    g135(.A1(new_n315), .A2(KEYINPUT70), .A3(G116), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT2), .B(G113), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(new_n324), .ZN(new_n328));
  OAI221_X1 g142(.A(new_n252), .B1(new_n326), .B2(new_n328), .C1(new_n284), .C2(new_n285), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT5), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(new_n315), .A3(G116), .ZN(new_n331));
  OAI211_X1 g145(.A(G113), .B(new_n331), .C1(new_n327), .C2(new_n330), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n323), .A2(new_n325), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n333), .A3(new_n237), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT88), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT88), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n332), .A2(new_n333), .A3(new_n336), .A4(new_n237), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n329), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(G110), .B(G122), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n329), .A2(new_n339), .A3(new_n335), .A4(new_n337), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT6), .ZN(new_n343));
  INV_X1    g157(.A(G125), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n221), .A2(new_n344), .A3(new_n199), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(new_n251), .B2(new_n344), .ZN(new_n346));
  INV_X1    g160(.A(G224), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n347), .A2(G953), .ZN(new_n348));
  OR2_X1    g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(new_n348), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT6), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n338), .A2(new_n352), .A3(new_n340), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n343), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n332), .A2(new_n333), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n262), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT89), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(new_n334), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n355), .A2(KEYINPUT89), .A3(new_n262), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n339), .B(KEYINPUT8), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT7), .ZN(new_n362));
  INV_X1    g176(.A(new_n348), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n346), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n361), .A2(new_n342), .A3(new_n364), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n349), .A2(new_n350), .B1(new_n362), .B2(new_n363), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n188), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n314), .B1(new_n354), .B2(new_n367), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n361), .A2(new_n342), .A3(new_n364), .ZN(new_n369));
  INV_X1    g183(.A(new_n366), .ZN(new_n370));
  AOI21_X1  g184(.A(G902), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n343), .A2(new_n351), .A3(new_n353), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(new_n313), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n312), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT9), .B(G234), .ZN(new_n375));
  OAI21_X1  g189(.A(G221), .B1(new_n375), .B2(G902), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n310), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G113), .B(G122), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(new_n227), .ZN(new_n379));
  XNOR2_X1  g193(.A(G125), .B(G140), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n206), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT90), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n380), .B(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n381), .B1(new_n383), .B2(new_n206), .ZN(new_n384));
  OR2_X1    g198(.A1(KEYINPUT72), .A2(G953), .ZN(new_n385));
  INV_X1    g199(.A(G237), .ZN(new_n386));
  NAND2_X1  g200(.A1(KEYINPUT72), .A2(G953), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n385), .A2(G214), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n209), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n191), .A2(G143), .A3(G214), .A4(new_n386), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(KEYINPUT18), .A3(G131), .ZN(new_n392));
  NAND2_X1  g206(.A1(KEYINPUT18), .A2(G131), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n389), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n384), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT91), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n395), .B(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(KEYINPUT92), .B1(new_n391), .B2(G131), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT92), .ZN(new_n399));
  AOI211_X1 g213(.A(new_n399), .B(new_n277), .C1(new_n389), .C2(new_n390), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT17), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n380), .A2(KEYINPUT16), .ZN(new_n402));
  OR3_X1    g216(.A1(new_n344), .A2(KEYINPUT16), .A3(G140), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G146), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(new_n403), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n206), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n401), .A2(KEYINPUT93), .A3(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n398), .A2(new_n400), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT17), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n389), .A2(new_n390), .A3(new_n277), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(KEYINPUT93), .B1(new_n401), .B2(new_n408), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n379), .B(new_n397), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n379), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n395), .B(KEYINPUT91), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n380), .A2(KEYINPUT19), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n419), .B1(new_n383), .B2(KEYINPUT19), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n405), .B1(new_n420), .B2(G146), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n410), .B2(new_n412), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n417), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n416), .A2(KEYINPUT94), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT94), .B1(new_n416), .B2(new_n423), .ZN(new_n425));
  NOR2_X1   g239(.A1(G475), .A2(G902), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n424), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT95), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n425), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n416), .A2(KEYINPUT94), .A3(new_n423), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n426), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT95), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n434), .A3(KEYINPUT20), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n416), .A2(new_n423), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n427), .A2(KEYINPUT20), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n430), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n397), .B1(new_n414), .B2(new_n415), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n417), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT96), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n441), .B(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n416), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n188), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G475), .ZN(new_n446));
  INV_X1    g260(.A(G122), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G116), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n230), .B1(new_n448), .B2(KEYINPUT14), .ZN(new_n449));
  XNOR2_X1  g263(.A(G116), .B(G122), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n449), .B(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G128), .B(G143), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT98), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n453), .A2(new_n270), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n453), .A2(new_n270), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n451), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n270), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT97), .B(KEYINPUT13), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(G128), .A3(new_n209), .ZN(new_n459));
  INV_X1    g273(.A(new_n452), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n459), .B(G134), .C1(new_n460), .C2(new_n458), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n450), .B(new_n230), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n457), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n456), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G217), .ZN(new_n465));
  NOR3_X1   g279(.A1(new_n375), .A2(new_n465), .A3(G953), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT100), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n464), .A2(KEYINPUT100), .A3(new_n467), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n456), .A2(new_n463), .A3(new_n466), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT99), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n472), .A2(new_n473), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n470), .B(new_n471), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G478), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(KEYINPUT15), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n476), .A2(new_n188), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n479), .B1(new_n476), .B2(new_n188), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G953), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G952), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n485), .B1(G234), .B2(G237), .ZN(new_n486));
  AOI211_X1 g300(.A(new_n188), .B(new_n191), .C1(G234), .C2(G237), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT21), .B(G898), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n439), .A2(new_n446), .A3(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n377), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n465), .B1(G234), .B2(new_n188), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT79), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n494), .A2(KEYINPUT25), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT22), .B(G137), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n497), .B(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n381), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(new_n404), .B2(G146), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n315), .A2(G128), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n315), .A2(G128), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT24), .B(G110), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n509), .B(new_n504), .C1(new_n502), .C2(KEYINPUT23), .ZN(new_n510));
  OAI22_X1  g324(.A1(new_n506), .A2(new_n508), .B1(new_n510), .B2(G110), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n501), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT77), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n501), .A2(KEYINPUT77), .A3(new_n511), .ZN(new_n515));
  INV_X1    g329(.A(G110), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT76), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n516), .B1(new_n510), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n518), .B1(new_n517), .B2(new_n510), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n405), .A2(new_n407), .B1(new_n506), .B2(new_n508), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n514), .A2(new_n515), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n499), .B1(new_n521), .B2(KEYINPUT78), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(KEYINPUT78), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n520), .A2(new_n519), .ZN(new_n524));
  INV_X1    g338(.A(new_n515), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT77), .B1(new_n501), .B2(new_n511), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT78), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n523), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n522), .B1(new_n530), .B2(new_n499), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n496), .B1(new_n531), .B2(new_n188), .ZN(new_n532));
  INV_X1    g346(.A(new_n499), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n533), .B1(new_n523), .B2(new_n529), .ZN(new_n534));
  NOR4_X1   g348(.A1(new_n534), .A2(G902), .A3(new_n522), .A4(new_n495), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n493), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT80), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n493), .A2(G902), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT80), .B1(new_n534), .B2(new_n522), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT67), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n272), .A3(G134), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT67), .B1(new_n270), .B2(G137), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n272), .A2(G134), .ZN(new_n546));
  OAI211_X1 g360(.A(G131), .B(new_n544), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n278), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n217), .A2(new_n222), .A3(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n326), .A2(new_n328), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n198), .A2(new_n244), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n220), .A2(KEYINPUT65), .A3(new_n246), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT65), .B1(new_n220), .B2(new_n246), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n279), .B(new_n552), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n550), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n548), .B1(new_n221), .B2(new_n199), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(new_n555), .B2(KEYINPUT66), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n249), .A2(new_n250), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT66), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n552), .A4(new_n279), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT30), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n550), .A2(KEYINPUT30), .A3(new_n555), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n551), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n556), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT75), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT31), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n191), .A2(G210), .A3(new_n386), .ZN(new_n569));
  XOR2_X1   g383(.A(KEYINPUT73), .B(KEYINPUT27), .Z(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT26), .B(G101), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n571), .B(new_n572), .Z(new_n573));
  NAND4_X1  g387(.A1(new_n566), .A2(new_n567), .A3(new_n568), .A4(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n555), .A2(KEYINPUT66), .ZN(new_n575));
  INV_X1    g389(.A(new_n557), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n561), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT30), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n550), .A2(KEYINPUT30), .A3(new_n555), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n565), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n556), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n581), .A2(new_n568), .A3(new_n573), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT75), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n574), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n581), .A2(new_n573), .A3(new_n582), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT31), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT74), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT74), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n586), .A2(new_n589), .A3(KEYINPUT31), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n582), .A2(KEYINPUT28), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT28), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n556), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n577), .A2(new_n565), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n573), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n585), .A2(new_n588), .A3(new_n590), .A4(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(G472), .A2(G902), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n599), .A2(KEYINPUT32), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT32), .B1(new_n599), .B2(new_n600), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n550), .A2(new_n555), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n594), .B1(new_n551), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n573), .A2(KEYINPUT29), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT29), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n607), .B1(new_n596), .B2(new_n597), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n566), .A2(new_n573), .ZN(new_n609));
  OAI221_X1 g423(.A(new_n188), .B1(new_n605), .B2(new_n606), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(G472), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n542), .B1(new_n603), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n492), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G101), .ZN(G3));
  INV_X1    g428(.A(new_n472), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT33), .B1(new_n615), .B2(KEYINPUT102), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(KEYINPUT102), .B2(new_n615), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n468), .B(KEYINPUT101), .Z(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n617), .A2(new_n618), .B1(new_n619), .B2(new_n476), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n477), .A2(G902), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n476), .A2(new_n188), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT103), .B(G478), .Z(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n620), .A2(new_n621), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n439), .B2(new_n446), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n599), .A2(new_n188), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n628), .A2(G472), .B1(new_n600), .B2(new_n599), .ZN(new_n629));
  INV_X1    g443(.A(new_n489), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n371), .A2(new_n372), .A3(new_n313), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n313), .B1(new_n371), .B2(new_n372), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n630), .B(new_n311), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(new_n542), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n629), .A2(new_n634), .A3(new_n376), .A4(new_n310), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n627), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT34), .B(G104), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  NOR2_X1   g452(.A1(new_n424), .A2(new_n425), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n437), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n430), .A2(new_n435), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n446), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n635), .A2(new_n482), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT35), .B(G107), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  NOR2_X1   g459(.A1(new_n533), .A2(KEYINPUT36), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n527), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n539), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n536), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n629), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n492), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT37), .B(G110), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  INV_X1    g468(.A(new_n649), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n603), .B2(new_n611), .ZN(new_n656));
  INV_X1    g470(.A(new_n377), .ZN(new_n657));
  INV_X1    g471(.A(G900), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n486), .B1(new_n487), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n641), .A2(new_n446), .A3(new_n483), .A4(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n656), .A2(new_n657), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  AND2_X1   g478(.A1(new_n310), .A2(new_n376), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n659), .B(KEYINPUT39), .Z(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n604), .A2(new_n551), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n597), .B1(new_n670), .B2(new_n556), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(KEYINPUT104), .Z(new_n672));
  INV_X1    g486(.A(new_n586), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n188), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(G472), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n603), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n631), .A2(new_n632), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n677), .A2(KEYINPUT38), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(KEYINPUT38), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n439), .A2(new_n446), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n649), .A2(new_n482), .A3(new_n312), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n668), .A2(new_n669), .A3(new_n676), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G143), .ZN(G45));
  AOI211_X1 g499(.A(new_n625), .B(new_n659), .C1(new_n439), .C2(new_n446), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n656), .A2(new_n686), .A3(new_n657), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  NOR2_X1   g502(.A1(new_n288), .A2(KEYINPUT87), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n293), .B1(new_n292), .B2(new_n287), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n297), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n303), .B1(new_n691), .B2(new_n194), .ZN(new_n692));
  OAI21_X1  g506(.A(G469), .B1(new_n692), .B2(G902), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n693), .A2(new_n376), .A3(new_n304), .ZN(new_n694));
  INV_X1    g508(.A(new_n542), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n588), .A2(new_n590), .A3(new_n598), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n574), .A2(new_n584), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n600), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT32), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n599), .A2(KEYINPUT32), .A3(new_n600), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n611), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n694), .A2(new_n695), .A3(new_n702), .ZN(new_n703));
  AOI211_X1 g517(.A(new_n489), .B(new_n312), .C1(new_n368), .C2(new_n373), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n626), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(KEYINPUT105), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  AOI211_X1 g520(.A(new_n625), .B(new_n633), .C1(new_n439), .C2(new_n446), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n612), .A2(new_n707), .A3(new_n708), .A4(new_n694), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT41), .B(G113), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  AND4_X1   g526(.A1(new_n446), .A2(new_n641), .A3(new_n704), .A4(new_n483), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n612), .A2(new_n713), .A3(new_n694), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  NAND4_X1  g529(.A1(new_n693), .A2(new_n374), .A3(new_n376), .A4(new_n304), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n491), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n656), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  AOI21_X1  g533(.A(new_n482), .B1(new_n439), .B2(new_n446), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n605), .A2(new_n597), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n585), .A2(new_n587), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n600), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(G472), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(new_n599), .B2(new_n188), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n724), .A2(new_n726), .A3(new_n542), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n720), .A2(new_n727), .A3(new_n694), .A4(new_n704), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G122), .ZN(G24));
  INV_X1    g543(.A(new_n726), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n649), .A3(new_n723), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n716), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n686), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  INV_X1    g548(.A(KEYINPUT42), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n308), .A2(KEYINPUT106), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT106), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n307), .A2(new_n737), .A3(G469), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n736), .A2(new_n304), .A3(new_n309), .A4(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n677), .A2(new_n311), .A3(new_n376), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n702), .A2(new_n739), .A3(new_n741), .A4(new_n695), .ZN(new_n742));
  INV_X1    g556(.A(new_n625), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n681), .A2(new_n743), .A3(new_n660), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n735), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n304), .A2(new_n309), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n307), .A2(new_n737), .A3(G469), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n737), .B1(new_n307), .B2(G469), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n740), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n612), .A2(new_n686), .A3(KEYINPUT42), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n745), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G131), .ZN(G33));
  INV_X1    g567(.A(KEYINPUT107), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n754), .B1(new_n742), .B2(new_n661), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n612), .A2(new_n662), .A3(new_n750), .A4(KEYINPUT107), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g571(.A(KEYINPUT108), .B(G134), .Z(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G36));
  NOR2_X1   g573(.A1(new_n681), .A2(new_n625), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT43), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n629), .A2(new_n655), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n376), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n692), .A2(G469), .A3(G902), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n295), .A2(new_n305), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n306), .A2(new_n194), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n307), .A2(KEYINPUT45), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(G469), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n309), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT46), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n767), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n774), .A2(KEYINPUT46), .A3(new_n309), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n766), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n631), .A2(new_n632), .A3(new_n312), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n779), .A2(new_n666), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n761), .A2(KEYINPUT44), .A3(new_n762), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n765), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  XOR2_X1   g597(.A(KEYINPUT109), .B(G137), .Z(new_n784));
  XNOR2_X1  g598(.A(new_n783), .B(new_n784), .ZN(G39));
  NAND2_X1  g599(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n779), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n780), .A2(new_n542), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n744), .A2(new_n702), .A3(new_n788), .ZN(new_n789));
  XOR2_X1   g603(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n790));
  OAI211_X1 g604(.A(new_n787), .B(new_n789), .C1(new_n779), .C2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G140), .ZN(G42));
  INV_X1    g606(.A(new_n716), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n761), .A2(new_n794), .A3(new_n486), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n794), .B1(new_n761), .B2(new_n486), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n793), .B(new_n727), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n694), .A2(new_n780), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n695), .A2(new_n486), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n798), .A2(new_n676), .A3(new_n799), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n800), .B(KEYINPUT117), .Z(new_n801));
  AOI21_X1  g615(.A(new_n485), .B1(new_n801), .B2(new_n626), .ZN(new_n802));
  INV_X1    g616(.A(new_n798), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n612), .B(new_n803), .C1(new_n795), .C2(new_n796), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n804), .A2(KEYINPUT48), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(KEYINPUT48), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n797), .B(new_n802), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n694), .A2(new_n312), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n808), .A2(KEYINPUT115), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(KEYINPUT115), .ZN(new_n810));
  NOR2_X1   g624(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n809), .A2(new_n810), .A3(new_n680), .A4(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n727), .B(new_n812), .C1(new_n795), .C2(new_n796), .ZN(new_n813));
  AND2_X1   g627(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n779), .A2(new_n790), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n816), .B1(new_n779), .B2(new_n786), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n693), .A2(new_n304), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n817), .B1(new_n766), .B2(new_n818), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n727), .B(new_n780), .C1(new_n795), .C2(new_n796), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT51), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n815), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n681), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n801), .A2(new_n823), .A3(new_n625), .ZN(new_n824));
  INV_X1    g638(.A(new_n731), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n825), .B(new_n803), .C1(new_n795), .C2(new_n796), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT118), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n807), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n817), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n818), .A2(new_n766), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n833), .B1(new_n817), .B2(new_n831), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n826), .B(new_n824), .C1(new_n835), .C2(new_n820), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n830), .B1(new_n836), .B2(new_n815), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n829), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n536), .A2(new_n376), .A3(new_n648), .A4(new_n660), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(new_n746), .B2(new_n749), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n840), .A2(new_n676), .A3(new_n374), .A4(new_n720), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n663), .A2(new_n687), .A3(new_n733), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT52), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n702), .A2(new_n649), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n377), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n845), .A2(new_n662), .B1(new_n686), .B2(new_n732), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n846), .A2(new_n847), .A3(new_n687), .A4(new_n841), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n686), .A2(new_n825), .A3(new_n750), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT112), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n480), .A2(new_n481), .A3(new_n659), .ZN(new_n852));
  AND4_X1   g666(.A1(new_n311), .A2(new_n852), .A3(new_n368), .A4(new_n373), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n310), .A2(new_n376), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(new_n642), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n851), .B1(new_n855), .B2(new_n656), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n844), .A2(new_n854), .A3(KEYINPUT112), .A4(new_n642), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n850), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n745), .A2(new_n751), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n702), .A2(new_n695), .ZN(new_n861));
  AOI211_X1 g675(.A(new_n491), .B(new_n377), .C1(new_n861), .C2(new_n650), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n439), .A2(new_n446), .A3(new_n483), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n635), .B1(new_n627), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT111), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n492), .B1(new_n612), .B2(new_n651), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n634), .A2(new_n310), .A3(new_n376), .ZN(new_n867));
  INV_X1    g681(.A(new_n863), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n867), .B(new_n629), .C1(new_n868), .C2(new_n626), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT111), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n866), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n865), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n714), .A2(new_n718), .A3(new_n728), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n873), .B1(new_n709), .B2(new_n706), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n860), .A2(new_n872), .A3(new_n757), .A4(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n876));
  INV_X1    g690(.A(new_n846), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT52), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n849), .B(new_n875), .C1(new_n876), .C2(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n714), .A2(new_n718), .A3(new_n728), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n866), .A2(new_n869), .A3(new_n870), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n870), .B1(new_n866), .B2(new_n869), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n710), .B(new_n880), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n855), .A2(new_n656), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT112), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n855), .A2(new_n851), .A3(new_n656), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n887), .A2(new_n752), .A3(new_n757), .A4(new_n850), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n843), .A2(new_n848), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT53), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT54), .B1(new_n879), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n876), .B1(new_n875), .B2(new_n849), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT54), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n880), .A2(new_n710), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n865), .B2(new_n871), .ZN(new_n896));
  INV_X1    g710(.A(new_n888), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n876), .B1(new_n877), .B2(KEYINPUT52), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n896), .A2(new_n890), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n893), .A2(new_n894), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n892), .A2(new_n900), .ZN(new_n901));
  OAI22_X1  g715(.A1(new_n838), .A2(new_n901), .B1(G952), .B2(G953), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n695), .A2(new_n311), .A3(new_n376), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT49), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n903), .B(new_n680), .C1(new_n904), .C2(new_n818), .ZN(new_n905));
  INV_X1    g719(.A(new_n676), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n818), .A2(new_n904), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n905), .A2(new_n906), .A3(new_n760), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n902), .A2(new_n908), .ZN(G75));
  NAND2_X1  g723(.A1(new_n893), .A2(new_n899), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n910), .A2(G210), .A3(G902), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT56), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n343), .A2(new_n353), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT119), .Z(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT55), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(new_n351), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n911), .A2(new_n912), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n916), .B1(new_n911), .B2(new_n912), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n191), .A2(G952), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(G51));
  AOI211_X1 g734(.A(new_n188), .B(new_n774), .C1(new_n893), .C2(new_n899), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n309), .B(KEYINPUT57), .Z(new_n922));
  AND3_X1   g736(.A1(new_n893), .A2(new_n894), .A3(new_n899), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n894), .B1(new_n893), .B2(new_n899), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n692), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n921), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT120), .B1(new_n927), .B2(new_n919), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT120), .ZN(new_n929));
  INV_X1    g743(.A(new_n919), .ZN(new_n930));
  AND4_X1   g744(.A1(new_n896), .A2(new_n890), .A3(new_n897), .A4(new_n898), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT54), .B1(new_n891), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n900), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n692), .B1(new_n933), .B2(new_n922), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n929), .B(new_n930), .C1(new_n934), .C2(new_n921), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n928), .A2(new_n935), .ZN(G54));
  NAND4_X1  g750(.A1(new_n910), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n937));
  INV_X1    g751(.A(new_n639), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(new_n919), .ZN(G60));
  NAND2_X1  g755(.A1(G478), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT59), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n620), .B1(new_n901), .B2(new_n943), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n933), .A2(new_n620), .A3(new_n943), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n944), .A2(new_n919), .A3(new_n945), .ZN(G63));
  NAND2_X1  g760(.A1(G217), .A2(G902), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT121), .Z(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT60), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n893), .B2(new_n899), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n647), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n538), .A2(new_n540), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n951), .B(new_n930), .C1(new_n952), .C2(new_n950), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT122), .ZN(new_n954));
  AOI21_X1  g768(.A(KEYINPUT61), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n953), .B(new_n955), .ZN(G66));
  INV_X1    g770(.A(new_n488), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n484), .B1(new_n957), .B2(G224), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n958), .B1(new_n883), .B2(new_n191), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n914), .B1(G898), .B2(new_n191), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT123), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n959), .B(new_n961), .ZN(G69));
  XOR2_X1   g776(.A(new_n564), .B(new_n420), .Z(new_n963));
  INV_X1    g777(.A(new_n191), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(G900), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n720), .A2(new_n374), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n779), .A2(new_n612), .A3(new_n666), .A4(new_n966), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n791), .A2(new_n752), .A3(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n687), .A2(new_n663), .A3(new_n733), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n968), .A2(new_n757), .A3(new_n783), .A4(new_n969), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n963), .B(new_n965), .C1(new_n970), .C2(new_n964), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT124), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n684), .A2(new_n969), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT62), .ZN(new_n974));
  INV_X1    g788(.A(new_n667), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n627), .A2(new_n863), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n975), .A2(new_n612), .A3(new_n976), .A4(new_n780), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n791), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n783), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n972), .B1(new_n974), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT62), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n973), .B(new_n981), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n982), .A2(KEYINPUT124), .A3(new_n783), .A4(new_n978), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n964), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n971), .B1(new_n984), .B2(new_n963), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n191), .B1(G227), .B2(G900), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(G72));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT63), .ZN(new_n989));
  INV_X1    g803(.A(new_n609), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n989), .B1(new_n990), .B2(new_n586), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n991), .B1(new_n879), .B2(new_n891), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT127), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n989), .B(KEYINPUT125), .Z(new_n994));
  OAI21_X1  g808(.A(new_n994), .B1(new_n970), .B2(new_n883), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n566), .A2(new_n597), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n993), .B1(new_n997), .B2(new_n930), .ZN(new_n998));
  AOI211_X1 g812(.A(KEYINPUT127), .B(new_n919), .C1(new_n995), .C2(new_n996), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n992), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n980), .A2(new_n983), .A3(new_n896), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n994), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n566), .A2(new_n597), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(KEYINPUT126), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT126), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1002), .A2(new_n1006), .A3(new_n1003), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1000), .B1(new_n1005), .B2(new_n1007), .ZN(G57));
endmodule


