//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n582, new_n583, new_n585, new_n586, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n641, new_n642, new_n643, new_n644,
    new_n647, new_n648, new_n650, new_n651, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  INV_X1    g031(.A(G2104), .ZN(new_n457));
  OAI21_X1  g032(.A(KEYINPUT67), .B1(new_n457), .B2(G2105), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n459));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n459), .A2(new_n460), .A3(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n460), .A2(G137), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n462), .A2(G101), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OR2_X1    g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  AND2_X1   g048(.A1(new_n463), .A2(KEYINPUT68), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n463), .A2(KEYINPUT68), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n460), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT69), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(G112), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G2105), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n476), .A2(G2105), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G136), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  AND2_X1   g061(.A1(G126), .A2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n463), .A2(new_n487), .ZN(new_n488));
  OR2_X1    g063(.A1(new_n460), .A2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n460), .A2(G138), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(new_n463), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n463), .A2(new_n494), .A3(new_n495), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n493), .B1(new_n497), .B2(new_n498), .ZN(G164));
  NOR2_X1   g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  OAI22_X1  g078(.A1(new_n500), .A2(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G88), .ZN(new_n505));
  OAI21_X1  g080(.A(G543), .B1(new_n502), .B2(new_n503), .ZN(new_n506));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  OAI22_X1  g082(.A1(new_n504), .A2(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI221_X1 g085(.A(KEYINPUT70), .B1(new_n506), .B2(new_n507), .C1(new_n504), .C2(new_n505), .ZN(new_n511));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n501), .A2(new_n500), .ZN(new_n513));
  INV_X1    g088(.A(G62), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n510), .A2(new_n511), .B1(G651), .B2(new_n515), .ZN(G166));
  OAI21_X1  g091(.A(KEYINPUT71), .B1(new_n501), .B2(new_n500), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT72), .B(KEYINPUT7), .Z(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n526), .B(new_n527), .ZN(new_n528));
  OR2_X1    g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n519), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G51), .ZN(new_n532));
  INV_X1    g107(.A(new_n504), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G89), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n525), .A2(new_n528), .A3(new_n532), .A4(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  NAND3_X1  g111(.A1(new_n517), .A2(new_n523), .A3(G64), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G651), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  XNOR2_X1  g116(.A(KEYINPUT73), .B(G52), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n504), .A2(new_n541), .B1(new_n506), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n540), .A2(KEYINPUT74), .A3(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT74), .ZN(new_n546));
  INV_X1    g121(.A(G651), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n537), .B2(new_n538), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n548), .B2(new_n543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n545), .A2(new_n549), .ZN(G171));
  OAI211_X1 g125(.A(G43), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n551));
  XOR2_X1   g126(.A(KEYINPUT75), .B(G81), .Z(new_n552));
  OAI211_X1 g127(.A(KEYINPUT76), .B(new_n551), .C1(new_n504), .C2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n529), .A2(new_n530), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n520), .A2(new_n522), .ZN(new_n556));
  XNOR2_X1  g131(.A(KEYINPUT75), .B(G81), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g133(.A(KEYINPUT76), .B1(new_n558), .B2(new_n551), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n517), .A2(new_n523), .A3(G56), .ZN(new_n561));
  NAND2_X1  g136(.A1(G68), .A2(G543), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n547), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(new_n520), .B2(new_n522), .ZN(new_n571));
  AND2_X1   g146(.A1(G78), .A2(G543), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n555), .A2(new_n556), .A3(G91), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(KEYINPUT77), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(new_n531), .B2(G53), .ZN(new_n578));
  OAI211_X1 g153(.A(G53), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n576), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n573), .B(new_n574), .C1(new_n578), .C2(new_n580), .ZN(G299));
  AND3_X1   g156(.A1(new_n545), .A2(KEYINPUT78), .A3(new_n549), .ZN(new_n582));
  AOI21_X1  g157(.A(KEYINPUT78), .B1(new_n545), .B2(new_n549), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(G301));
  NAND2_X1  g159(.A1(new_n510), .A2(new_n511), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n515), .A2(G651), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(G303));
  NAND2_X1  g162(.A1(new_n517), .A2(new_n523), .ZN(new_n588));
  INV_X1    g163(.A(G74), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n547), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(G87), .ZN(new_n591));
  INV_X1    g166(.A(G49), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n504), .A2(new_n591), .B1(new_n506), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G288));
  OAI21_X1  g170(.A(G61), .B1(new_n501), .B2(new_n500), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  AOI211_X1 g172(.A(KEYINPUT79), .B(new_n547), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(G86), .ZN(new_n599));
  INV_X1    g174(.A(G48), .ZN(new_n600));
  OAI22_X1  g175(.A1(new_n504), .A2(new_n599), .B1(new_n506), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n596), .A2(new_n597), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G651), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n602), .A2(new_n606), .ZN(G305));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n517), .A2(new_n523), .A3(G60), .ZN(new_n609));
  NAND2_X1  g184(.A1(G72), .A2(G543), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G651), .ZN(new_n612));
  INV_X1    g187(.A(G85), .ZN(new_n613));
  INV_X1    g188(.A(G47), .ZN(new_n614));
  OAI22_X1  g189(.A1(new_n504), .A2(new_n613), .B1(new_n506), .B2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n608), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n547), .B1(new_n609), .B2(new_n610), .ZN(new_n618));
  NOR3_X1   g193(.A1(new_n618), .A2(KEYINPUT80), .A3(new_n615), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(G290));
  INV_X1    g196(.A(G66), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(new_n520), .B2(new_n522), .ZN(new_n623));
  NAND2_X1  g198(.A1(G79), .A2(G543), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(KEYINPUT81), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n627), .B(new_n624), .C1(new_n513), .C2(new_n622), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n626), .A2(G651), .A3(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT10), .ZN(new_n630));
  INV_X1    g205(.A(G92), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n504), .B2(new_n631), .ZN(new_n632));
  NAND4_X1  g207(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT10), .A4(G92), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n531), .A2(G54), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n629), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n636), .A2(G868), .ZN(new_n637));
  INV_X1    g212(.A(G301), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(G868), .ZN(G284));
  AOI21_X1  g214(.A(new_n637), .B1(new_n638), .B2(G868), .ZN(G321));
  NAND2_X1  g215(.A1(G286), .A2(G868), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n578), .A2(new_n580), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n573), .A2(new_n574), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n641), .B1(G868), .B2(new_n644), .ZN(G297));
  XNOR2_X1  g220(.A(G297), .B(KEYINPUT82), .ZN(G280));
  INV_X1    g221(.A(new_n636), .ZN(new_n647));
  INV_X1    g222(.A(G559), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n647), .B1(new_n648), .B2(G860), .ZN(G148));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(G868), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(G868), .B2(new_n564), .ZN(G323));
  XNOR2_X1  g227(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g228(.A1(new_n483), .A2(G135), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n477), .A2(G123), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n460), .A2(G111), .ZN(new_n656));
  OAI21_X1  g231(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n654), .B(new_n655), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(G2096), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n462), .A2(new_n463), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT12), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT13), .Z(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(G2100), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(G2100), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n659), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT83), .ZN(G156));
  XOR2_X1   g241(.A(G2443), .B(G2446), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT85), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2451), .ZN(new_n669));
  XOR2_X1   g244(.A(G1341), .B(G1348), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT15), .B(G2435), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2438), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2427), .B(G2430), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT86), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n676), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n677), .A2(new_n678), .A3(KEYINPUT14), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n671), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(G2454), .Z(new_n682));
  OR2_X1    g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n682), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n683), .A2(G14), .A3(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G401));
  XNOR2_X1  g261(.A(G2084), .B(G2090), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT87), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G2067), .B(G2678), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT88), .ZN(new_n691));
  XNOR2_X1  g266(.A(G2072), .B(G2078), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT17), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n689), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(new_n692), .B2(new_n691), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT90), .Z(new_n696));
  NAND3_X1  g271(.A1(new_n689), .A2(new_n692), .A3(new_n691), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n697), .B(new_n698), .Z(new_n699));
  OR3_X1    g274(.A1(new_n691), .A2(new_n688), .A3(new_n693), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n696), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G2096), .B(G2100), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G227));
  XNOR2_X1  g279(.A(G1971), .B(G1976), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT19), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(G1961), .B(G1966), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT91), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1956), .B(G2474), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n707), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT20), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n707), .B1(new_n709), .B2(new_n711), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n709), .A2(new_n711), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n713), .B(new_n716), .C1(new_n706), .C2(new_n715), .ZN(new_n717));
  XNOR2_X1  g292(.A(G1991), .B(G1996), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT92), .ZN(new_n721));
  XNOR2_X1  g296(.A(G1981), .B(G1986), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT93), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n721), .B(new_n723), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n719), .A2(new_n724), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(G229));
  INV_X1    g302(.A(G16), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G23), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n594), .B2(new_n728), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT33), .B(G1976), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NOR3_X1   g307(.A1(new_n605), .A2(new_n598), .A3(new_n601), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G16), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G6), .B2(G16), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT32), .B(G1981), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n732), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n728), .A2(KEYINPUT96), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n728), .A2(KEYINPUT96), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G22), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT97), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G166), .B2(new_n742), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G1971), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n736), .A2(new_n737), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n745), .A2(G1971), .ZN(new_n748));
  AND4_X1   g323(.A1(new_n738), .A2(new_n746), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT34), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  INV_X1    g327(.A(G29), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G25), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT94), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n483), .A2(G131), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n477), .A2(G119), .ZN(new_n757));
  INV_X1    g332(.A(G95), .ZN(new_n758));
  AND3_X1   g333(.A1(new_n758), .A2(new_n460), .A3(KEYINPUT95), .ZN(new_n759));
  AOI21_X1  g334(.A(KEYINPUT95), .B1(new_n758), .B2(new_n460), .ZN(new_n760));
  OAI221_X1 g335(.A(G2104), .B1(G107), .B2(new_n460), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n756), .A2(new_n757), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n755), .B1(new_n762), .B2(G29), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT35), .B(G1991), .Z(new_n764));
  XOR2_X1   g339(.A(new_n763), .B(new_n764), .Z(new_n765));
  NOR2_X1   g340(.A1(new_n741), .A2(G24), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n620), .B2(new_n741), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(G1986), .Z(new_n768));
  NAND4_X1  g343(.A1(new_n751), .A2(new_n752), .A3(new_n765), .A4(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT36), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n753), .A2(G35), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G162), .B2(new_n753), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G2090), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT105), .B(KEYINPUT29), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G5), .A2(G16), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G171), .B2(G16), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1961), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n483), .A2(G139), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT100), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n463), .A2(G127), .ZN(new_n782));
  INV_X1    g357(.A(G115), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n457), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT101), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n460), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n785), .B2(new_n784), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT25), .Z(new_n789));
  NAND3_X1  g364(.A1(new_n781), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(G29), .ZN(new_n792));
  NOR2_X1   g367(.A1(G29), .A2(G33), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT99), .Z(new_n794));
  AOI22_X1  g369(.A1(new_n792), .A2(new_n794), .B1(KEYINPUT102), .B2(G2072), .ZN(new_n795));
  OR3_X1    g370(.A1(new_n795), .A2(KEYINPUT102), .A3(G2072), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(KEYINPUT102), .B2(G2072), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n779), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(G168), .A2(new_n728), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n728), .B2(G21), .ZN(new_n800));
  INV_X1    g375(.A(G1966), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT104), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n753), .A2(G26), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT28), .Z(new_n805));
  NAND2_X1  g380(.A1(new_n483), .A2(G140), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n477), .A2(G128), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n460), .A2(G116), .ZN(new_n808));
  OAI21_X1  g383(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n806), .B(new_n807), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n805), .B1(new_n810), .B2(G29), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G2067), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n742), .A2(G19), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT98), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n564), .B2(new_n742), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G1341), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n728), .A2(G4), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n647), .B2(new_n728), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G1348), .ZN(new_n819));
  NOR4_X1   g394(.A1(new_n803), .A2(new_n812), .A3(new_n816), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n753), .A2(G32), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n483), .A2(G141), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n477), .A2(G129), .ZN(new_n823));
  NAND3_X1  g398(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT26), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  AOI22_X1  g402(.A1(G105), .A2(new_n462), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n822), .A2(new_n823), .A3(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n821), .B1(new_n830), .B2(new_n753), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT27), .B(G1996), .Z(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT103), .ZN(new_n834));
  INV_X1    g409(.A(G28), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n835), .A2(KEYINPUT30), .ZN(new_n836));
  AOI21_X1  g411(.A(G29), .B1(new_n835), .B2(KEYINPUT30), .ZN(new_n837));
  OR2_X1    g412(.A1(KEYINPUT31), .A2(G11), .ZN(new_n838));
  NAND2_X1  g413(.A1(KEYINPUT31), .A2(G11), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n836), .A2(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI221_X1 g415(.A(new_n840), .B1(new_n753), .B2(new_n658), .C1(new_n800), .C2(new_n801), .ZN(new_n841));
  INV_X1    g416(.A(G34), .ZN(new_n842));
  AOI21_X1  g417(.A(G29), .B1(new_n842), .B2(KEYINPUT24), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(KEYINPUT24), .B2(new_n842), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n472), .B2(new_n753), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(G2084), .Z(new_n846));
  NOR2_X1   g421(.A1(G27), .A2(G29), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(G164), .B2(G29), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(G2078), .ZN(new_n849));
  NOR3_X1   g424(.A1(new_n841), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n742), .A2(G20), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT23), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n644), .B2(new_n728), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(G1956), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(new_n831), .B2(new_n832), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n834), .A2(new_n850), .A3(new_n855), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n776), .A2(new_n798), .A3(new_n820), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n771), .A2(new_n857), .ZN(G311));
  OR2_X1    g433(.A1(new_n771), .A2(new_n857), .ZN(G150));
  INV_X1    g434(.A(G93), .ZN(new_n860));
  INV_X1    g435(.A(G55), .ZN(new_n861));
  OAI22_X1  g436(.A1(new_n504), .A2(new_n860), .B1(new_n506), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(G80), .A2(G543), .ZN(new_n863));
  INV_X1    g438(.A(G67), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n588), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n862), .B1(new_n865), .B2(G651), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(G860), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT107), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT37), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT106), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n560), .B2(new_n563), .ZN(new_n872));
  INV_X1    g447(.A(new_n563), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n873), .B(KEYINPUT106), .C1(new_n559), .C2(new_n554), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n867), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n564), .A2(KEYINPUT106), .A3(new_n866), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n647), .A2(G559), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n881), .A2(KEYINPUT39), .ZN(new_n882));
  INV_X1    g457(.A(G860), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(new_n881), .B2(KEYINPUT39), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n870), .B1(new_n882), .B2(new_n884), .ZN(G145));
  XNOR2_X1  g460(.A(new_n658), .B(G160), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n485), .ZN(new_n887));
  AOI22_X1  g462(.A1(new_n463), .A2(new_n487), .B1(new_n489), .B2(new_n491), .ZN(new_n888));
  INV_X1    g463(.A(new_n498), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n888), .B1(new_n889), .B2(new_n496), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT108), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g467(.A(KEYINPUT108), .B(new_n888), .C1(new_n889), .C2(new_n496), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n810), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n810), .A2(new_n894), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n895), .A2(new_n829), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n829), .B1(new_n895), .B2(new_n896), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n790), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n810), .B(new_n894), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n830), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n895), .A2(new_n829), .A3(new_n896), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n791), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n904));
  INV_X1    g479(.A(G118), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n904), .B1(new_n905), .B2(G2105), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n906), .B1(new_n477), .B2(G130), .ZN(new_n907));
  INV_X1    g482(.A(G142), .ZN(new_n908));
  INV_X1    g483(.A(new_n483), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n661), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n762), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n907), .B(new_n661), .C1(new_n908), .C2(new_n909), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n913), .B1(new_n912), .B2(new_n914), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n899), .A2(new_n903), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT109), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n899), .A2(new_n903), .ZN(new_n921));
  INV_X1    g496(.A(new_n917), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n919), .A3(new_n922), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n887), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT40), .ZN(new_n927));
  INV_X1    g502(.A(G37), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n918), .A2(new_n887), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n917), .B1(new_n899), .B2(new_n903), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n926), .A2(new_n927), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n887), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n930), .B1(new_n919), .B2(new_n918), .ZN(new_n934));
  INV_X1    g509(.A(new_n925), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n931), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT40), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n932), .A2(new_n938), .ZN(G395));
  XNOR2_X1  g514(.A(new_n877), .B(new_n650), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n636), .A2(new_n644), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT110), .ZN(new_n942));
  NAND4_X1  g517(.A1(G299), .A2(new_n629), .A3(new_n635), .A4(new_n634), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n647), .A2(KEYINPUT110), .A3(G299), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n940), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT41), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n949), .B1(new_n944), .B2(new_n945), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n941), .A2(new_n943), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n951), .B1(new_n952), .B2(new_n949), .ZN(new_n953));
  AOI211_X1 g528(.A(KEYINPUT111), .B(KEYINPUT41), .C1(new_n941), .C2(new_n943), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n950), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n948), .B1(new_n955), .B2(new_n940), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n956), .A2(KEYINPUT42), .ZN(new_n957));
  OAI21_X1  g532(.A(G166), .B1(new_n617), .B2(new_n619), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT80), .B1(new_n618), .B2(new_n615), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n612), .A2(new_n608), .A3(new_n616), .ZN(new_n960));
  NAND3_X1  g535(.A1(G303), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n962));
  INV_X1    g537(.A(new_n593), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT112), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n590), .A2(new_n965), .A3(new_n593), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n733), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n962), .A2(new_n963), .A3(KEYINPUT112), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n965), .B1(new_n590), .B2(new_n593), .ZN(new_n969));
  NAND3_X1  g544(.A1(G305), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  AND4_X1   g545(.A1(new_n958), .A2(new_n961), .A3(new_n967), .A4(new_n970), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n958), .A2(new_n961), .B1(new_n967), .B2(new_n970), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n956), .A2(KEYINPUT42), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n957), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n973), .B1(new_n957), .B2(new_n974), .ZN(new_n976));
  OAI21_X1  g551(.A(G868), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(G868), .B2(new_n866), .ZN(G295));
  OAI21_X1  g553(.A(new_n977), .B1(G868), .B2(new_n866), .ZN(G331));
  INV_X1    g554(.A(KEYINPUT78), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT74), .B1(new_n540), .B2(new_n544), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n548), .A2(new_n546), .A3(new_n543), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n545), .A2(KEYINPUT78), .A3(new_n549), .ZN(new_n984));
  AOI21_X1  g559(.A(G286), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(G171), .A2(G168), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n876), .B(new_n875), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(G168), .B1(new_n582), .B2(new_n583), .ZN(new_n988));
  INV_X1    g563(.A(new_n986), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(new_n877), .A3(new_n989), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n987), .A2(KEYINPUT41), .A3(new_n990), .A4(new_n952), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(new_n971), .B2(new_n972), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n958), .A2(new_n961), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n967), .A2(new_n970), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n958), .A2(new_n961), .A3(new_n967), .A4(new_n970), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(KEYINPUT113), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n993), .A2(new_n998), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n991), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n987), .A2(KEYINPUT41), .A3(new_n990), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n946), .ZN(new_n1002));
  AOI21_X1  g577(.A(G37), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n988), .A2(new_n877), .A3(new_n989), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n877), .B1(new_n988), .B2(new_n989), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n946), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n955), .A2(new_n987), .A3(new_n990), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT114), .B1(new_n1008), .B2(new_n973), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n1010));
  INV_X1    g585(.A(new_n973), .ZN(new_n1011));
  AOI211_X1 g586(.A(new_n1010), .B(new_n1011), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1003), .B(KEYINPUT43), .C1(new_n1009), .C2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1006), .A2(new_n1007), .A3(new_n999), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n928), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n955), .A2(new_n987), .A3(new_n990), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n947), .B1(new_n987), .B2(new_n990), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n973), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n1010), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1008), .A2(KEYINPUT114), .A3(new_n973), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1015), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1013), .B1(new_n1021), .B2(KEYINPUT43), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT44), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT43), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1003), .B(new_n1024), .C1(new_n1009), .C2(new_n1012), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1023), .A2(new_n1028), .ZN(G397));
  XOR2_X1   g604(.A(new_n762), .B(new_n764), .Z(new_n1030));
  INV_X1    g605(.A(G1384), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n894), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT45), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n465), .A2(new_n471), .A3(G40), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1030), .A2(new_n1036), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1035), .A2(G1996), .A3(new_n829), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1036), .A2(G1996), .A3(new_n829), .ZN(new_n1039));
  OR2_X1    g614(.A1(new_n1039), .A2(KEYINPUT115), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(KEYINPUT115), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1038), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n810), .B(G2067), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n1036), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1044), .B(KEYINPUT116), .ZN(new_n1045));
  AND2_X1   g620(.A1(G290), .A2(G1986), .ZN(new_n1046));
  NOR2_X1   g621(.A1(G290), .A2(G1986), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1036), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AND4_X1   g623(.A1(new_n1037), .A2(new_n1042), .A3(new_n1045), .A4(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(G303), .A2(KEYINPUT118), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1050));
  INV_X1    g625(.A(G8), .ZN(new_n1051));
  NOR2_X1   g626(.A1(G166), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1050), .B1(KEYINPUT55), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT118), .B1(new_n1052), .B2(KEYINPUT55), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1033), .A2(G1384), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n892), .A2(new_n893), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n890), .A2(new_n1031), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n1033), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1057), .A2(new_n1059), .A3(new_n1034), .ZN(new_n1060));
  INV_X1    g635(.A(G1971), .ZN(new_n1061));
  NOR2_X1   g636(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n890), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n1034), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT50), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(new_n890), .B2(new_n1031), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT117), .B(G2090), .Z(new_n1068));
  AOI22_X1  g643(.A1(new_n1060), .A2(new_n1061), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1055), .B1(new_n1069), .B2(new_n1051), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G305), .A2(G1981), .ZN(new_n1071));
  INV_X1    g646(.A(G1981), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n733), .A2(new_n1072), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1071), .A2(new_n1073), .A3(KEYINPUT49), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT49), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1034), .A2(new_n1031), .A3(new_n890), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G8), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n594), .A2(G1976), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(G8), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT52), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1082), .B1(new_n594), .B2(G1976), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1081), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1078), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1088), .B(G8), .C1(new_n1054), .C2(new_n1053), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1056), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1034), .B1(G164), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT45), .B1(new_n890), .B2(new_n1031), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n801), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1058), .A2(KEYINPUT50), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n465), .A2(new_n471), .A3(G40), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1095), .B1(new_n890), .B2(new_n1062), .ZN(new_n1096));
  XOR2_X1   g671(.A(KEYINPUT119), .B(G2084), .Z(new_n1097));
  NAND3_X1  g672(.A1(new_n1094), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1093), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(G8), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(G286), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1070), .A2(new_n1085), .A3(new_n1089), .A4(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT120), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT63), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT63), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1102), .A2(KEYINPUT120), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1089), .ZN(new_n1108));
  OR2_X1    g683(.A1(G288), .A2(G1976), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1073), .B1(new_n1078), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1077), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1108), .A2(new_n1085), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1070), .A2(new_n1085), .A3(new_n1089), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(new_n1060), .B2(G2078), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1116));
  INV_X1    g691(.A(G1961), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1114), .A2(G2078), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1115), .A2(new_n1118), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(G301), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT54), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1057), .A2(new_n1034), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(new_n1126), .A3(new_n1120), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1127), .A2(new_n1115), .A3(new_n1118), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1124), .B1(new_n1128), .B2(G171), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1113), .B1(new_n1123), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1076), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT58), .B(G1341), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1060), .A2(G1996), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n564), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT59), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1133), .A2(new_n1136), .A3(new_n564), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(G1956), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1116), .A2(new_n1139), .ZN(new_n1140));
  XOR2_X1   g715(.A(G299), .B(KEYINPUT57), .Z(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT56), .B(G2072), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1140), .B(new_n1141), .C1(new_n1060), .C2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1146), .B1(new_n1147), .B2(new_n1144), .ZN(new_n1148));
  AOI21_X1  g723(.A(G1348), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1076), .A2(G2067), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n636), .B1(new_n1151), .B2(KEYINPUT60), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n1153));
  NOR4_X1   g728(.A1(new_n1149), .A2(new_n1150), .A3(new_n1153), .A4(new_n647), .ZN(new_n1154));
  OAI22_X1  g729(.A1(new_n1152), .A2(new_n1154), .B1(KEYINPUT60), .B2(new_n1151), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1138), .A2(new_n1148), .A3(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1126), .A2(new_n1059), .A3(new_n1142), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1141), .B1(new_n1157), .B2(new_n1140), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1151), .A2(new_n636), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1144), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1156), .A2(new_n1160), .ZN(new_n1161));
  XOR2_X1   g736(.A(KEYINPUT125), .B(KEYINPUT54), .Z(new_n1162));
  NOR2_X1   g737(.A1(new_n1128), .A2(new_n638), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1122), .A2(G301), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1162), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1130), .A2(new_n1161), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1099), .A2(KEYINPUT122), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT122), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1093), .A2(new_n1098), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(G168), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT51), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1172), .A2(new_n1051), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1171), .A2(KEYINPUT124), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n1175));
  AOI21_X1  g750(.A(G286), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1173), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n1100), .B(new_n1172), .C1(new_n1051), .C2(G168), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1174), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1167), .A2(G8), .A3(G286), .A4(new_n1169), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1181), .B(new_n1182), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g759(.A(new_n1107), .B(new_n1112), .C1(new_n1166), .C2(new_n1184), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1164), .A2(new_n1070), .A3(new_n1085), .A4(new_n1089), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1180), .A2(KEYINPUT62), .A3(new_n1183), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1186), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1049), .B1(new_n1185), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n913), .A2(new_n764), .ZN(new_n1193));
  XOR2_X1   g768(.A(new_n1193), .B(KEYINPUT126), .Z(new_n1194));
  NAND3_X1  g769(.A1(new_n1042), .A2(new_n1045), .A3(new_n1194), .ZN(new_n1195));
  OR2_X1    g770(.A1(new_n810), .A2(G2067), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1035), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  OR2_X1    g772(.A1(new_n1043), .A2(new_n829), .ZN(new_n1198));
  OR3_X1    g773(.A1(new_n1035), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1199));
  OAI21_X1  g774(.A(KEYINPUT46), .B1(new_n1035), .B2(G1996), .ZN(new_n1200));
  AOI22_X1  g775(.A1(new_n1198), .A2(new_n1036), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT47), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1036), .A2(new_n1047), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1203), .B(KEYINPUT48), .ZN(new_n1204));
  AND4_X1   g779(.A1(new_n1037), .A2(new_n1042), .A3(new_n1045), .A4(new_n1204), .ZN(new_n1205));
  NOR3_X1   g780(.A1(new_n1197), .A2(new_n1202), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1192), .A2(new_n1206), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g782(.A1(new_n685), .A2(new_n726), .A3(new_n725), .ZN(new_n1209));
  NAND2_X1  g783(.A1(new_n703), .A2(G319), .ZN(new_n1210));
  OR2_X1    g784(.A1(new_n1210), .A2(KEYINPUT127), .ZN(new_n1211));
  NAND2_X1  g785(.A1(new_n1210), .A2(KEYINPUT127), .ZN(new_n1212));
  AOI21_X1  g786(.A(new_n1209), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g787(.A1(new_n936), .A2(new_n937), .ZN(new_n1214));
  AND3_X1   g788(.A1(new_n1213), .A2(new_n1026), .A3(new_n1214), .ZN(G308));
  NAND3_X1  g789(.A1(new_n1213), .A2(new_n1026), .A3(new_n1214), .ZN(G225));
endmodule


