//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT65), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  INV_X1    g0009(.A(G226), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  OAI22_X1  g0011(.A1(new_n202), .A2(new_n210), .B1(new_n205), .B2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G58), .B2(G232), .ZN(new_n213));
  INV_X1    g0013(.A(G97), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G107), .ZN(new_n216));
  INV_X1    g0016(.A(G264), .ZN(new_n217));
  OAI22_X1  g0017(.A1(new_n214), .A2(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(G87), .B2(G250), .ZN(new_n219));
  XOR2_X1   g0019(.A(KEYINPUT66), .B(G238), .Z(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G68), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n213), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G116), .ZN(new_n223));
  INV_X1    g0023(.A(G270), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT67), .Z(new_n228));
  NOR2_X1   g0028(.A1(new_n209), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT0), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  INV_X1    g0032(.A(G20), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  NOR3_X1   g0034(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(new_n226), .B2(KEYINPUT1), .ZN(new_n236));
  NAND3_X1  g0036(.A1(new_n228), .A2(new_n231), .A3(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(KEYINPUT68), .Z(G361));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G264), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n224), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n241), .B(KEYINPUT69), .Z(new_n242));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  INV_X1    g0043(.A(G232), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT2), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n210), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n242), .B(new_n247), .ZN(G358));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(new_n205), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G97), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(new_n216), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(new_n223), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n251), .B(new_n254), .Z(G351));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G150), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n233), .A2(G33), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT8), .B(G58), .ZN(new_n259));
  OAI221_X1 g0059(.A(new_n257), .B1(new_n258), .B2(new_n259), .C1(new_n204), .C2(new_n233), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n234), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n233), .A2(G1), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G13), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n260), .A2(new_n262), .B1(new_n202), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n262), .A2(new_n263), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G50), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n266), .A2(KEYINPUT9), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(KEYINPUT9), .B1(new_n266), .B2(new_n268), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n234), .B1(G33), .B2(G41), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT70), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G41), .A2(G45), .ZN(new_n278));
  OAI21_X1  g0078(.A(KEYINPUT70), .B1(new_n278), .B2(G1), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n272), .A2(new_n277), .A3(G274), .A4(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NOR2_X1   g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT71), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT71), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT3), .ZN(new_n286));
  INV_X1    g0086(.A(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n285), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(G1698), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT73), .ZN(new_n292));
  OAI21_X1  g0092(.A(KEYINPUT71), .B1(new_n282), .B2(new_n283), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n288), .A2(new_n285), .A3(new_n289), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT73), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(new_n296), .A3(G1698), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n292), .A2(G223), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n295), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G77), .ZN(new_n300));
  INV_X1    g0100(.A(G1698), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT72), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT72), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G1698), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n295), .A2(G222), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n298), .A2(new_n300), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n281), .B1(new_n307), .B2(new_n271), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n271), .A2(new_n275), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(new_n210), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n270), .B1(new_n313), .B2(G200), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT76), .ZN(new_n315));
  AOI211_X1 g0115(.A(new_n281), .B(new_n311), .C1(new_n307), .C2(new_n271), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(G190), .ZN(new_n317));
  AND4_X1   g0117(.A1(new_n315), .A2(new_n308), .A3(G190), .A4(new_n312), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n269), .B(new_n314), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT10), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G190), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT76), .B1(new_n313), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n316), .A2(new_n315), .A3(G190), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n325), .A2(KEYINPUT10), .A3(new_n269), .A4(new_n314), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT13), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT77), .B1(new_n291), .B2(new_n244), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n295), .A2(G226), .A3(new_n305), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT77), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n295), .A2(new_n330), .A3(G232), .A4(G1698), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n287), .A2(new_n214), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n328), .A2(new_n329), .A3(new_n331), .A4(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n271), .ZN(new_n335));
  INV_X1    g0135(.A(G238), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n280), .B1(new_n310), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n327), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  AOI211_X1 g0140(.A(KEYINPUT13), .B(new_n337), .C1(new_n334), .C2(new_n271), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(new_n342), .A3(G190), .ZN(new_n343));
  OAI21_X1  g0143(.A(G200), .B1(new_n339), .B2(new_n341), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n256), .A2(G50), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT78), .ZN(new_n346));
  INV_X1    g0146(.A(G68), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n345), .A2(new_n346), .B1(G20), .B2(new_n347), .ZN(new_n348));
  OAI221_X1 g0148(.A(new_n348), .B1(new_n346), .B2(new_n345), .C1(new_n205), .C2(new_n258), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n349), .A2(KEYINPUT11), .A3(new_n262), .ZN(new_n350));
  INV_X1    g0150(.A(new_n267), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n350), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n264), .A2(G68), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n353), .B(KEYINPUT12), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT11), .B1(new_n349), .B2(new_n262), .ZN(new_n355));
  NOR3_X1   g0155(.A1(new_n352), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n343), .A2(new_n344), .A3(new_n356), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT74), .B(G179), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n316), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n266), .A2(new_n268), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n360), .B(new_n361), .C1(G169), .C2(new_n316), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n321), .A2(new_n326), .A3(new_n357), .A4(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(G169), .B1(new_n339), .B2(new_n341), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT14), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n340), .A2(new_n342), .A3(G179), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT14), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n367), .B(G169), .C1(new_n339), .C2(new_n341), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n365), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n356), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n259), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n372), .A2(new_n256), .B1(G20), .B2(G77), .ZN(new_n373));
  XNOR2_X1  g0173(.A(KEYINPUT15), .B(G87), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n373), .B1(new_n258), .B2(new_n374), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n375), .A2(new_n262), .B1(G77), .B2(new_n267), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n264), .A2(G77), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n377), .B(KEYINPUT75), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n292), .A2(new_n220), .A3(new_n297), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n295), .A2(G232), .A3(new_n305), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n380), .B(new_n381), .C1(new_n216), .C2(new_n295), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n281), .B1(new_n382), .B2(new_n271), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n310), .A2(new_n211), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n379), .B1(new_n386), .B2(new_n358), .ZN(new_n387));
  AOI21_X1  g0187(.A(G169), .B1(new_n383), .B2(new_n385), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n386), .A2(G200), .ZN(new_n391));
  INV_X1    g0191(.A(new_n379), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n383), .A2(G190), .A3(new_n385), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n371), .A2(new_n390), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT16), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n293), .A2(new_n294), .A3(new_n233), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT7), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n288), .A2(KEYINPUT7), .A3(new_n233), .A4(new_n289), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT79), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n282), .A2(new_n283), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT79), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n402), .A2(new_n403), .A3(KEYINPUT7), .A4(new_n233), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n347), .B1(new_n399), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(G58), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n407), .A2(new_n347), .ZN(new_n408));
  OAI21_X1  g0208(.A(G20), .B1(new_n408), .B2(new_n201), .ZN(new_n409));
  INV_X1    g0209(.A(G159), .ZN(new_n410));
  INV_X1    g0210(.A(new_n256), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n396), .B1(new_n406), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT80), .ZN(new_n414));
  INV_X1    g0214(.A(new_n262), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n288), .A2(new_n289), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n398), .B1(new_n416), .B2(G20), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n400), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n412), .B1(new_n418), .B2(G68), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n415), .B1(new_n419), .B2(KEYINPUT16), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT80), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n421), .B(new_n396), .C1(new_n406), .C2(new_n412), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n414), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n372), .B(KEYINPUT81), .C1(G1), .C2(new_n233), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT81), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n259), .B2(new_n263), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n424), .A2(new_n264), .A3(new_n415), .A4(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n264), .B2(new_n372), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n428), .B(KEYINPUT82), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(G223), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n302), .B2(new_n304), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n210), .A2(new_n301), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n416), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G87), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n272), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(new_n281), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n309), .A2(G232), .ZN(new_n438));
  AOI21_X1  g0238(.A(G169), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n438), .ZN(new_n440));
  NOR4_X1   g0240(.A1(new_n436), .A2(new_n281), .A3(new_n440), .A4(new_n358), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT83), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  XNOR2_X1  g0242(.A(KEYINPUT72), .B(G1698), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n443), .A2(new_n431), .B1(new_n210), .B2(new_n301), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n444), .A2(new_n416), .B1(G33), .B2(G87), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n280), .B(new_n438), .C1(new_n445), .C2(new_n272), .ZN(new_n446));
  INV_X1    g0246(.A(G169), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT83), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n448), .B(new_n449), .C1(new_n358), .C2(new_n446), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n442), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n430), .A2(KEYINPUT18), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT84), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT84), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n430), .A2(new_n451), .A3(new_n454), .A4(KEYINPUT18), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n430), .A2(new_n451), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT18), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n453), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n446), .A2(G200), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n437), .A2(G190), .A3(new_n438), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n423), .A2(new_n429), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  XNOR2_X1  g0262(.A(new_n462), .B(KEYINPUT17), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n363), .A2(new_n395), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G283), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n416), .A2(new_n305), .A3(G244), .ZN(new_n468));
  XOR2_X1   g0268(.A(KEYINPUT85), .B(KEYINPUT4), .Z(new_n469));
  AOI21_X1  g0269(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g0270(.A1(KEYINPUT4), .A2(G244), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n295), .A2(new_n305), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n295), .A2(G250), .A3(G1698), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n470), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n271), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT5), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT86), .B1(new_n476), .B2(G41), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT86), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n478), .A2(new_n273), .A3(KEYINPUT5), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n274), .A2(G1), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n476), .A2(G41), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n477), .A2(new_n479), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n482), .A2(G257), .A3(new_n272), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G274), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n482), .A2(new_n485), .A3(new_n271), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n475), .A2(G190), .A3(new_n484), .A4(new_n487), .ZN(new_n488));
  AOI211_X1 g0288(.A(new_n483), .B(new_n486), .C1(new_n474), .C2(new_n271), .ZN(new_n489));
  INV_X1    g0289(.A(G200), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n265), .A2(new_n214), .ZN(new_n492));
  INV_X1    g0292(.A(G1), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G33), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n415), .A2(new_n264), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G97), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n216), .B1(new_n399), .B2(new_n405), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n411), .A2(new_n205), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT6), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n214), .A2(new_n216), .ZN(new_n501));
  NOR2_X1   g0301(.A1(G97), .A2(G107), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n216), .A2(KEYINPUT6), .A3(G97), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(new_n233), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n498), .A2(new_n499), .A3(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n492), .B(new_n497), .C1(new_n507), .C2(new_n415), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n491), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n475), .A2(new_n358), .A3(new_n484), .A4(new_n487), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n489), .B2(new_n447), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n508), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT87), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT87), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n511), .A2(new_n514), .A3(new_n508), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n509), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n482), .A2(new_n272), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G264), .ZN(new_n518));
  INV_X1    g0318(.A(G250), .ZN(new_n519));
  OAI22_X1  g0319(.A1(new_n443), .A2(new_n519), .B1(new_n215), .B2(new_n301), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n520), .A2(new_n416), .B1(G33), .B2(G294), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n518), .B(new_n487), .C1(new_n272), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G169), .ZN(new_n523));
  INV_X1    g0323(.A(G179), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(new_n522), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT89), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT23), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT23), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT89), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n527), .A2(new_n529), .A3(G20), .A4(new_n216), .ZN(new_n530));
  OAI211_X1 g0330(.A(KEYINPUT89), .B(new_n528), .C1(new_n233), .C2(G107), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(KEYINPUT22), .A2(G87), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n416), .A2(new_n534), .B1(G33), .B2(G116), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n532), .B1(new_n535), .B2(G20), .ZN(new_n536));
  INV_X1    g0336(.A(G87), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(G20), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT22), .B1(new_n295), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(KEYINPUT90), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n538), .B1(new_n284), .B2(new_n290), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT22), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(G33), .A2(G116), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n402), .B2(new_n533), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n545), .A2(new_n233), .B1(new_n530), .B2(new_n531), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT90), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n543), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n540), .A2(new_n548), .A3(KEYINPUT24), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT24), .ZN(new_n550));
  OAI211_X1 g0350(.A(KEYINPUT90), .B(new_n550), .C1(new_n536), .C2(new_n539), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n262), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n265), .A2(KEYINPUT25), .A3(new_n216), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT25), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n264), .B2(G107), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n496), .A2(G107), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n552), .A2(KEYINPUT91), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT91), .B1(new_n552), .B2(new_n556), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n525), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT19), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n258), .B2(new_n214), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n416), .A2(new_n233), .A3(G68), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n537), .A2(new_n214), .A3(new_n216), .ZN(new_n563));
  XNOR2_X1  g0363(.A(new_n563), .B(KEYINPUT88), .ZN(new_n564));
  AOI21_X1  g0364(.A(G20), .B1(new_n332), .B2(KEYINPUT19), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n561), .B(new_n562), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n262), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n265), .A2(new_n374), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  OR3_X1    g0370(.A1(new_n271), .A2(new_n519), .A3(new_n480), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n305), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n544), .B1(new_n573), .B2(new_n402), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n572), .B1(new_n574), .B2(new_n271), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n480), .A2(G274), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(G190), .A3(new_n576), .ZN(new_n577));
  OAI22_X1  g0377(.A1(new_n443), .A2(new_n336), .B1(new_n211), .B2(new_n301), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n578), .A2(new_n416), .B1(G33), .B2(G116), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n576), .B(new_n571), .C1(new_n579), .C2(new_n272), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G200), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n496), .A2(G87), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n570), .A2(new_n577), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n495), .A2(new_n374), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n569), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n575), .A2(new_n359), .A3(new_n576), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n580), .A2(new_n447), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n583), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n215), .B1(new_n302), .B2(new_n304), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n217), .A2(new_n301), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n416), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n293), .A2(new_n294), .A3(G303), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n486), .B1(new_n594), .B2(new_n271), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n482), .A2(G270), .A3(new_n272), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(G190), .A3(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n264), .A2(G116), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n415), .A2(new_n264), .A3(G116), .A4(new_n494), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n261), .A2(new_n234), .B1(G20), .B2(new_n223), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n466), .B(new_n233), .C1(G33), .C2(new_n214), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(KEYINPUT20), .A3(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT20), .B1(new_n602), .B2(new_n603), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n600), .B(new_n601), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n272), .B1(new_n592), .B2(new_n593), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n609), .A2(new_n486), .A3(new_n596), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n598), .B(new_n608), .C1(new_n490), .C2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(G179), .A3(new_n607), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT21), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n607), .A2(G169), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n613), .B1(new_n610), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n594), .A2(new_n271), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n616), .A2(new_n487), .A3(new_n597), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n223), .A2(G20), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n603), .A2(new_n262), .A3(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT20), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n599), .B1(new_n621), .B2(new_n604), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n447), .B1(new_n622), .B2(new_n601), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n617), .A2(new_n623), .A3(KEYINPUT21), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n611), .A2(new_n612), .A3(new_n615), .A4(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n589), .A2(new_n625), .ZN(new_n626));
  OR2_X1    g0426(.A1(new_n521), .A2(new_n272), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n627), .A2(new_n322), .A3(new_n487), .A4(new_n518), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n522), .A2(new_n490), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(new_n629), .A3(KEYINPUT92), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT92), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n522), .A2(new_n631), .A3(new_n490), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n630), .A2(new_n552), .A3(new_n556), .A4(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n559), .A2(new_n626), .A3(new_n633), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n465), .A2(new_n516), .A3(new_n634), .ZN(G372));
  AND3_X1   g0435(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT93), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT93), .B1(new_n586), .B2(new_n587), .ZN(new_n637));
  OAI22_X1  g0437(.A1(new_n636), .A2(new_n637), .B1(new_n584), .B2(new_n569), .ZN(new_n638));
  INV_X1    g0438(.A(new_n512), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n639), .A2(new_n638), .A3(new_n640), .A4(new_n583), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n511), .A2(new_n514), .A3(new_n508), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n514), .B1(new_n511), .B2(new_n508), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n642), .A2(new_n643), .A3(new_n589), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n638), .B(new_n641), .C1(new_n644), .C2(new_n640), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n638), .A2(new_n633), .A3(new_n583), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n552), .A2(new_n556), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n525), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n615), .A2(new_n624), .A3(new_n612), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(KEYINPUT94), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT94), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n648), .A2(new_n652), .A3(new_n649), .ZN(new_n653));
  AND4_X1   g0453(.A1(new_n516), .A2(new_n646), .A3(new_n651), .A4(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n465), .B1(new_n645), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n362), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n458), .A2(new_n452), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n389), .B1(new_n369), .B2(new_n370), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n463), .A2(new_n357), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n321), .A2(new_n326), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n656), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n655), .A2(new_n662), .ZN(G369));
  INV_X1    g0463(.A(new_n633), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT91), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n647), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n552), .A2(KEYINPUT91), .A3(new_n556), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n664), .B1(new_n668), .B2(new_n525), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT97), .ZN(new_n670));
  INV_X1    g0470(.A(G13), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G20), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT27), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(new_n673), .A3(new_n493), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n493), .A2(new_n233), .A3(G13), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n674), .A2(new_n676), .A3(G213), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT95), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g0479(.A(KEYINPUT96), .B(G343), .Z(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n670), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n677), .B(KEYINPUT95), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n683), .A2(KEYINPUT97), .A3(new_n680), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n668), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n669), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n559), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n685), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT100), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT99), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n615), .A2(new_n624), .A3(new_n612), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n608), .B1(new_n682), .B2(new_n684), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT98), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n695), .B(new_n696), .C1(new_n625), .C2(new_n694), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n694), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n649), .A2(new_n611), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n696), .B1(new_n700), .B2(new_n695), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n692), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n490), .B1(new_n595), .B2(new_n597), .ZN(new_n703));
  NOR4_X1   g0503(.A1(new_n609), .A2(new_n596), .A3(new_n486), .A4(new_n322), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n703), .A2(new_n704), .A3(new_n607), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n693), .A2(new_n705), .A3(new_n694), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n693), .A2(new_n694), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT98), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n708), .A2(KEYINPUT99), .A3(new_n697), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n702), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n691), .B1(new_n710), .B2(G330), .ZN(new_n711));
  INV_X1    g0511(.A(G330), .ZN(new_n712));
  AOI211_X1 g0512(.A(KEYINPUT100), .B(new_n712), .C1(new_n702), .C2(new_n709), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n690), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n649), .A2(new_n685), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n559), .A2(new_n633), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n685), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n647), .A2(new_n525), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT101), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n716), .A2(KEYINPUT101), .A3(new_n718), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n714), .A2(new_n723), .ZN(G399));
  NAND2_X1  g0524(.A1(new_n564), .A2(new_n223), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n229), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G41), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n726), .A2(G1), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n232), .B2(new_n729), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT28), .ZN(new_n732));
  INV_X1    g0532(.A(new_n638), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n733), .B1(new_n644), .B2(new_n640), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n559), .A2(new_n649), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(new_n516), .A3(new_n646), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n638), .A2(new_n583), .ZN(new_n737));
  OAI21_X1  g0537(.A(KEYINPUT26), .B1(new_n737), .B2(new_n512), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n734), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n717), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT29), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT29), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n742), .B(new_n717), .C1(new_n654), .C2(new_n645), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n617), .A2(new_n524), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n518), .B1(new_n521), .B2(new_n272), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n580), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n744), .A2(new_n489), .A3(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT30), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n617), .A2(new_n522), .A3(new_n359), .A4(new_n580), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n750), .A2(new_n489), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n747), .A2(new_n748), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n749), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n685), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT31), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n753), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n669), .A2(new_n516), .A3(new_n626), .A4(new_n717), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT102), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n634), .A2(KEYINPUT102), .A3(new_n516), .A4(new_n717), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n758), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n741), .B(new_n743), .C1(new_n712), .C2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n732), .B1(new_n765), .B2(G1), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT103), .Z(G364));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n708), .A2(new_n697), .A3(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n233), .A2(G190), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n490), .A2(G179), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G283), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G179), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G329), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n774), .A2(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G294), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n776), .A2(G190), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n299), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n233), .A2(new_n322), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(new_n773), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n779), .B(new_n784), .C1(G303), .C2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n358), .A2(new_n490), .A3(new_n772), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G311), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n358), .A2(G20), .A3(G200), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n322), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n358), .A2(new_n490), .A3(new_n785), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n793), .A2(G326), .B1(new_n795), .B2(G322), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n792), .A2(G190), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT33), .B(G317), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n788), .A2(new_n791), .A3(new_n796), .A4(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n777), .ZN(new_n801));
  XOR2_X1   g0601(.A(KEYINPUT104), .B(G159), .Z(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT32), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n774), .A2(new_n216), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n783), .A2(new_n214), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n797), .A2(G68), .B1(new_n790), .B2(G77), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n793), .A2(G50), .B1(G87), .B2(new_n787), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n807), .A2(new_n808), .A3(new_n809), .A4(new_n295), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n794), .A2(new_n407), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n800), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n234), .B1(G20), .B2(new_n447), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n727), .A2(new_n416), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n232), .A2(G45), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(new_n251), .C2(new_n274), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n295), .A2(G355), .A3(new_n229), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n816), .B(new_n817), .C1(G116), .C2(new_n229), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n770), .A2(new_n813), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n812), .A2(new_n813), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n493), .B1(new_n672), .B2(G45), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n728), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n771), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n711), .A2(new_n713), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n823), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n710), .B2(G330), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n824), .B1(new_n826), .B2(new_n828), .ZN(G396));
  OAI21_X1  g0629(.A(new_n717), .B1(new_n654), .B2(new_n645), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n387), .A2(new_n388), .A3(new_n685), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n685), .A2(new_n379), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT105), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n394), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n831), .B1(new_n390), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n830), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n836), .B(new_n717), .C1(new_n654), .C2(new_n645), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n712), .B2(new_n763), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n761), .A2(new_n762), .ZN(new_n842));
  INV_X1    g0642(.A(new_n758), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n844), .A2(new_n838), .A3(G330), .A4(new_n839), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n823), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n793), .A2(G303), .B1(new_n795), .B2(G294), .ZN(new_n847));
  INV_X1    g0647(.A(new_n797), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n847), .B1(new_n775), .B2(new_n848), .ZN(new_n849));
  AOI22_X1  g0649(.A1(G107), .A2(new_n787), .B1(new_n801), .B2(G311), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n850), .B(new_n299), .C1(new_n214), .C2(new_n783), .ZN(new_n851));
  INV_X1    g0651(.A(new_n774), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n851), .B1(G87), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n849), .B(new_n854), .C1(G116), .C2(new_n790), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n793), .A2(G137), .B1(new_n790), .B2(new_n802), .ZN(new_n857));
  INV_X1    g0657(.A(G143), .ZN(new_n858));
  INV_X1    g0658(.A(G150), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n857), .B1(new_n858), .B2(new_n794), .C1(new_n859), .C2(new_n848), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT34), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n852), .A2(G68), .ZN(new_n862));
  INV_X1    g0662(.A(G132), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n416), .B1(new_n777), .B2(new_n863), .C1(new_n202), .C2(new_n786), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(G58), .B2(new_n782), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n861), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n856), .A2(new_n866), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n837), .A2(new_n768), .B1(new_n813), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n813), .A2(new_n768), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n205), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n827), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n846), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT106), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR3_X1   g0674(.A1(new_n846), .A2(KEYINPUT106), .A3(new_n871), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n874), .A2(new_n875), .ZN(G384));
  OAI21_X1  g0676(.A(new_n420), .B1(KEYINPUT16), .B2(new_n419), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n429), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n683), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n464), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n430), .A2(new_n683), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n456), .A2(new_n882), .A3(new_n883), .A4(new_n462), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n878), .B1(new_n451), .B2(new_n683), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n885), .A2(new_n462), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n884), .B1(new_n886), .B2(new_n883), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n881), .A2(KEYINPUT38), .A3(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT38), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n879), .B1(new_n459), .B2(new_n463), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n883), .B1(new_n885), .B2(new_n462), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n456), .A2(new_n882), .A3(new_n462), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n891), .B1(new_n893), .B2(new_n883), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n889), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n888), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n356), .A2(new_n717), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n371), .A2(new_n357), .A3(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n357), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n370), .B(new_n685), .C1(new_n900), .C2(new_n369), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n902), .A2(new_n837), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n755), .A2(KEYINPUT108), .ZN(new_n904));
  OR2_X1    g0704(.A1(new_n754), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n754), .A2(new_n904), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n842), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n896), .A2(new_n903), .A3(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT40), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n462), .A2(KEYINPUT17), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n462), .A2(KEYINPUT17), .ZN(new_n913));
  INV_X1    g0713(.A(new_n452), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT18), .B1(new_n430), .B2(new_n451), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n912), .A2(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n882), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n892), .A2(KEYINPUT37), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n884), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n888), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n923), .A2(new_n903), .A3(KEYINPUT40), .A4(new_n908), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n911), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n908), .A2(new_n465), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n925), .B(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n927), .A2(new_n712), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n369), .A2(new_n370), .A3(new_n717), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n890), .A2(new_n894), .A3(new_n889), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n931), .A2(new_n921), .A3(KEYINPUT39), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT39), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n888), .B2(new_n895), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n930), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n657), .A2(new_n683), .ZN(new_n936));
  INV_X1    g0736(.A(new_n831), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n902), .B1(new_n937), .B2(new_n839), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n936), .B1(new_n938), .B2(new_n896), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n743), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n742), .B1(new_n739), .B2(new_n717), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n465), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n662), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n940), .B(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n928), .B(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n493), .B2(new_n672), .ZN(new_n947));
  OAI21_X1  g0747(.A(G77), .B1(new_n407), .B2(new_n347), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n948), .A2(new_n232), .B1(G50), .B2(new_n347), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(G1), .A3(new_n671), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT35), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n233), .B(new_n234), .C1(new_n505), .C2(new_n951), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n952), .B(G116), .C1(new_n951), .C2(new_n505), .ZN(new_n953));
  XOR2_X1   g0753(.A(KEYINPUT107), .B(KEYINPUT36), .Z(new_n954));
  XNOR2_X1  g0754(.A(new_n953), .B(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n947), .A2(new_n950), .A3(new_n955), .ZN(G367));
  AOI22_X1  g0756(.A1(new_n797), .A2(new_n802), .B1(new_n790), .B2(G50), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n859), .B2(new_n794), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n783), .A2(new_n347), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(new_n299), .ZN(new_n960));
  AOI22_X1  g0760(.A1(G58), .A2(new_n787), .B1(new_n852), .B2(G77), .ZN(new_n961));
  INV_X1    g0761(.A(G137), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n960), .B(new_n961), .C1(new_n962), .C2(new_n777), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n958), .B(new_n963), .C1(G143), .C2(new_n793), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT114), .Z(new_n965));
  NOR2_X1   g0765(.A1(new_n786), .A2(new_n223), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT46), .ZN(new_n967));
  INV_X1    g0767(.A(new_n793), .ZN(new_n968));
  INV_X1    g0768(.A(G311), .ZN(new_n969));
  INV_X1    g0769(.A(G317), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n968), .A2(new_n969), .B1(new_n970), .B2(new_n777), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n967), .B(new_n971), .C1(G107), .C2(new_n782), .ZN(new_n972));
  INV_X1    g0772(.A(G303), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n775), .A2(new_n789), .B1(new_n794), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(new_n797), .B2(G294), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n972), .B(new_n975), .C1(new_n214), .C2(new_n774), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n965), .B1(new_n416), .B2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(KEYINPUT115), .B(KEYINPUT47), .Z(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n827), .B1(new_n979), .B2(new_n813), .ZN(new_n980));
  INV_X1    g0780(.A(new_n814), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n819), .B1(new_n229), .B2(new_n374), .C1(new_n241), .C2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n717), .B1(new_n570), .B2(new_n582), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n638), .A2(new_n983), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n638), .A2(new_n583), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n984), .B1(new_n985), .B2(new_n983), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT109), .Z(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n770), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n980), .A2(new_n982), .A3(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT45), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT111), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n508), .A2(new_n685), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n516), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n639), .A2(new_n685), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n991), .B1(new_n723), .B2(new_n995), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n716), .A2(KEYINPUT101), .A3(new_n718), .ZN(new_n997));
  AOI21_X1  g0797(.A(KEYINPUT101), .B1(new_n716), .B2(new_n718), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n991), .B(new_n995), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n990), .B1(new_n996), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(KEYINPUT111), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1003), .A2(KEYINPUT45), .A3(new_n999), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT44), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n723), .B2(new_n995), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n995), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1007), .A2(new_n721), .A3(KEYINPUT44), .A4(new_n722), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1001), .A2(new_n1004), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n714), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n716), .B1(new_n690), .B2(new_n715), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n825), .B2(KEYINPUT112), .ZN(new_n1014));
  AND3_X1   g0814(.A1(new_n708), .A2(KEYINPUT99), .A3(new_n697), .ZN(new_n1015));
  AOI21_X1  g0815(.A(KEYINPUT99), .B1(new_n708), .B2(new_n697), .ZN(new_n1016));
  OAI21_X1  g0816(.A(G330), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(KEYINPUT100), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n710), .A2(new_n691), .A3(G330), .ZN(new_n1019));
  AND4_X1   g0819(.A1(KEYINPUT112), .A2(new_n1018), .A3(new_n1019), .A4(new_n1013), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n1014), .A2(new_n764), .A3(new_n1020), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1001), .A2(new_n714), .A3(new_n1004), .A4(new_n1009), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1012), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n765), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n728), .B(KEYINPUT41), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(KEYINPUT113), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT113), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1024), .A2(new_n1028), .A3(new_n1025), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n822), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT110), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n987), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT43), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n987), .A2(new_n1031), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n993), .A2(new_n716), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT42), .Z(new_n1037));
  NAND2_X1  g0837(.A1(new_n995), .A2(new_n688), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n513), .A2(new_n515), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n685), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1035), .B(new_n1041), .C1(new_n1033), .C2(new_n987), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n1041), .B2(new_n1035), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1011), .A2(new_n995), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1043), .B(new_n1044), .Z(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n989), .B1(new_n1030), .B2(new_n1046), .ZN(G387));
  INV_X1    g0847(.A(new_n1021), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n764), .B1(new_n1014), .B2(new_n1020), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n728), .B(KEYINPUT118), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1048), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  OR3_X1    g0852(.A1(new_n1014), .A2(new_n821), .A3(new_n1020), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n783), .A2(new_n374), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n402), .B1(new_n852), .B2(G97), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n787), .A2(G77), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n801), .A2(G150), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n797), .A2(new_n372), .B1(new_n790), .B2(G68), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n202), .B2(new_n794), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1058), .B(new_n1060), .C1(G159), .C2(new_n793), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT116), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n793), .A2(G322), .B1(new_n790), .B2(G303), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n970), .B2(new_n794), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G311), .B2(new_n797), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT48), .Z(new_n1066));
  AOI22_X1  g0866(.A1(new_n787), .A2(G294), .B1(new_n782), .B2(G283), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT117), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1069), .A2(KEYINPUT49), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(KEYINPUT49), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n416), .B1(new_n801), .B2(G326), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n774), .A2(new_n223), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1062), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n827), .B1(new_n1075), .B2(new_n813), .ZN(new_n1076));
  OAI21_X1  g0876(.A(KEYINPUT50), .B1(new_n259), .B2(G50), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n259), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1078), .A2(G45), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n726), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(G68), .B2(G77), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n814), .B1(new_n247), .B2(new_n274), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n725), .A2(new_n229), .A3(new_n295), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n229), .A2(G107), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n819), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n770), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1076), .B(new_n1086), .C1(new_n690), .C2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1052), .A2(new_n1053), .A3(new_n1088), .ZN(G393));
  NAND3_X1  g0889(.A1(new_n1012), .A2(new_n822), .A3(new_n1022), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n995), .A2(new_n1087), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n1091), .A2(KEYINPUT119), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n254), .A2(new_n814), .B1(G97), .B2(new_n727), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n819), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1091), .A2(KEYINPUT119), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n416), .B1(new_n777), .B2(new_n858), .C1(new_n537), .C2(new_n774), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n848), .A2(new_n202), .B1(new_n259), .B2(new_n789), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1096), .B(new_n1097), .C1(G77), .C2(new_n782), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n793), .A2(G150), .B1(new_n795), .B2(G159), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(KEYINPUT120), .B(KEYINPUT51), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1099), .B(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1098), .B(new_n1101), .C1(new_n347), .C2(new_n786), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT121), .Z(new_n1103));
  AOI22_X1  g0903(.A1(new_n793), .A2(G317), .B1(new_n795), .B2(G311), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT52), .Z(new_n1105));
  AOI21_X1  g0905(.A(new_n295), .B1(G322), .B2(new_n801), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n805), .B1(G283), .B2(new_n787), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n797), .A2(G303), .B1(new_n790), .B2(G294), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n223), .B2(new_n783), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT122), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1103), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n827), .B1(new_n1112), .B2(new_n813), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1092), .A2(new_n1094), .A3(new_n1095), .A4(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1090), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT123), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1090), .A2(KEYINPUT123), .A3(new_n1114), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1023), .A2(new_n1051), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1012), .A2(new_n1022), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n1048), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1117), .A2(new_n1118), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(G390));
  NAND3_X1  g0923(.A1(new_n908), .A2(G330), .A3(new_n465), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n943), .A2(new_n1124), .A3(new_n662), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n899), .A2(new_n901), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n836), .A2(G330), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n908), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n902), .B1(new_n763), .B2(new_n1127), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n839), .A2(new_n937), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n844), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n761), .A2(new_n762), .B1(new_n905), .B2(new_n906), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n902), .B1(new_n1135), .B2(new_n1127), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n390), .A2(new_n835), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n739), .A2(new_n717), .A3(new_n1137), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n1138), .A2(new_n937), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1134), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1125), .B1(new_n1133), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(KEYINPUT38), .B1(new_n881), .B2(new_n887), .ZN(new_n1142));
  OAI21_X1  g0942(.A(KEYINPUT39), .B1(new_n1142), .B2(new_n931), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n922), .A2(new_n888), .A3(new_n933), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(new_n930), .C2(new_n938), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n929), .B1(new_n931), .B2(new_n921), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n902), .B1(new_n1138), .B2(new_n937), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1134), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1145), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1129), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1141), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n930), .B1(new_n1132), .B2(new_n1126), .ZN(new_n1154));
  NOR3_X1   g0954(.A1(new_n1154), .A2(new_n932), .A3(new_n934), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1129), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n943), .A2(new_n1124), .A3(new_n662), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1134), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1129), .A2(new_n1130), .B1(new_n937), .B2(new_n839), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1145), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1157), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1153), .A2(new_n1051), .A3(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1143), .A2(new_n768), .A3(new_n1144), .ZN(new_n1165));
  INV_X1    g0965(.A(G125), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n295), .B1(new_n1166), .B2(new_n777), .ZN(new_n1167));
  OR3_X1    g0967(.A1(new_n786), .A2(KEYINPUT53), .A3(new_n859), .ZN(new_n1168));
  OAI21_X1  g0968(.A(KEYINPUT53), .B1(new_n786), .B2(new_n859), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1168), .B(new_n1169), .C1(new_n410), .C2(new_n783), .ZN(new_n1170));
  XOR2_X1   g0970(.A(KEYINPUT54), .B(G143), .Z(new_n1171));
  AOI211_X1 g0971(.A(new_n1167), .B(new_n1170), .C1(new_n790), .C2(new_n1171), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n848), .A2(new_n962), .B1(new_n863), .B2(new_n794), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G128), .B2(new_n793), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1172), .B(new_n1174), .C1(new_n202), .C2(new_n774), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n789), .A2(new_n214), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n862), .B1(new_n537), .B2(new_n786), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n299), .B1(new_n205), .B2(new_n783), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(G294), .C2(new_n801), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n797), .A2(G107), .B1(new_n795), .B2(G116), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(new_n775), .C2(new_n968), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1175), .B1(new_n1176), .B2(new_n1181), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT124), .Z(new_n1183));
  AOI21_X1  g0983(.A(new_n827), .B1(new_n1183), .B2(new_n813), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1165), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n259), .B2(new_n869), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1157), .A2(new_n1162), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1186), .B1(new_n1187), .B2(new_n822), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1164), .A2(new_n1188), .ZN(G378));
  INV_X1    g0989(.A(KEYINPUT57), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n911), .A2(G330), .A3(new_n924), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT125), .B(KEYINPUT56), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n321), .A2(new_n326), .A3(new_n362), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(KEYINPUT55), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT55), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n321), .A2(new_n326), .A3(new_n1196), .A4(new_n362), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n361), .A2(new_n683), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1198), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1193), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1198), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(new_n1192), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1201), .A2(new_n1206), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1207), .A2(new_n935), .A3(new_n939), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1207), .B1(new_n935), .B2(new_n939), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1191), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1207), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n940), .A2(new_n1211), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n911), .A2(G330), .A3(new_n924), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1207), .A2(new_n935), .A3(new_n939), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1210), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1125), .B1(new_n1187), .B2(new_n1141), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1190), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1153), .A2(new_n1158), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1219), .A2(KEYINPUT57), .A3(new_n1215), .A4(new_n1210), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1218), .A2(new_n1220), .A3(new_n1051), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1210), .A2(new_n822), .A3(new_n1215), .ZN(new_n1222));
  INV_X1    g1022(.A(G128), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n848), .A2(new_n863), .B1(new_n1223), .B2(new_n794), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n787), .A2(new_n1171), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n859), .B2(new_n783), .C1(new_n968), .C2(new_n1166), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1224), .B(new_n1226), .C1(G137), .C2(new_n790), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT59), .ZN(new_n1228));
  AOI21_X1  g1028(.A(G41), .B1(new_n801), .B2(G124), .ZN(new_n1229));
  AOI21_X1  g1029(.A(G33), .B1(new_n852), .B2(new_n802), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n202), .B1(new_n282), .B2(G41), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n848), .A2(new_n214), .B1(new_n216), .B2(new_n794), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(G116), .B2(new_n793), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1056), .B1(new_n407), .B2(new_n774), .C1(new_n775), .C2(new_n777), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(new_n1235), .A2(G41), .A3(new_n416), .A4(new_n959), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1234), .B(new_n1236), .C1(new_n374), .C2(new_n789), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(KEYINPUT58), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1231), .A2(new_n1232), .A3(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n827), .B1(new_n1239), .B2(new_n813), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n869), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1240), .B1(G50), .B2(new_n1241), .C1(new_n1211), .C2(new_n769), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1222), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1221), .A2(new_n1244), .ZN(G375));
  OAI21_X1  g1045(.A(new_n822), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n786), .A2(new_n214), .B1(new_n774), .B2(new_n205), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1054), .A2(new_n299), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1247), .B(new_n1248), .C1(G303), .C2(new_n801), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n797), .A2(G116), .B1(new_n790), .B2(G107), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n775), .B2(new_n794), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1249), .B(new_n1252), .C1(new_n780), .C2(new_n968), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1253), .B(KEYINPUT126), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n968), .A2(new_n863), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n797), .A2(new_n1171), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n787), .A2(G159), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n416), .B1(new_n777), .B2(new_n1223), .C1(new_n407), .C2(new_n774), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(G50), .B2(new_n782), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(G137), .A2(new_n795), .B1(new_n790), .B2(G150), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1256), .A2(new_n1257), .A3(new_n1259), .A4(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1254), .B1(new_n1255), .B2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n827), .B1(new_n1262), .B2(new_n813), .ZN(new_n1263));
  OAI221_X1 g1063(.A(new_n1263), .B1(G68), .B2(new_n1241), .C1(new_n1126), .C2(new_n769), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1246), .A2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1133), .A2(new_n1125), .A3(new_n1140), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1161), .A2(new_n1266), .A3(new_n1025), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(G381));
  NOR3_X1   g1068(.A1(G387), .A2(G390), .A3(G381), .ZN(new_n1269));
  AND4_X1   g1069(.A1(new_n1188), .A2(new_n1222), .A3(new_n1164), .A4(new_n1242), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1221), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1269), .A2(new_n1272), .A3(new_n1273), .ZN(G407));
  OAI211_X1 g1074(.A(G407), .B(G213), .C1(new_n680), .C2(new_n1271), .ZN(G409));
  AND2_X1   g1075(.A1(new_n681), .A2(G213), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1219), .A2(new_n1025), .A3(new_n1215), .A4(new_n1210), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1276), .B1(new_n1270), .B2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1161), .B1(new_n1157), .B2(new_n1162), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1215), .B(new_n1210), .C1(new_n1279), .C2(new_n1125), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1050), .B1(new_n1280), .B2(new_n1190), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1243), .B1(new_n1281), .B2(new_n1220), .ZN(new_n1282));
  INV_X1    g1082(.A(G378), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1278), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT60), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1050), .B1(new_n1266), .B2(new_n1285), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1133), .A2(new_n1125), .A3(KEYINPUT60), .A4(new_n1140), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1286), .A2(new_n1161), .A3(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(G384), .A2(new_n1288), .A3(new_n1265), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(G384), .B1(new_n1265), .B2(new_n1288), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(KEYINPUT62), .B1(new_n1284), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1276), .A2(G2897), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1288), .A2(new_n1265), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1298), .B1(new_n874), .B2(new_n875), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(new_n1289), .A3(new_n1295), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT61), .B1(new_n1284), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(G375), .A2(G378), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT62), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1303), .A2(new_n1304), .A3(new_n1278), .A4(new_n1292), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1294), .A2(new_n1302), .A3(new_n1305), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(G393), .B(G396), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(G387), .A2(new_n1122), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1028), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1025), .ZN(new_n1310));
  AOI211_X1 g1110(.A(KEYINPUT113), .B(new_n1310), .C1(new_n1023), .C2(new_n765), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n821), .B1(new_n1309), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1045), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1313), .A2(new_n989), .A3(G390), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1308), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT127), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1307), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(G390), .B1(new_n1313), .B2(new_n989), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n989), .ZN(new_n1319));
  AOI211_X1 g1119(.A(new_n1319), .B(new_n1122), .C1(new_n1312), .C2(new_n1045), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1316), .B(new_n1307), .C1(new_n1318), .C2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1317), .A2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1316), .B1(new_n1318), .B2(new_n1320), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1307), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1303), .A2(KEYINPUT63), .A3(new_n1278), .A4(new_n1292), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1326), .A2(new_n1321), .A3(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT61), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT63), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1330), .B1(new_n1284), .B2(new_n1301), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1284), .A2(new_n1293), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1329), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1333));
  OAI22_X1  g1133(.A1(new_n1306), .A2(new_n1323), .B1(new_n1328), .B2(new_n1333), .ZN(G405));
  NAND2_X1  g1134(.A1(new_n1303), .A2(new_n1271), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(new_n1292), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1303), .A2(new_n1271), .A3(new_n1293), .ZN(new_n1337));
  AND4_X1   g1137(.A1(new_n1326), .A2(new_n1336), .A3(new_n1321), .A4(new_n1337), .ZN(new_n1338));
  AOI22_X1  g1138(.A1(new_n1326), .A2(new_n1321), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1338), .A2(new_n1339), .ZN(G402));
endmodule


