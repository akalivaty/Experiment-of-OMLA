//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n555, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1140, new_n1141, new_n1142,
    new_n1143;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT67), .Z(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n461), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n469), .A2(new_n464), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n472), .B1(new_n463), .B2(G2104), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n470), .A2(G137), .A3(new_n471), .A4(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n461), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n468), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT71), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n473), .A2(new_n469), .A3(G2105), .A4(new_n464), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT70), .Z(new_n485));
  NAND3_X1  g060(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI211_X1 g062(.A(new_n481), .B(new_n485), .C1(G136), .C2(new_n487), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n473), .A2(new_n469), .A3(new_n490), .A4(new_n464), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n462), .A2(new_n464), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n489), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n491), .A2(KEYINPUT4), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G114), .C2(new_n471), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n482), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n494), .A2(new_n498), .ZN(G164));
  XNOR2_X1  g074(.A(KEYINPUT6), .B(G651), .ZN(new_n500));
  XNOR2_X1  g075(.A(KEYINPUT5), .B(G543), .ZN(new_n501));
  AND3_X1   g076(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT72), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT72), .B1(new_n500), .B2(new_n501), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G88), .ZN(new_n505));
  NAND2_X1  g080(.A1(G75), .A2(G543), .ZN(new_n506));
  XNOR2_X1  g081(.A(new_n506), .B(KEYINPUT73), .ZN(new_n507));
  INV_X1    g082(.A(G62), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n507), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n512), .A2(G651), .B1(G50), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n505), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND3_X1  g095(.A1(new_n501), .A2(G63), .A3(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n500), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G51), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n524), .A2(KEYINPUT74), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n504), .A2(G89), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XOR2_X1   g102(.A(new_n527), .B(KEYINPUT7), .Z(new_n528));
  AOI21_X1  g103(.A(new_n528), .B1(new_n524), .B2(KEYINPUT74), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n525), .A2(new_n526), .A3(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  AOI22_X1  g106(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G651), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n535));
  INV_X1    g110(.A(new_n516), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n514), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n535), .B1(new_n537), .B2(new_n511), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT72), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n538), .A2(G90), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n517), .A2(G52), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT75), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n540), .A2(KEYINPUT75), .A3(new_n541), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n534), .B1(new_n544), .B2(new_n545), .ZN(G171));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n511), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n549), .A2(G651), .B1(G43), .B2(new_n517), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n538), .A2(G81), .A3(new_n539), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT76), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OR3_X1    g135(.A1(new_n522), .A2(KEYINPUT9), .A3(new_n560), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT9), .B1(new_n522), .B2(new_n560), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n511), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n561), .A2(new_n562), .B1(G651), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT77), .B1(new_n502), .B2(new_n503), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n538), .A2(new_n568), .A3(new_n539), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(G91), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(new_n545), .ZN(new_n572));
  AOI21_X1  g147(.A(KEYINPUT75), .B1(new_n540), .B2(new_n541), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n572), .A2(new_n573), .B1(new_n533), .B2(new_n532), .ZN(G301));
  NAND3_X1  g149(.A1(new_n567), .A2(G87), .A3(new_n569), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n501), .A2(G74), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(new_n517), .B2(G49), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(G288));
  NAND3_X1  g153(.A1(new_n567), .A2(G86), .A3(new_n569), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n511), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(G48), .B2(new_n517), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n579), .A2(new_n583), .ZN(G305));
  NAND2_X1  g159(.A1(G72), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G60), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n511), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G651), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n538), .A2(G85), .A3(new_n539), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT78), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n517), .A2(G47), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n590), .B1(new_n589), .B2(new_n591), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n588), .B1(new_n592), .B2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n567), .A2(G92), .A3(new_n569), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n567), .A2(KEYINPUT10), .A3(G92), .A4(new_n569), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n501), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT79), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n533), .B1(new_n601), .B2(new_n602), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n603), .A2(new_n604), .B1(G54), .B2(new_n517), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n595), .B1(new_n607), .B2(G868), .ZN(G284));
  XOR2_X1   g183(.A(G284), .B(KEYINPUT80), .Z(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G299), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G297));
  OAI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(new_n614), .B2(G860), .ZN(G148));
  NOR2_X1   g190(.A1(new_n552), .A2(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n607), .A2(new_n614), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n616), .B1(new_n619), .B2(G868), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n492), .A2(new_n475), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(G2100), .Z(new_n626));
  AND2_X1   g201(.A1(new_n487), .A2(G135), .ZN(new_n627));
  INV_X1    g202(.A(G123), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n471), .A2(G111), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  OAI22_X1  g205(.A1(new_n482), .A2(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(G2096), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(G2096), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n626), .A2(new_n634), .A3(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT84), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2451), .ZN(new_n639));
  XOR2_X1   g214(.A(G1341), .B(G1348), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(new_n646), .A3(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n641), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2454), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n648), .A2(new_n650), .ZN(new_n652));
  AND3_X1   g227(.A1(new_n651), .A2(G14), .A3(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2072), .B(G2078), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT17), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n657), .B2(new_n654), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n658), .B1(KEYINPUT85), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n661), .B1(KEYINPUT85), .B2(new_n660), .ZN(new_n662));
  INV_X1    g237(.A(new_n654), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n663), .A2(new_n659), .A3(new_n656), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT18), .Z(new_n665));
  NAND3_X1  g240(.A1(new_n655), .A2(new_n659), .A3(new_n657), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n662), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2096), .B(G2100), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(G1971), .B(G1976), .Z(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1956), .B(G2474), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT20), .Z(new_n678));
  NAND2_X1  g253(.A1(new_n673), .A2(new_n674), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n672), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n672), .A2(new_n679), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n678), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G229));
  OAI21_X1  g263(.A(KEYINPUT97), .B1(G16), .B2(G21), .ZN(new_n689));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NOR2_X1   g265(.A1(G286), .A2(new_n690), .ZN(new_n691));
  MUX2_X1   g266(.A(new_n689), .B(KEYINPUT97), .S(new_n691), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT98), .ZN(new_n693));
  INV_X1    g268(.A(G1966), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT100), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n693), .A2(new_n694), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT31), .B(G11), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT30), .B(G28), .Z(new_n699));
  XOR2_X1   g274(.A(KEYINPUT87), .B(G29), .Z(new_n700));
  OAI221_X1 g275(.A(new_n698), .B1(G29), .B2(new_n699), .C1(new_n633), .C2(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT99), .Z(new_n702));
  INV_X1    g277(.A(G1961), .ZN(new_n703));
  NOR2_X1   g278(.A1(G171), .A2(new_n690), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G5), .B2(new_n690), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n702), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n697), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n696), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(KEYINPUT101), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT101), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n696), .A2(new_n710), .A3(new_n707), .ZN(new_n711));
  INV_X1    g286(.A(new_n700), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n712), .A2(G35), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G162), .B2(new_n712), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT29), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G2090), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G33), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT25), .Z(new_n720));
  INV_X1    g295(.A(G139), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n492), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n722));
  OAI221_X1 g297(.A(new_n720), .B1(new_n486), .B2(new_n721), .C1(new_n471), .C2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT95), .Z(new_n724));
  OAI21_X1  g299(.A(new_n718), .B1(new_n724), .B2(new_n717), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(G2072), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(G2072), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n690), .A2(G19), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n553), .B2(new_n690), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(G1341), .Z(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT24), .B(G34), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n700), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT96), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n477), .B2(new_n717), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G2084), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n726), .A2(new_n727), .A3(new_n730), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n690), .A2(G20), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT23), .Z(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G299), .B2(G16), .ZN(new_n739));
  INV_X1    g314(.A(G1956), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n717), .A2(G32), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT26), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n745), .A2(new_n746), .B1(G105), .B2(new_n475), .ZN(new_n747));
  INV_X1    g322(.A(G129), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n482), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n487), .B2(G141), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n742), .B1(new_n750), .B2(new_n717), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT27), .B(G1996), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n700), .A2(G27), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G164), .B2(new_n700), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(G2078), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  OR3_X1    g332(.A1(new_n736), .A2(new_n741), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n607), .A2(G16), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G4), .B2(G16), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT93), .B(G1348), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n705), .A2(new_n703), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n700), .A2(G26), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT28), .ZN(new_n765));
  INV_X1    g340(.A(G128), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n471), .A2(G116), .ZN(new_n767));
  OAI21_X1  g342(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n768));
  OAI22_X1  g343(.A1(new_n482), .A2(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n487), .B2(G140), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n765), .B1(new_n770), .B2(new_n717), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT94), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G2067), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n762), .A2(new_n763), .A3(new_n773), .ZN(new_n774));
  NOR3_X1   g349(.A1(new_n716), .A2(new_n758), .A3(new_n774), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n709), .A2(new_n711), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n690), .A2(G23), .ZN(new_n777));
  INV_X1    g352(.A(G288), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(new_n690), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n779), .A2(KEYINPUT91), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n779), .A2(KEYINPUT91), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT33), .B(G1976), .Z(new_n782));
  OR3_X1    g357(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n690), .A2(G22), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G166), .B2(new_n690), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1971), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n690), .A2(G6), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G305), .B2(G16), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT32), .B(G1981), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n788), .A2(new_n790), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n786), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n782), .B1(new_n780), .B2(new_n781), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n783), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT92), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT34), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n487), .A2(G131), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT88), .Z(new_n802));
  OAI21_X1  g377(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n803));
  INV_X1    g378(.A(G107), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(G2105), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n483), .B2(G119), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  MUX2_X1   g382(.A(G25), .B(new_n807), .S(new_n712), .Z(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT89), .Z(new_n809));
  XOR2_X1   g384(.A(KEYINPUT35), .B(G1991), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT90), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n809), .A2(new_n812), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n690), .A2(G24), .ZN(new_n815));
  INV_X1    g390(.A(G290), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(new_n690), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1986), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n813), .A2(new_n814), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n799), .A2(new_n800), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT36), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT36), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n799), .A2(new_n822), .A3(new_n800), .A4(new_n819), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n776), .B1(new_n821), .B2(new_n823), .ZN(G311));
  NAND2_X1  g399(.A1(new_n821), .A2(new_n823), .ZN(new_n825));
  INV_X1    g400(.A(new_n776), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(G150));
  NAND2_X1  g402(.A1(G80), .A2(G543), .ZN(new_n828));
  INV_X1    g403(.A(G67), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n511), .B2(new_n829), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n830), .A2(G651), .B1(G55), .B2(new_n517), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n538), .A2(G93), .A3(new_n539), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G860), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT37), .Z(new_n835));
  NOR2_X1   g410(.A1(new_n606), .A2(new_n614), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT103), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n836), .B(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n552), .A2(new_n833), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n550), .A2(new_n831), .A3(new_n551), .A4(new_n832), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n839), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n844), .A2(KEYINPUT39), .ZN(new_n845));
  INV_X1    g420(.A(G860), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n844), .B2(KEYINPUT39), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n835), .B1(new_n845), .B2(new_n847), .ZN(G145));
  XNOR2_X1  g423(.A(new_n770), .B(G164), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n750), .ZN(new_n850));
  MUX2_X1   g425(.A(new_n723), .B(new_n724), .S(new_n850), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n483), .A2(G130), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT104), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n853), .A2(new_n471), .A3(G118), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n471), .B2(G118), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n855), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n852), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(G142), .B2(new_n487), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n624), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n807), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n851), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n632), .B(new_n477), .ZN(new_n862));
  XNOR2_X1  g437(.A(G162), .B(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(G37), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n863), .B2(new_n861), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g441(.A1(G305), .A2(G303), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  AOI22_X1  g443(.A1(new_n579), .A2(new_n583), .B1(new_n505), .B2(new_n518), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT106), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n868), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(KEYINPUT106), .B1(new_n867), .B2(new_n869), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT105), .ZN(new_n874));
  NAND2_X1  g449(.A1(G288), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n575), .A2(KEYINPUT105), .A3(new_n577), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(G290), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(G290), .B1(new_n875), .B2(new_n876), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n872), .B(new_n873), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n879), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n867), .A2(KEYINPUT106), .A3(new_n869), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(new_n882), .A3(new_n877), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n884), .A2(KEYINPUT42), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n880), .A2(new_n883), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT107), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n885), .B(new_n888), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n840), .A2(new_n841), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n619), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n617), .B(KEYINPUT81), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n842), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n600), .A2(new_n611), .A3(new_n605), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n611), .B1(new_n600), .B2(new_n605), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n606), .A2(G299), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n600), .A2(new_n611), .A3(new_n605), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n899), .A2(KEYINPUT41), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n894), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n896), .A2(new_n897), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n906), .B1(new_n891), .B2(new_n893), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT108), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n907), .B1(new_n894), .B2(new_n903), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n889), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n911), .A2(new_n889), .ZN(new_n913));
  OAI21_X1  g488(.A(G868), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G868), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n833), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(G295));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n916), .ZN(G331));
  NAND2_X1  g493(.A1(new_n890), .A2(G301), .ZN(new_n919));
  NAND2_X1  g494(.A1(G171), .A2(new_n842), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(new_n920), .A3(G168), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n890), .A2(G301), .ZN(new_n922));
  NOR2_X1   g497(.A1(G171), .A2(new_n842), .ZN(new_n923));
  OAI21_X1  g498(.A(G286), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n898), .A2(new_n901), .A3(new_n921), .A4(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n921), .ZN(new_n926));
  AOI21_X1  g501(.A(G168), .B1(new_n919), .B2(new_n920), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n905), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n884), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n925), .A2(new_n928), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n886), .ZN(new_n932));
  INV_X1    g507(.A(G37), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n930), .B1(new_n934), .B2(KEYINPUT110), .ZN(new_n935));
  XNOR2_X1  g510(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n932), .A2(new_n938), .A3(new_n933), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n935), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n932), .A2(new_n929), .A3(new_n933), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n936), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n935), .A2(new_n946), .A3(new_n936), .A4(new_n939), .ZN(new_n947));
  AOI22_X1  g522(.A1(new_n925), .A2(new_n928), .B1(new_n883), .B2(new_n880), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT110), .B1(new_n948), .B2(G37), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n939), .A2(new_n949), .A3(new_n936), .A4(new_n929), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT111), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT44), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT112), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n957));
  AOI211_X1 g532(.A(new_n957), .B(new_n954), .C1(new_n947), .C2(new_n951), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n945), .B1(new_n956), .B2(new_n958), .ZN(G397));
  INV_X1    g534(.A(G1384), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(new_n494), .B2(new_n498), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n468), .A2(G40), .A3(new_n474), .A4(new_n476), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n962), .A2(KEYINPUT45), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n750), .B(G1996), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n770), .B(G2067), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n968), .A2(new_n812), .A3(new_n802), .A4(new_n806), .ZN(new_n969));
  INV_X1    g544(.A(G2067), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n770), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n965), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G1996), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n964), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT46), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n967), .A2(new_n750), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n975), .B1(new_n965), .B2(new_n976), .ZN(new_n977));
  XOR2_X1   g552(.A(new_n977), .B(KEYINPUT47), .Z(new_n978));
  NOR3_X1   g553(.A1(new_n965), .A2(G1986), .A3(G290), .ZN(new_n979));
  OR2_X1    g554(.A1(new_n979), .A2(KEYINPUT48), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n807), .B(new_n812), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n968), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n982), .A2(new_n964), .B1(new_n979), .B2(KEYINPUT48), .ZN(new_n983));
  AOI211_X1 g558(.A(new_n972), .B(new_n978), .C1(new_n980), .C2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT127), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n984), .B(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT62), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n963), .B1(new_n961), .B2(KEYINPUT50), .ZN(new_n988));
  INV_X1    g563(.A(G2084), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n990), .B(new_n960), .C1(new_n494), .C2(new_n498), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n988), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n962), .A2(KEYINPUT45), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n963), .B1(new_n961), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n992), .B(G168), .C1(new_n997), .C2(G1966), .ZN(new_n998));
  INV_X1    g573(.A(new_n992), .ZN(new_n999));
  AOI21_X1  g574(.A(G1966), .B1(new_n993), .B2(new_n995), .ZN(new_n1000));
  OAI21_X1  g575(.A(G286), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n998), .A2(new_n1001), .A3(G8), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT51), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT123), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n998), .A2(new_n1005), .A3(G8), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1003), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1004), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n987), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1009), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1011), .A2(KEYINPUT62), .A3(new_n1007), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n778), .A2(G1976), .ZN(new_n1013));
  XOR2_X1   g588(.A(KEYINPUT114), .B(G1976), .Z(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT52), .B1(G288), .B2(new_n1014), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n961), .A2(new_n963), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1013), .A2(new_n1015), .A3(G8), .A4(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(G8), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1018), .B1(G1976), .B2(new_n778), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1017), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1981), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n579), .A2(new_n1022), .A3(new_n583), .ZN(new_n1023));
  INV_X1    g598(.A(new_n583), .ZN(new_n1024));
  XOR2_X1   g599(.A(KEYINPUT115), .B(G86), .Z(new_n1025));
  NOR3_X1   g600(.A1(new_n502), .A2(new_n503), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(G1981), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1023), .A2(KEYINPUT49), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT49), .B1(new_n1023), .B2(new_n1027), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n1028), .A2(new_n1029), .A3(new_n1018), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1021), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(G303), .A2(G8), .ZN(new_n1032));
  XOR2_X1   g607(.A(new_n1032), .B(KEYINPUT55), .Z(new_n1033));
  AOI21_X1  g608(.A(G1971), .B1(new_n993), .B2(new_n995), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n988), .A2(new_n991), .ZN(new_n1035));
  OAI22_X1  g610(.A1(new_n1034), .A2(KEYINPUT113), .B1(G2090), .B2(new_n1035), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1034), .A2(KEYINPUT113), .ZN(new_n1037));
  OAI211_X1 g612(.A(G8), .B(new_n1033), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G8), .ZN(new_n1039));
  INV_X1    g614(.A(G2090), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n991), .B(KEYINPUT117), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n988), .A2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n988), .A2(new_n1042), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1040), .B(new_n1041), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1034), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1039), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1031), .B(new_n1038), .C1(new_n1033), .C2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n996), .A2(G2078), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n1049), .A2(KEYINPUT53), .B1(new_n1035), .B2(new_n703), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT124), .B1(new_n1049), .B2(KEYINPUT53), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT124), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1052), .B(new_n1053), .C1(new_n996), .C2(G2078), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1050), .A2(new_n1051), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G171), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1048), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1010), .A2(new_n1012), .A3(new_n1057), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1030), .A2(G1976), .A3(G288), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1023), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1031), .ZN(new_n1062));
  OAI22_X1  g637(.A1(new_n1061), .A2(new_n1018), .B1(new_n1062), .B2(new_n1038), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT63), .ZN(new_n1064));
  OAI211_X1 g639(.A(G8), .B(G168), .C1(new_n999), .C2(new_n1000), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1064), .B1(new_n1048), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(G8), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1033), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1065), .A2(new_n1064), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1069), .A2(new_n1031), .A3(new_n1038), .A4(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1063), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1041), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT56), .B(G2072), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1073), .A2(new_n740), .B1(new_n997), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1077), .B1(new_n566), .B2(new_n570), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1075), .A2(KEYINPUT118), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT118), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1035), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(G1348), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1016), .A2(G2067), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n607), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n611), .A2(new_n1077), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1078), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT119), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n1075), .A2(new_n1093), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1081), .A2(new_n1083), .B1(new_n1087), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT60), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1097));
  OAI221_X1 g672(.A(KEYINPUT60), .B1(G2067), .B2(new_n1016), .C1(new_n1084), .C2(G1348), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(new_n607), .A3(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1100), .A2(KEYINPUT60), .A3(new_n606), .ZN(new_n1101));
  NOR2_X1   g676(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT58), .B(G1341), .Z(new_n1103));
  NAND2_X1  g678(.A1(new_n1016), .A2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n996), .B2(G1996), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1102), .B1(new_n1105), .B2(new_n553), .ZN(new_n1106));
  NAND2_X1  g681(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1107));
  XOR2_X1   g682(.A(new_n1107), .B(KEYINPUT121), .Z(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  AOI211_X1 g685(.A(new_n1102), .B(new_n1108), .C1(new_n1105), .C2(new_n553), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1099), .B(new_n1101), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1075), .A2(KEYINPUT122), .A3(new_n1079), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT61), .B1(new_n1075), .B2(new_n1093), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1075), .A2(new_n1079), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1112), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  OAI22_X1  g694(.A1(new_n1080), .A2(new_n1082), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1095), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1050), .A2(new_n1051), .A3(G301), .A4(new_n1054), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT54), .B1(new_n1056), .B2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1125), .A2(new_n1048), .ZN(new_n1126));
  NAND2_X1  g701(.A1(G171), .A2(KEYINPUT125), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n1129));
  OAI221_X1 g704(.A(KEYINPUT54), .B1(new_n1055), .B2(new_n1128), .C1(new_n1056), .C2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1126), .A2(new_n1011), .A3(new_n1007), .A4(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1058), .B(new_n1072), .C1(new_n1123), .C2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT126), .ZN(new_n1133));
  XNOR2_X1  g708(.A(G290), .B(G1986), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n964), .B1(new_n982), .B2(new_n1134), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1132), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1133), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n986), .B1(new_n1136), .B2(new_n1137), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g713(.A(new_n458), .ZN(new_n1140));
  OR2_X1    g714(.A1(G227), .A2(new_n1140), .ZN(new_n1141));
  NOR3_X1   g715(.A1(G229), .A2(G401), .A3(new_n1141), .ZN(new_n1142));
  AND2_X1   g716(.A1(new_n1142), .A2(new_n865), .ZN(new_n1143));
  NAND2_X1  g717(.A1(new_n1143), .A2(new_n943), .ZN(G225));
  INV_X1    g718(.A(G225), .ZN(G308));
endmodule


