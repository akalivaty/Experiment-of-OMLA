

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769;

  NOR2_X1 U371 ( .A1(G953), .A2(G237), .ZN(n496) );
  XNOR2_X1 U372 ( .A(n758), .B(n412), .ZN(n458) );
  INV_X2 U373 ( .A(G953), .ZN(n760) );
  XOR2_X1 U374 ( .A(KEYINPUT91), .B(G119), .Z(n349) );
  AND2_X1 U375 ( .A1(n392), .A2(n385), .ZN(n395) );
  NAND2_X1 U376 ( .A1(n725), .A2(n720), .ZN(n638) );
  INV_X1 U377 ( .A(n409), .ZN(n473) );
  BUF_X1 U378 ( .A(n737), .Z(n743) );
  NOR2_X1 U379 ( .A1(n362), .A2(n562), .ZN(n360) );
  INV_X1 U380 ( .A(n542), .ZN(n350) );
  AND2_X1 U381 ( .A1(n589), .A2(n590), .ZN(n378) );
  INV_X1 U382 ( .A(n447), .ZN(n548) );
  XNOR2_X1 U383 ( .A(n458), .B(n419), .ZN(n733) );
  XNOR2_X1 U384 ( .A(n466), .B(n465), .ZN(n749) );
  XOR2_X1 U385 ( .A(G113), .B(G104), .Z(n493) );
  XOR2_X1 U386 ( .A(G122), .B(G107), .Z(n512) );
  NOR2_X1 U387 ( .A1(n629), .A2(n549), .ZN(n370) );
  XNOR2_X1 U388 ( .A(G128), .B(G119), .ZN(n424) );
  XNOR2_X1 U389 ( .A(G146), .B(G125), .ZN(n472) );
  NAND2_X1 U390 ( .A1(n381), .A2(n380), .ZN(n681) );
  INV_X1 U391 ( .A(n750), .ZN(n381) );
  NAND2_X1 U392 ( .A1(n366), .A2(n365), .ZN(n369) );
  INV_X1 U393 ( .A(KEYINPUT0), .ZN(n394) );
  AND2_X1 U394 ( .A1(n573), .A2(n572), .ZN(n604) );
  XNOR2_X1 U395 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U396 ( .A(n518), .B(G478), .ZN(n555) );
  NAND2_X1 U397 ( .A1(n767), .A2(n713), .ZN(n542) );
  NAND2_X1 U398 ( .A1(n373), .A2(KEYINPUT84), .ZN(n372) );
  AND2_X1 U399 ( .A1(n377), .A2(n375), .ZN(n374) );
  OR2_X1 U400 ( .A1(G237), .A2(G902), .ZN(n485) );
  NAND2_X1 U401 ( .A1(n411), .A2(n410), .ZN(n513) );
  XNOR2_X1 U402 ( .A(n397), .B(n396), .ZN(n478) );
  XNOR2_X1 U403 ( .A(n473), .B(n475), .ZN(n396) );
  XNOR2_X1 U404 ( .A(n474), .B(n352), .ZN(n397) );
  NOR2_X1 U405 ( .A1(n569), .A2(n586), .ZN(n570) );
  XNOR2_X1 U406 ( .A(KEYINPUT15), .B(G902), .ZN(n676) );
  INV_X1 U407 ( .A(n633), .ZN(n391) );
  NOR2_X1 U408 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U409 ( .A(n420), .B(G469), .ZN(n552) );
  NOR2_X1 U410 ( .A1(n733), .A2(G902), .ZN(n420) );
  XNOR2_X1 U411 ( .A(n552), .B(KEYINPUT1), .ZN(n528) );
  INV_X1 U412 ( .A(KEYINPUT48), .ZN(n620) );
  XNOR2_X1 U413 ( .A(G116), .B(G101), .ZN(n448) );
  XNOR2_X1 U414 ( .A(KEYINPUT24), .B(G137), .ZN(n431) );
  XNOR2_X1 U415 ( .A(G110), .B(KEYINPUT23), .ZN(n423) );
  XNOR2_X1 U416 ( .A(G143), .B(G122), .ZN(n494) );
  XOR2_X1 U417 ( .A(G131), .B(KEYINPUT103), .Z(n498) );
  XNOR2_X1 U418 ( .A(n472), .B(n429), .ZN(n759) );
  XNOR2_X1 U419 ( .A(KEYINPUT10), .B(G140), .ZN(n429) );
  XOR2_X1 U420 ( .A(KEYINPUT79), .B(G140), .Z(n416) );
  XNOR2_X1 U421 ( .A(G101), .B(G110), .ZN(n415) );
  XOR2_X1 U422 ( .A(G107), .B(G104), .Z(n414) );
  OR2_X1 U423 ( .A1(n702), .A2(G902), .ZN(n439) );
  INV_X1 U424 ( .A(G902), .ZN(n459) );
  BUF_X1 U425 ( .A(n552), .Z(n586) );
  XNOR2_X1 U426 ( .A(n370), .B(KEYINPUT34), .ZN(n519) );
  NAND2_X1 U427 ( .A1(n384), .A2(n556), .ZN(n725) );
  AND2_X1 U428 ( .A1(n392), .A2(n356), .ZN(n351) );
  NAND2_X1 U429 ( .A1(n369), .A2(n367), .ZN(n629) );
  AND2_X1 U430 ( .A1(G224), .A2(n760), .ZN(n352) );
  AND2_X1 U431 ( .A1(n706), .A2(n559), .ZN(n353) );
  BUF_X1 U432 ( .A(n528), .Z(n645) );
  AND2_X1 U433 ( .A1(n718), .A2(n592), .ZN(n354) );
  AND2_X1 U434 ( .A1(n731), .A2(n729), .ZN(n355) );
  AND2_X1 U435 ( .A1(n388), .A2(n390), .ZN(n356) );
  XOR2_X1 U436 ( .A(KEYINPUT109), .B(KEYINPUT33), .Z(n357) );
  XNOR2_X1 U437 ( .A(KEYINPUT62), .B(n684), .ZN(n358) );
  XNOR2_X2 U438 ( .A(n359), .B(n563), .ZN(n750) );
  NAND2_X1 U439 ( .A1(n361), .A2(n360), .ZN(n359) );
  NAND2_X1 U440 ( .A1(n363), .A2(n364), .ZN(n361) );
  NAND2_X1 U441 ( .A1(n560), .A2(n353), .ZN(n362) );
  NAND2_X1 U442 ( .A1(n541), .A2(n540), .ZN(n363) );
  NAND2_X1 U443 ( .A1(n538), .A2(n537), .ZN(n364) );
  INV_X1 U444 ( .A(n357), .ZN(n365) );
  NAND2_X1 U445 ( .A1(n548), .A2(n595), .ZN(n366) );
  NAND2_X1 U446 ( .A1(n548), .A2(n368), .ZN(n367) );
  AND2_X1 U447 ( .A1(n595), .A2(n357), .ZN(n368) );
  XNOR2_X2 U448 ( .A(n395), .B(n394), .ZN(n549) );
  XNOR2_X2 U449 ( .A(n513), .B(n371), .ZN(n758) );
  INV_X1 U450 ( .A(n407), .ZN(n371) );
  OR2_X2 U451 ( .A1(n718), .A2(n591), .ZN(n589) );
  NOR2_X1 U452 ( .A1(n376), .A2(n354), .ZN(n375) );
  XNOR2_X1 U453 ( .A(n621), .B(n620), .ZN(n628) );
  NAND2_X1 U454 ( .A1(n628), .A2(n355), .ZN(n382) );
  XNOR2_X2 U455 ( .A(G128), .B(G143), .ZN(n409) );
  NAND2_X1 U456 ( .A1(n473), .A2(n408), .ZN(n411) );
  NAND2_X1 U457 ( .A1(n374), .A2(n372), .ZN(n593) );
  INV_X1 U458 ( .A(n379), .ZN(n373) );
  NOR2_X1 U459 ( .A1(n589), .A2(n590), .ZN(n376) );
  NAND2_X1 U460 ( .A1(n379), .A2(n378), .ZN(n377) );
  XNOR2_X1 U461 ( .A(n579), .B(n578), .ZN(n379) );
  NAND2_X1 U462 ( .A1(n382), .A2(n673), .ZN(n398) );
  INV_X1 U463 ( .A(n382), .ZN(n380) );
  XNOR2_X1 U464 ( .A(n382), .B(n762), .ZN(n761) );
  NAND2_X1 U465 ( .A1(n383), .A2(n555), .ZN(n720) );
  INV_X1 U466 ( .A(n556), .ZN(n383) );
  INV_X1 U467 ( .A(n555), .ZN(n384) );
  AND2_X1 U468 ( .A1(n388), .A2(n386), .ZN(n385) );
  NOR2_X1 U469 ( .A1(n492), .A2(n387), .ZN(n386) );
  INV_X1 U470 ( .A(n390), .ZN(n387) );
  NAND2_X1 U471 ( .A1(n625), .A2(n389), .ZN(n388) );
  NOR2_X1 U472 ( .A1(n391), .A2(n486), .ZN(n389) );
  NAND2_X1 U473 ( .A1(n486), .A2(n391), .ZN(n390) );
  NAND2_X1 U474 ( .A1(n393), .A2(n486), .ZN(n392) );
  INV_X1 U475 ( .A(n625), .ZN(n393) );
  AND2_X1 U476 ( .A1(n398), .A2(n674), .ZN(n399) );
  NAND2_X1 U477 ( .A1(n750), .A2(n673), .ZN(n400) );
  NAND2_X1 U478 ( .A1(n400), .A2(n399), .ZN(n678) );
  XNOR2_X2 U479 ( .A(n533), .B(n532), .ZN(n767) );
  NOR2_X1 U480 ( .A1(n638), .A2(n591), .ZN(n576) );
  XNOR2_X1 U481 ( .A(n453), .B(n452), .ZN(n454) );
  INV_X1 U482 ( .A(KEYINPUT66), .ZN(n543) );
  XNOR2_X1 U483 ( .A(n455), .B(n454), .ZN(n456) );
  NOR2_X1 U484 ( .A1(n602), .A2(n727), .ZN(n619) );
  NAND2_X1 U485 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U486 ( .A1(n534), .A2(n529), .ZN(n531) );
  XNOR2_X1 U487 ( .A(n508), .B(n507), .ZN(n556) );
  INV_X1 U488 ( .A(n747), .ZN(n687) );
  NAND2_X1 U489 ( .A1(n604), .A2(n575), .ZN(n700) );
  XNOR2_X1 U490 ( .A(n672), .B(n671), .ZN(G75) );
  INV_X1 U491 ( .A(G137), .ZN(n401) );
  NAND2_X1 U492 ( .A1(n401), .A2(KEYINPUT4), .ZN(n404) );
  INV_X1 U493 ( .A(KEYINPUT4), .ZN(n402) );
  NAND2_X1 U494 ( .A1(n402), .A2(G137), .ZN(n403) );
  NAND2_X1 U495 ( .A1(n404), .A2(n403), .ZN(n406) );
  XNOR2_X1 U496 ( .A(G131), .B(KEYINPUT70), .ZN(n405) );
  XNOR2_X1 U497 ( .A(n406), .B(n405), .ZN(n407) );
  INV_X1 U498 ( .A(G134), .ZN(n408) );
  NAND2_X1 U499 ( .A1(n409), .A2(G134), .ZN(n410) );
  INV_X1 U500 ( .A(G146), .ZN(n412) );
  NAND2_X1 U501 ( .A1(G227), .A2(n760), .ZN(n413) );
  XNOR2_X1 U502 ( .A(n414), .B(n413), .ZN(n418) );
  XNOR2_X1 U503 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U504 ( .A(n418), .B(n417), .Z(n419) );
  INV_X1 U505 ( .A(n528), .ZN(n445) );
  NAND2_X1 U506 ( .A1(n760), .A2(G234), .ZN(n422) );
  XNOR2_X1 U507 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n421) );
  XNOR2_X1 U508 ( .A(n422), .B(n421), .ZN(n509) );
  NAND2_X1 U509 ( .A1(n509), .A2(G221), .ZN(n428) );
  XNOR2_X1 U510 ( .A(n424), .B(n423), .ZN(n426) );
  XNOR2_X1 U511 ( .A(KEYINPUT97), .B(KEYINPUT78), .ZN(n425) );
  XNOR2_X1 U512 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U513 ( .A(n428), .B(n427), .ZN(n434) );
  XNOR2_X1 U514 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n430) );
  XNOR2_X1 U515 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U516 ( .A(n759), .B(n432), .ZN(n433) );
  XNOR2_X1 U517 ( .A(n434), .B(n433), .ZN(n702) );
  NAND2_X1 U518 ( .A1(n676), .A2(G234), .ZN(n435) );
  XNOR2_X1 U519 ( .A(n435), .B(KEYINPUT20), .ZN(n440) );
  NAND2_X1 U520 ( .A1(n440), .A2(G217), .ZN(n437) );
  XNOR2_X1 U521 ( .A(KEYINPUT77), .B(KEYINPUT25), .ZN(n436) );
  XNOR2_X1 U522 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X2 U523 ( .A(n439), .B(n438), .ZN(n544) );
  NAND2_X1 U524 ( .A1(n440), .A2(G221), .ZN(n443) );
  XOR2_X1 U525 ( .A(KEYINPUT21), .B(KEYINPUT98), .Z(n441) );
  XNOR2_X1 U526 ( .A(KEYINPUT99), .B(n441), .ZN(n442) );
  XNOR2_X1 U527 ( .A(n443), .B(n442), .ZN(n647) );
  XOR2_X1 U528 ( .A(n647), .B(KEYINPUT100), .Z(n525) );
  NAND2_X1 U529 ( .A1(n544), .A2(n525), .ZN(n568) );
  INV_X1 U530 ( .A(n568), .ZN(n444) );
  NAND2_X1 U531 ( .A1(n445), .A2(n444), .ZN(n446) );
  XNOR2_X1 U532 ( .A(n446), .B(KEYINPUT74), .ZN(n447) );
  XNOR2_X1 U533 ( .A(n349), .B(n448), .ZN(n449) );
  XNOR2_X1 U534 ( .A(KEYINPUT3), .B(n449), .ZN(n462) );
  XOR2_X1 U535 ( .A(KEYINPUT75), .B(KEYINPUT101), .Z(n451) );
  NAND2_X1 U536 ( .A1(n496), .A2(G210), .ZN(n450) );
  XNOR2_X1 U537 ( .A(n451), .B(n450), .ZN(n455) );
  XNOR2_X1 U538 ( .A(G113), .B(KEYINPUT5), .ZN(n453) );
  INV_X1 U539 ( .A(KEYINPUT102), .ZN(n452) );
  XNOR2_X1 U540 ( .A(n462), .B(n456), .ZN(n457) );
  XNOR2_X1 U541 ( .A(n458), .B(n457), .ZN(n684) );
  NAND2_X1 U542 ( .A1(n684), .A2(n459), .ZN(n460) );
  XNOR2_X2 U543 ( .A(n460), .B(G472), .ZN(n651) );
  INV_X1 U544 ( .A(KEYINPUT6), .ZN(n461) );
  XNOR2_X1 U545 ( .A(n651), .B(n461), .ZN(n595) );
  INV_X1 U546 ( .A(n462), .ZN(n466) );
  XNOR2_X1 U547 ( .A(n512), .B(n493), .ZN(n464) );
  XOR2_X1 U548 ( .A(G110), .B(KEYINPUT16), .Z(n463) );
  XNOR2_X1 U549 ( .A(n464), .B(n463), .ZN(n465) );
  INV_X1 U550 ( .A(n749), .ZN(n477) );
  INV_X1 U551 ( .A(KEYINPUT18), .ZN(n467) );
  NAND2_X1 U552 ( .A1(KEYINPUT80), .A2(n467), .ZN(n470) );
  INV_X1 U553 ( .A(KEYINPUT80), .ZN(n468) );
  NAND2_X1 U554 ( .A1(n468), .A2(KEYINPUT18), .ZN(n469) );
  NAND2_X1 U555 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U556 ( .A(n472), .B(n471), .ZN(n474) );
  XNOR2_X1 U557 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n475) );
  INV_X1 U558 ( .A(n478), .ZN(n476) );
  NAND2_X1 U559 ( .A1(n477), .A2(n476), .ZN(n480) );
  NAND2_X1 U560 ( .A1(n478), .A2(n749), .ZN(n479) );
  NAND2_X1 U561 ( .A1(n480), .A2(n479), .ZN(n691) );
  NAND2_X1 U562 ( .A1(n691), .A2(n676), .ZN(n484) );
  AND2_X1 U563 ( .A1(G210), .A2(n485), .ZN(n482) );
  XOR2_X1 U564 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n481) );
  XNOR2_X1 U565 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X2 U566 ( .A(n484), .B(n483), .ZN(n625) );
  NAND2_X1 U567 ( .A1(G214), .A2(n485), .ZN(n633) );
  XOR2_X1 U568 ( .A(KEYINPUT19), .B(KEYINPUT68), .Z(n486) );
  XOR2_X1 U569 ( .A(KEYINPUT73), .B(KEYINPUT14), .Z(n488) );
  NAND2_X1 U570 ( .A1(G234), .A2(G237), .ZN(n487) );
  XNOR2_X1 U571 ( .A(n488), .B(n487), .ZN(n664) );
  NAND2_X1 U572 ( .A1(G952), .A2(n760), .ZN(n565) );
  NOR2_X1 U573 ( .A1(G898), .A2(n760), .ZN(n748) );
  NAND2_X1 U574 ( .A1(G902), .A2(n748), .ZN(n489) );
  NAND2_X1 U575 ( .A1(n565), .A2(n489), .ZN(n490) );
  NAND2_X1 U576 ( .A1(n664), .A2(n490), .ZN(n491) );
  XNOR2_X1 U577 ( .A(KEYINPUT94), .B(n491), .ZN(n492) );
  XNOR2_X1 U578 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U579 ( .A(n495), .B(n759), .Z(n504) );
  NAND2_X1 U580 ( .A1(G214), .A2(n496), .ZN(n497) );
  XNOR2_X1 U581 ( .A(n498), .B(n497), .ZN(n502) );
  XOR2_X1 U582 ( .A(KEYINPUT11), .B(KEYINPUT104), .Z(n500) );
  XNOR2_X1 U583 ( .A(KEYINPUT105), .B(KEYINPUT12), .ZN(n499) );
  XNOR2_X1 U584 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U585 ( .A(n502), .B(n501), .Z(n503) );
  XNOR2_X1 U586 ( .A(n504), .B(n503), .ZN(n738) );
  NOR2_X1 U587 ( .A1(G902), .A2(n738), .ZN(n508) );
  XNOR2_X1 U588 ( .A(KEYINPUT106), .B(KEYINPUT13), .ZN(n506) );
  INV_X1 U589 ( .A(G475), .ZN(n505) );
  XOR2_X1 U590 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n511) );
  NAND2_X1 U591 ( .A1(G217), .A2(n509), .ZN(n510) );
  XNOR2_X1 U592 ( .A(n511), .B(n510), .ZN(n517) );
  XOR2_X1 U593 ( .A(KEYINPUT107), .B(n512), .Z(n515) );
  XNOR2_X1 U594 ( .A(G116), .B(n513), .ZN(n514) );
  XNOR2_X1 U595 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U596 ( .A(n517), .B(n516), .ZN(n744) );
  NOR2_X1 U597 ( .A1(G902), .A2(n744), .ZN(n518) );
  NOR2_X1 U598 ( .A1(n556), .A2(n555), .ZN(n574) );
  NAND2_X1 U599 ( .A1(n519), .A2(n574), .ZN(n521) );
  INV_X1 U600 ( .A(KEYINPUT35), .ZN(n520) );
  XNOR2_X2 U601 ( .A(n521), .B(n520), .ZN(n561) );
  NOR2_X1 U602 ( .A1(n561), .A2(KEYINPUT89), .ZN(n523) );
  INV_X1 U603 ( .A(KEYINPUT44), .ZN(n522) );
  NOR2_X1 U604 ( .A1(n523), .A2(n522), .ZN(n538) );
  INV_X1 U605 ( .A(n549), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n556), .A2(n555), .ZN(n637) );
  INV_X1 U607 ( .A(n637), .ZN(n524) );
  AND2_X1 U608 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U609 ( .A1(n551), .A2(n526), .ZN(n527) );
  XNOR2_X1 U610 ( .A(n527), .B(KEYINPUT22), .ZN(n534) );
  OR2_X1 U611 ( .A1(n645), .A2(n544), .ZN(n529) );
  XNOR2_X1 U612 ( .A(n595), .B(KEYINPUT81), .ZN(n530) );
  NAND2_X1 U613 ( .A1(n531), .A2(n530), .ZN(n533) );
  XOR2_X1 U614 ( .A(KEYINPUT67), .B(KEYINPUT32), .Z(n532) );
  INV_X1 U615 ( .A(n534), .ZN(n547) );
  NOR2_X1 U616 ( .A1(n651), .A2(n544), .ZN(n535) );
  AND2_X1 U617 ( .A1(n645), .A2(n535), .ZN(n536) );
  NAND2_X1 U618 ( .A1(n547), .A2(n536), .ZN(n713) );
  NAND2_X1 U619 ( .A1(n542), .A2(KEYINPUT66), .ZN(n537) );
  NAND2_X1 U620 ( .A1(n350), .A2(n561), .ZN(n541) );
  NOR2_X1 U621 ( .A1(KEYINPUT89), .A2(KEYINPUT44), .ZN(n539) );
  AND2_X1 U622 ( .A1(n539), .A2(KEYINPUT66), .ZN(n540) );
  NAND2_X1 U623 ( .A1(n350), .A2(n543), .ZN(n560) );
  INV_X1 U624 ( .A(n544), .ZN(n648) );
  NOR2_X1 U625 ( .A1(n595), .A2(n648), .ZN(n545) );
  AND2_X1 U626 ( .A1(n545), .A2(n645), .ZN(n546) );
  NAND2_X1 U627 ( .A1(n547), .A2(n546), .ZN(n706) );
  NAND2_X1 U628 ( .A1(n548), .A2(n651), .ZN(n656) );
  NOR2_X1 U629 ( .A1(n656), .A2(n549), .ZN(n550) );
  XNOR2_X1 U630 ( .A(n550), .B(KEYINPUT31), .ZN(n724) );
  INV_X1 U631 ( .A(n651), .ZN(n583) );
  NAND2_X1 U632 ( .A1(n583), .A2(n444), .ZN(n553) );
  NOR2_X1 U633 ( .A1(n553), .A2(n586), .ZN(n554) );
  NAND2_X1 U634 ( .A1(n551), .A2(n554), .ZN(n710) );
  NAND2_X1 U635 ( .A1(n724), .A2(n710), .ZN(n557) );
  NAND2_X1 U636 ( .A1(n557), .A2(n638), .ZN(n558) );
  XNOR2_X1 U637 ( .A(n558), .B(KEYINPUT108), .ZN(n559) );
  AND2_X1 U638 ( .A1(n561), .A2(KEYINPUT89), .ZN(n562) );
  INV_X1 U639 ( .A(KEYINPUT45), .ZN(n563) );
  NOR2_X1 U640 ( .A1(G900), .A2(n760), .ZN(n564) );
  NAND2_X1 U641 ( .A1(n564), .A2(G902), .ZN(n566) );
  NAND2_X1 U642 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U643 ( .A1(n664), .A2(n567), .ZN(n580) );
  OR2_X1 U644 ( .A1(n568), .A2(n580), .ZN(n569) );
  XNOR2_X1 U645 ( .A(n570), .B(KEYINPUT76), .ZN(n573) );
  AND2_X1 U646 ( .A1(n651), .A2(n633), .ZN(n571) );
  XNOR2_X1 U647 ( .A(n571), .B(KEYINPUT30), .ZN(n572) );
  AND2_X1 U648 ( .A1(n574), .A2(n625), .ZN(n575) );
  INV_X1 U649 ( .A(KEYINPUT47), .ZN(n591) );
  XNOR2_X1 U650 ( .A(n576), .B(KEYINPUT85), .ZN(n577) );
  NAND2_X1 U651 ( .A1(n700), .A2(n577), .ZN(n579) );
  INV_X1 U652 ( .A(KEYINPUT82), .ZN(n578) );
  INV_X1 U653 ( .A(KEYINPUT28), .ZN(n585) );
  NOR2_X1 U654 ( .A1(n580), .A2(n647), .ZN(n581) );
  XOR2_X1 U655 ( .A(KEYINPUT71), .B(n581), .Z(n594) );
  NAND2_X1 U656 ( .A1(n594), .A2(n648), .ZN(n582) );
  XNOR2_X1 U657 ( .A(n585), .B(n584), .ZN(n588) );
  XOR2_X1 U658 ( .A(n586), .B(KEYINPUT111), .Z(n587) );
  NOR2_X1 U659 ( .A1(n588), .A2(n587), .ZN(n613) );
  AND2_X1 U660 ( .A1(n613), .A2(n351), .ZN(n718) );
  INV_X1 U661 ( .A(KEYINPUT84), .ZN(n590) );
  AND2_X1 U662 ( .A1(n638), .A2(n591), .ZN(n592) );
  XNOR2_X1 U663 ( .A(n593), .B(KEYINPUT72), .ZN(n602) );
  NAND2_X1 U664 ( .A1(n594), .A2(n633), .ZN(n597) );
  INV_X1 U665 ( .A(n720), .ZN(n717) );
  NAND2_X1 U666 ( .A1(n717), .A2(n595), .ZN(n596) );
  NOR2_X1 U667 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U668 ( .A1(n598), .A2(n648), .ZN(n622) );
  NAND2_X1 U669 ( .A1(n622), .A2(n625), .ZN(n600) );
  INV_X1 U670 ( .A(KEYINPUT36), .ZN(n599) );
  XNOR2_X1 U671 ( .A(n600), .B(n599), .ZN(n601) );
  AND2_X1 U672 ( .A1(n601), .A2(n445), .ZN(n727) );
  INV_X1 U673 ( .A(KEYINPUT38), .ZN(n603) );
  XNOR2_X1 U674 ( .A(n625), .B(n603), .ZN(n634) );
  NAND2_X1 U675 ( .A1(n604), .A2(n634), .ZN(n607) );
  INV_X1 U676 ( .A(KEYINPUT88), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n605), .B(KEYINPUT39), .ZN(n606) );
  XNOR2_X1 U678 ( .A(n607), .B(n606), .ZN(n627) );
  INV_X1 U679 ( .A(n627), .ZN(n608) );
  NAND2_X1 U680 ( .A1(n608), .A2(n717), .ZN(n609) );
  XNOR2_X1 U681 ( .A(n609), .B(KEYINPUT40), .ZN(n690) );
  NAND2_X1 U682 ( .A1(n634), .A2(n633), .ZN(n639) );
  NOR2_X1 U683 ( .A1(n637), .A2(n639), .ZN(n612) );
  XNOR2_X1 U684 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n610) );
  XNOR2_X1 U685 ( .A(n610), .B(KEYINPUT112), .ZN(n611) );
  XNOR2_X1 U686 ( .A(n612), .B(n611), .ZN(n630) );
  AND2_X1 U687 ( .A1(n630), .A2(n613), .ZN(n615) );
  INV_X1 U688 ( .A(KEYINPUT42), .ZN(n614) );
  XNOR2_X1 U689 ( .A(n615), .B(n614), .ZN(n769) );
  NAND2_X1 U690 ( .A1(n690), .A2(n769), .ZN(n617) );
  XOR2_X1 U691 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n616) );
  XNOR2_X1 U692 ( .A(n617), .B(n616), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n622), .B(KEYINPUT110), .ZN(n623) );
  NAND2_X1 U695 ( .A1(n623), .A2(n645), .ZN(n624) );
  XNOR2_X1 U696 ( .A(n624), .B(KEYINPUT43), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n626), .A2(n393), .ZN(n731) );
  OR2_X1 U698 ( .A1(n627), .A2(n725), .ZN(n729) );
  XNOR2_X1 U699 ( .A(n681), .B(n680), .ZN(n632) );
  INV_X1 U700 ( .A(n630), .ZN(n659) );
  OR2_X1 U701 ( .A1(n629), .A2(n659), .ZN(n631) );
  NAND2_X1 U702 ( .A1(n632), .A2(n631), .ZN(n668) );
  NOR2_X1 U703 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U704 ( .A(KEYINPUT119), .B(n635), .Z(n636) );
  NOR2_X1 U705 ( .A1(n637), .A2(n636), .ZN(n642) );
  INV_X1 U706 ( .A(n638), .ZN(n640) );
  NOR2_X1 U707 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U708 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U709 ( .A(n643), .B(KEYINPUT120), .ZN(n644) );
  NOR2_X1 U710 ( .A1(n629), .A2(n644), .ZN(n661) );
  NAND2_X1 U711 ( .A1(n645), .A2(n568), .ZN(n646) );
  XNOR2_X1 U712 ( .A(n646), .B(KEYINPUT50), .ZN(n654) );
  NAND2_X1 U713 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U714 ( .A(n649), .B(KEYINPUT49), .ZN(n650) );
  NOR2_X1 U715 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U716 ( .A(KEYINPUT118), .B(n652), .ZN(n653) );
  NAND2_X1 U717 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U718 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U719 ( .A(KEYINPUT51), .B(n657), .ZN(n658) );
  NOR2_X1 U720 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U721 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U722 ( .A(n662), .B(KEYINPUT52), .Z(n663) );
  XNOR2_X1 U723 ( .A(KEYINPUT121), .B(n663), .ZN(n666) );
  NAND2_X1 U724 ( .A1(n664), .A2(G952), .ZN(n665) );
  NOR2_X1 U725 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U726 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U727 ( .A(KEYINPUT122), .B(n669), .ZN(n670) );
  NAND2_X1 U728 ( .A1(n670), .A2(n760), .ZN(n672) );
  XNOR2_X1 U729 ( .A(KEYINPUT53), .B(KEYINPUT123), .ZN(n671) );
  NAND2_X1 U730 ( .A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(n673) );
  INV_X1 U731 ( .A(n676), .ZN(n674) );
  INV_X1 U732 ( .A(KEYINPUT2), .ZN(n680) );
  NOR2_X1 U733 ( .A1(n680), .A2(KEYINPUT86), .ZN(n675) );
  NAND2_X1 U734 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X2 U735 ( .A(n679), .B(KEYINPUT65), .ZN(n683) );
  NOR2_X1 U736 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X4 U737 ( .A1(n683), .A2(n682), .ZN(n737) );
  NAND2_X1 U738 ( .A1(n737), .A2(G472), .ZN(n685) );
  XNOR2_X1 U739 ( .A(n685), .B(n358), .ZN(n688) );
  INV_X1 U740 ( .A(G952), .ZN(n686) );
  AND2_X1 U741 ( .A1(n686), .A2(G953), .ZN(n747) );
  NAND2_X1 U742 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U743 ( .A(n689), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U744 ( .A(n690), .B(G131), .ZN(G33) );
  NAND2_X1 U745 ( .A1(n737), .A2(G210), .ZN(n696) );
  XOR2_X1 U746 ( .A(KEYINPUT90), .B(KEYINPUT54), .Z(n693) );
  XNOR2_X1 U747 ( .A(KEYINPUT55), .B(KEYINPUT83), .ZN(n692) );
  XNOR2_X1 U748 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U749 ( .A(n691), .B(n694), .ZN(n695) );
  XNOR2_X1 U750 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X2 U751 ( .A1(n697), .A2(n747), .ZN(n699) );
  XOR2_X1 U752 ( .A(KEYINPUT87), .B(KEYINPUT56), .Z(n698) );
  XNOR2_X1 U753 ( .A(n699), .B(n698), .ZN(G51) );
  XNOR2_X1 U754 ( .A(n700), .B(G143), .ZN(G45) );
  XNOR2_X1 U755 ( .A(n561), .B(G122), .ZN(G24) );
  NAND2_X1 U756 ( .A1(n743), .A2(G217), .ZN(n704) );
  XOR2_X1 U757 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n701) );
  XNOR2_X1 U758 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U759 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U760 ( .A1(n705), .A2(n747), .ZN(G66) );
  XNOR2_X1 U761 ( .A(G101), .B(n706), .ZN(G3) );
  NOR2_X1 U762 ( .A1(n720), .A2(n710), .ZN(n707) );
  XOR2_X1 U763 ( .A(G104), .B(n707), .Z(G6) );
  XOR2_X1 U764 ( .A(KEYINPUT114), .B(KEYINPUT26), .Z(n709) );
  XNOR2_X1 U765 ( .A(G107), .B(KEYINPUT27), .ZN(n708) );
  XNOR2_X1 U766 ( .A(n709), .B(n708), .ZN(n712) );
  NOR2_X1 U767 ( .A1(n725), .A2(n710), .ZN(n711) );
  XOR2_X1 U768 ( .A(n712), .B(n711), .Z(G9) );
  XNOR2_X1 U769 ( .A(G110), .B(n713), .ZN(G12) );
  XOR2_X1 U770 ( .A(G128), .B(KEYINPUT29), .Z(n716) );
  INV_X1 U771 ( .A(n718), .ZN(n714) );
  OR2_X1 U772 ( .A1(n714), .A2(n725), .ZN(n715) );
  XNOR2_X1 U773 ( .A(n716), .B(n715), .ZN(G30) );
  NAND2_X1 U774 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U775 ( .A(n719), .B(G146), .ZN(G48) );
  NOR2_X1 U776 ( .A1(n720), .A2(n724), .ZN(n722) );
  XNOR2_X1 U777 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n721) );
  XNOR2_X1 U778 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U779 ( .A(G113), .B(n723), .ZN(G15) );
  NOR2_X1 U780 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U781 ( .A(G116), .B(n726), .Z(G18) );
  XNOR2_X1 U782 ( .A(G125), .B(n727), .ZN(n728) );
  XNOR2_X1 U783 ( .A(n728), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U784 ( .A(G134), .B(n729), .Z(n730) );
  XNOR2_X1 U785 ( .A(n730), .B(KEYINPUT117), .ZN(G36) );
  XNOR2_X1 U786 ( .A(G140), .B(n731), .ZN(G42) );
  NAND2_X1 U787 ( .A1(n743), .A2(G469), .ZN(n735) );
  XOR2_X1 U788 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n732) );
  XNOR2_X1 U789 ( .A(n733), .B(n732), .ZN(n734) );
  XNOR2_X1 U790 ( .A(n735), .B(n734), .ZN(n736) );
  NOR2_X1 U791 ( .A1(n747), .A2(n736), .ZN(G54) );
  NAND2_X1 U792 ( .A1(n737), .A2(G475), .ZN(n740) );
  XOR2_X1 U793 ( .A(KEYINPUT59), .B(n738), .Z(n739) );
  XNOR2_X1 U794 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X2 U795 ( .A1(n741), .A2(n747), .ZN(n742) );
  XNOR2_X1 U796 ( .A(n742), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U797 ( .A1(n743), .A2(G478), .ZN(n745) );
  XNOR2_X1 U798 ( .A(n745), .B(n744), .ZN(n746) );
  NOR2_X1 U799 ( .A1(n747), .A2(n746), .ZN(G63) );
  NOR2_X1 U800 ( .A1(n749), .A2(n748), .ZN(n757) );
  OR2_X1 U801 ( .A1(n750), .A2(G953), .ZN(n755) );
  NAND2_X1 U802 ( .A1(G953), .A2(G224), .ZN(n751) );
  XNOR2_X1 U803 ( .A(KEYINPUT61), .B(n751), .ZN(n752) );
  NAND2_X1 U804 ( .A1(n752), .A2(G898), .ZN(n753) );
  XNOR2_X1 U805 ( .A(n753), .B(KEYINPUT126), .ZN(n754) );
  NAND2_X1 U806 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U807 ( .A(n757), .B(n756), .ZN(G69) );
  XOR2_X1 U808 ( .A(n758), .B(n759), .Z(n762) );
  NAND2_X1 U809 ( .A1(n761), .A2(n760), .ZN(n766) );
  XNOR2_X1 U810 ( .A(n762), .B(G227), .ZN(n763) );
  NAND2_X1 U811 ( .A1(n763), .A2(G900), .ZN(n764) );
  NAND2_X1 U812 ( .A1(n764), .A2(G953), .ZN(n765) );
  NAND2_X1 U813 ( .A1(n766), .A2(n765), .ZN(G72) );
  XOR2_X1 U814 ( .A(n767), .B(G119), .Z(n768) );
  XNOR2_X1 U815 ( .A(KEYINPUT127), .B(n768), .ZN(G21) );
  XNOR2_X1 U816 ( .A(G137), .B(n769), .ZN(G39) );
endmodule

