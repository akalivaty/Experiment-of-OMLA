//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT2), .B(G113), .Z(new_n188));
  XNOR2_X1  g002(.A(G116), .B(G119), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n192));
  INV_X1    g006(.A(G134), .ZN(new_n193));
  NOR3_X1   g007(.A1(new_n192), .A2(new_n193), .A3(G137), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(KEYINPUT65), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G134), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n197), .A3(G137), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n194), .B1(new_n198), .B2(KEYINPUT66), .ZN(new_n199));
  INV_X1    g013(.A(G131), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT66), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n195), .A2(new_n197), .A3(new_n201), .A4(G137), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT65), .B(G134), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n192), .B1(new_n203), .B2(G137), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n199), .A2(new_n200), .A3(new_n202), .A4(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OAI211_X1 g024(.A(KEYINPUT67), .B(KEYINPUT1), .C1(new_n208), .C2(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G128), .ZN(new_n212));
  AOI21_X1  g026(.A(KEYINPUT67), .B1(new_n207), .B2(KEYINPUT1), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n210), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT64), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(new_n206), .A3(G143), .ZN(new_n217));
  INV_X1    g031(.A(G128), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n215), .A2(new_n217), .A3(new_n209), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(G137), .B1(new_n195), .B2(new_n197), .ZN(new_n222));
  INV_X1    g036(.A(G137), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(G134), .ZN(new_n224));
  OAI21_X1  g038(.A(G131), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n205), .A2(new_n221), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n198), .A2(KEYINPUT66), .ZN(new_n228));
  INV_X1    g042(.A(new_n194), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n202), .B1(new_n222), .B2(KEYINPUT11), .ZN(new_n231));
  OAI21_X1  g045(.A(G131), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n205), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n215), .A2(new_n217), .A3(new_n209), .A4(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT0), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n218), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n210), .A2(new_n238), .A3(new_n234), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n227), .B1(new_n233), .B2(new_n241), .ZN(new_n242));
  AOI211_X1 g056(.A(KEYINPUT68), .B(new_n240), .C1(new_n232), .C2(new_n205), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n226), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT30), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n233), .A2(new_n241), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT30), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n246), .A2(new_n247), .A3(new_n226), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n191), .B1(new_n245), .B2(new_n249), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n191), .B(new_n226), .C1(new_n242), .C2(new_n243), .ZN(new_n251));
  NOR2_X1   g065(.A1(G237), .A2(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G210), .ZN(new_n253));
  XOR2_X1   g067(.A(new_n253), .B(KEYINPUT27), .Z(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(G101), .ZN(new_n255));
  XOR2_X1   g069(.A(new_n254), .B(new_n255), .Z(new_n256));
  NAND2_X1  g070(.A1(new_n251), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT31), .B1(new_n250), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n256), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n246), .A2(new_n226), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n190), .B1(new_n260), .B2(KEYINPUT69), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n246), .A2(new_n262), .A3(new_n226), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT28), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n260), .A2(new_n190), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n265), .B1(new_n251), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n259), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n257), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT31), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n248), .B1(new_n244), .B2(KEYINPUT30), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n269), .B(new_n270), .C1(new_n191), .C2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n258), .A2(new_n268), .A3(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(G472), .A2(G902), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n187), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n273), .A2(new_n187), .A3(new_n274), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n244), .A2(new_n190), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(KEYINPUT70), .A3(new_n251), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n244), .A2(new_n279), .A3(new_n190), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n278), .A2(KEYINPUT28), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n264), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n256), .A2(KEYINPUT29), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n256), .B1(new_n264), .B2(new_n267), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n251), .B(new_n259), .C1(new_n271), .C2(new_n191), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT29), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n284), .A2(new_n287), .A3(G902), .ZN(new_n288));
  INV_X1    g102(.A(G472), .ZN(new_n289));
  OAI22_X1  g103(.A1(new_n275), .A2(new_n276), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT16), .ZN(new_n293));
  INV_X1    g107(.A(G140), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n294), .A3(G125), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(G125), .ZN(new_n296));
  INV_X1    g110(.A(G125), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G140), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n295), .B1(new_n299), .B2(new_n293), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n206), .ZN(new_n301));
  OAI211_X1 g115(.A(G146), .B(new_n295), .C1(new_n299), .C2(new_n293), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT23), .B1(new_n218), .B2(G119), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n306));
  INV_X1    g120(.A(G119), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n306), .B1(new_n307), .B2(G128), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n305), .B(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G110), .ZN(new_n310));
  XOR2_X1   g124(.A(G119), .B(G128), .Z(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT24), .B(G110), .ZN(new_n312));
  OAI22_X1  g126(.A1(new_n309), .A2(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n292), .B1(new_n304), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n311), .A2(new_n312), .ZN(new_n315));
  INV_X1    g129(.A(new_n309), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n315), .B1(new_n316), .B2(G110), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(KEYINPUT73), .A3(new_n303), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n311), .A2(new_n312), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n320), .B1(new_n316), .B2(G110), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n296), .A2(new_n298), .A3(new_n206), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n302), .A3(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT22), .B(G137), .ZN(new_n324));
  INV_X1    g138(.A(G221), .ZN(new_n325));
  INV_X1    g139(.A(G234), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n325), .A2(new_n326), .A3(G953), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n324), .B(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n319), .A2(new_n323), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n329), .B1(new_n319), .B2(new_n323), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G902), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(KEYINPUT25), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n319), .A2(new_n323), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n328), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n319), .A2(new_n323), .A3(new_n329), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n333), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT25), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(G217), .B1(new_n326), .B2(G902), .ZN(new_n342));
  XOR2_X1   g156(.A(new_n342), .B(KEYINPUT71), .Z(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(new_n333), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(KEYINPUT74), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n332), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n291), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n343), .B1(new_n334), .B2(new_n340), .ZN(new_n350));
  INV_X1    g164(.A(new_n348), .ZN(new_n351));
  NOR3_X1   g165(.A1(new_n350), .A2(KEYINPUT75), .A3(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n290), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(G214), .B1(G237), .B2(G902), .ZN(new_n355));
  XNOR2_X1  g169(.A(G110), .B(G122), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT85), .B(KEYINPUT8), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT3), .ZN(new_n359));
  INV_X1    g173(.A(G104), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n359), .B1(new_n360), .B2(G107), .ZN(new_n361));
  INV_X1    g175(.A(G107), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(KEYINPUT3), .A3(G104), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G101), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT76), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n366), .B1(new_n362), .B2(G104), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n360), .A2(KEYINPUT76), .A3(G107), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n364), .A2(new_n365), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT78), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n370), .B1(new_n362), .B2(G104), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n362), .A2(G104), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n360), .A2(KEYINPUT78), .A3(G107), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G101), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n369), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n189), .A2(KEYINPUT5), .ZN(new_n377));
  INV_X1    g191(.A(G116), .ZN(new_n378));
  NOR3_X1   g192(.A1(new_n378), .A2(KEYINPUT5), .A3(G119), .ZN(new_n379));
  INV_X1    g193(.A(G113), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n377), .A2(new_n381), .B1(new_n188), .B2(new_n189), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n376), .A2(new_n382), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n358), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n364), .A2(new_n367), .A3(new_n368), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n365), .A2(KEYINPUT77), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(KEYINPUT4), .A3(new_n369), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT77), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n387), .A2(new_n391), .A3(new_n392), .A4(G101), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n390), .A2(new_n190), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n356), .A3(new_n383), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT7), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT84), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n240), .A2(new_n397), .A3(G125), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n214), .A2(new_n297), .A3(new_n220), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n397), .B1(new_n240), .B2(G125), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n396), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n386), .A2(new_n395), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G224), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(G953), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n400), .A2(new_n405), .A3(new_n401), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n396), .A2(KEYINPUT86), .ZN(new_n407));
  INV_X1    g221(.A(new_n401), .ZN(new_n408));
  NAND2_X1  g222(.A1(KEYINPUT86), .A2(KEYINPUT7), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n408), .A2(new_n399), .A3(new_n398), .A4(new_n409), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n406), .A2(new_n407), .B1(new_n410), .B2(new_n405), .ZN(new_n411));
  AOI21_X1  g225(.A(G902), .B1(new_n403), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n394), .A2(new_n383), .ZN(new_n413));
  INV_X1    g227(.A(new_n356), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(KEYINPUT6), .A3(new_n395), .ZN(new_n416));
  INV_X1    g230(.A(new_n406), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n405), .B1(new_n400), .B2(new_n401), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n413), .A2(new_n420), .A3(new_n414), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n416), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(G210), .B1(G237), .B2(G902), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n412), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n423), .B1(new_n412), .B2(new_n422), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n355), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(G234), .A2(G237), .ZN(new_n427));
  INV_X1    g241(.A(G953), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(G952), .A3(new_n428), .ZN(new_n429));
  XOR2_X1   g243(.A(new_n429), .B(KEYINPUT94), .Z(new_n430));
  NAND3_X1  g244(.A1(new_n427), .A2(G902), .A3(G953), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(G898), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(KEYINPUT9), .B(G234), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(G217), .A3(new_n428), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT92), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n441), .B1(G128), .B2(new_n208), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n218), .A2(KEYINPUT92), .A3(G143), .ZN(new_n443));
  OR2_X1    g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n218), .A2(G143), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n203), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n444), .A2(new_n203), .A3(new_n445), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OR2_X1    g264(.A1(new_n378), .A2(G122), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n362), .B1(new_n451), .B2(KEYINPUT14), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n378), .A2(G122), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n452), .B(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n450), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT93), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT13), .ZN(new_n459));
  OAI22_X1  g273(.A1(new_n442), .A2(new_n443), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(KEYINPUT93), .B2(KEYINPUT13), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n444), .A2(new_n458), .A3(new_n459), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n462), .A3(new_n445), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n463), .A2(G134), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n454), .A2(new_n362), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n451), .A2(new_n453), .A3(G107), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n449), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n440), .B(new_n457), .C1(new_n464), .C2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n467), .B1(new_n463), .B2(G134), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n455), .B1(new_n448), .B2(new_n449), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n439), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n333), .ZN(new_n473));
  INV_X1    g287(.A(G478), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(KEYINPUT15), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n473), .B(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT88), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n299), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n296), .A2(new_n298), .A3(KEYINPUT88), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(KEYINPUT19), .A3(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n481), .B(new_n206), .C1(KEYINPUT19), .C2(new_n299), .ZN(new_n482));
  INV_X1    g296(.A(G237), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(new_n428), .A3(G214), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n485), .A3(new_n208), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n252), .B(G214), .C1(KEYINPUT87), .C2(G143), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(G131), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n486), .A2(new_n200), .A3(new_n487), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n482), .A2(new_n302), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(KEYINPUT18), .A2(G131), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n488), .B(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n479), .A2(G146), .A3(new_n480), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n322), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(G113), .B(G122), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(new_n360), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n492), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G475), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n333), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(KEYINPUT89), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n488), .A2(KEYINPUT17), .A3(G131), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n505), .A2(new_n301), .A3(new_n302), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT17), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n489), .A2(new_n507), .A3(new_n490), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n506), .A2(new_n508), .B1(new_n494), .B2(new_n496), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n501), .B(new_n504), .C1(new_n509), .C2(new_n500), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT20), .ZN(new_n511));
  INV_X1    g325(.A(new_n508), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n505), .A2(new_n301), .A3(new_n302), .ZN(new_n513));
  INV_X1    g327(.A(new_n493), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n488), .B(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n496), .ZN(new_n516));
  OAI22_X1  g330(.A1(new_n512), .A2(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n499), .B1(new_n494), .B2(new_n496), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n517), .A2(new_n499), .B1(new_n518), .B2(new_n492), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT20), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n520), .A3(new_n504), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n511), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT91), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n499), .A2(KEYINPUT90), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n509), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n333), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n509), .A2(new_n524), .ZN(new_n527));
  OAI21_X1  g341(.A(G475), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n522), .A2(new_n523), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n523), .B1(new_n522), .B2(new_n528), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n436), .B(new_n477), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT95), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n510), .A2(KEYINPUT20), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n520), .B1(new_n519), .B2(new_n504), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n528), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT91), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n522), .A2(new_n523), .A3(new_n528), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n539), .A2(KEYINPUT95), .A3(new_n436), .A4(new_n477), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n426), .B1(new_n533), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT83), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT82), .ZN(new_n543));
  XNOR2_X1  g357(.A(G110), .B(G140), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n428), .A2(G227), .ZN(new_n545));
  XOR2_X1   g359(.A(new_n544), .B(new_n545), .Z(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT81), .B1(new_n376), .B2(new_n221), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n215), .A2(new_n217), .A3(new_n209), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n549), .B1(new_n218), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n220), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n376), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n369), .A2(new_n375), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT81), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n554), .A2(new_n555), .A3(new_n220), .A4(new_n214), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n548), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n233), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT12), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n557), .A2(KEYINPUT12), .A3(new_n233), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT10), .ZN(new_n563));
  AND4_X1   g377(.A1(new_n215), .A2(new_n217), .A3(new_n209), .A4(new_n219), .ZN(new_n564));
  OR2_X1    g378(.A1(new_n550), .A2(new_n218), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n564), .B1(new_n565), .B2(new_n549), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n563), .B1(new_n566), .B2(new_n554), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n390), .A2(new_n241), .A3(new_n393), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n233), .A2(KEYINPUT80), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT80), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n232), .A2(new_n571), .A3(new_n205), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT79), .ZN(new_n574));
  INV_X1    g388(.A(new_n221), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n369), .A2(KEYINPUT10), .A3(new_n375), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n376), .A2(KEYINPUT79), .A3(new_n221), .A4(KEYINPUT10), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n569), .A2(new_n573), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n547), .B1(new_n562), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n569), .A2(new_n573), .A3(new_n579), .ZN(new_n582));
  INV_X1    g396(.A(new_n233), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n569), .B2(new_n579), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n582), .A2(new_n584), .A3(new_n546), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n543), .B1(new_n581), .B2(new_n585), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n557), .A2(KEYINPUT12), .A3(new_n233), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT12), .B1(new_n557), .B2(new_n233), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n580), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n546), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n569), .A2(new_n579), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n580), .B(new_n547), .C1(new_n591), .C2(new_n583), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n590), .A2(KEYINPUT82), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n586), .A2(G469), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(G469), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(new_n333), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n546), .B1(new_n582), .B2(new_n584), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n580), .B(new_n547), .C1(new_n587), .C2(new_n588), .ZN(new_n598));
  AOI21_X1  g412(.A(G902), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n596), .B1(new_n599), .B2(new_n595), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n325), .B1(new_n438), .B2(new_n333), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n542), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  AOI211_X1 g418(.A(KEYINPUT83), .B(new_n602), .C1(new_n594), .C2(new_n600), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n541), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n354), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(new_n365), .ZN(G3));
  NOR2_X1   g422(.A1(new_n604), .A2(new_n605), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n273), .A2(new_n333), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n610), .A2(G472), .B1(new_n274), .B2(new_n273), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n353), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(new_n613), .B(KEYINPUT96), .Z(new_n614));
  NAND2_X1  g428(.A1(G478), .A2(G902), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n615), .B1(new_n473), .B2(G478), .ZN(new_n616));
  OAI21_X1  g430(.A(KEYINPUT33), .B1(new_n440), .B2(KEYINPUT98), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n472), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n617), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n468), .A2(new_n471), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n474), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(new_n537), .A3(new_n538), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n426), .A2(KEYINPUT97), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT97), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n625), .B(new_n355), .C1(new_n424), .C2(new_n425), .ZN(new_n626));
  AOI211_X1 g440(.A(new_n435), .B(new_n623), .C1(new_n624), .C2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n614), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT99), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT34), .B(G104), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  INV_X1    g446(.A(new_n477), .ZN(new_n633));
  INV_X1    g447(.A(new_n536), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI211_X1 g449(.A(new_n435), .B(new_n635), .C1(new_n624), .C2(new_n626), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n614), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT35), .B(G107), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  INV_X1    g454(.A(new_n347), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n328), .A2(KEYINPUT36), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n335), .B(new_n642), .Z(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n345), .B1(new_n641), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n611), .A2(new_n645), .ZN(new_n646));
  OR2_X1    g460(.A1(new_n606), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT37), .B(G110), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G12));
  AOI21_X1  g463(.A(new_n350), .B1(new_n347), .B2(new_n643), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n273), .A2(new_n274), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(KEYINPUT32), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n273), .A2(new_n187), .A3(new_n274), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n285), .A2(new_n286), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n333), .B1(new_n655), .B2(KEYINPUT29), .ZN(new_n656));
  OAI21_X1  g470(.A(G472), .B1(new_n656), .B2(new_n284), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n650), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n601), .A2(new_n603), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(KEYINPUT83), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n601), .A2(new_n542), .A3(new_n603), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n624), .A2(new_n626), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n430), .B1(G900), .B2(new_n431), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n634), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n477), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n658), .A2(new_n662), .A3(new_n663), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  NOR2_X1   g482(.A1(new_n424), .A2(new_n425), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT38), .ZN(new_n670));
  INV_X1    g484(.A(new_n355), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n529), .A2(new_n530), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n633), .ZN(new_n673));
  NOR4_X1   g487(.A1(new_n670), .A2(new_n671), .A3(new_n645), .A4(new_n673), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n278), .A2(new_n280), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n333), .B1(new_n675), .B2(new_n256), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n251), .B1(new_n271), .B2(new_n191), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n256), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(G472), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT100), .B1(new_n654), .B2(new_n680), .ZN(new_n681));
  OAI211_X1 g495(.A(KEYINPUT100), .B(new_n680), .C1(new_n276), .C2(new_n275), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n674), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT101), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n664), .B(KEYINPUT39), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n687), .B1(new_n604), .B2(new_n605), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT40), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n674), .B(KEYINPUT101), .C1(new_n681), .C2(new_n683), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n686), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G143), .ZN(G45));
  INV_X1    g507(.A(new_n623), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n664), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n658), .A2(new_n662), .A3(new_n663), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G146), .ZN(G48));
  OR2_X1    g512(.A1(new_n599), .A2(new_n595), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n599), .A2(new_n595), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n699), .A2(new_n603), .A3(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n290), .A2(new_n627), .A3(new_n353), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT41), .B(G113), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  NAND4_X1  g519(.A1(new_n290), .A2(new_n636), .A3(new_n353), .A4(new_n702), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G116), .ZN(G18));
  AOI21_X1  g521(.A(new_n701), .B1(new_n533), .B2(new_n540), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n290), .A2(new_n663), .A3(new_n708), .A4(new_n645), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G119), .ZN(G21));
  AND2_X1   g524(.A1(new_n281), .A2(new_n282), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n258), .B(new_n272), .C1(new_n711), .C2(new_n256), .ZN(new_n712));
  AOI22_X1  g526(.A1(new_n712), .A2(new_n274), .B1(G472), .B2(new_n610), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n350), .A2(new_n351), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n673), .B1(new_n624), .B2(new_n626), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n701), .A2(new_n435), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n713), .A2(new_n714), .A3(new_n715), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G122), .ZN(G24));
  AOI21_X1  g532(.A(new_n701), .B1(new_n624), .B2(new_n626), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(new_n713), .A3(new_n645), .A4(new_n696), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G125), .ZN(G27));
  NAND3_X1  g535(.A1(new_n590), .A2(G469), .A3(new_n592), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n600), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n602), .A2(new_n671), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n723), .A2(new_n669), .A3(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n290), .A2(new_n353), .A3(new_n726), .A4(new_n696), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT42), .ZN(new_n728));
  INV_X1    g542(.A(new_n714), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n654), .B2(new_n657), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n725), .A2(new_n695), .A3(new_n728), .ZN(new_n731));
  AOI22_X1  g545(.A1(new_n727), .A2(new_n728), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(new_n200), .ZN(G33));
  NAND4_X1  g547(.A1(new_n290), .A2(new_n353), .A3(new_n726), .A4(new_n666), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT102), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n714), .A2(new_n291), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT75), .B1(new_n350), .B2(new_n351), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n738), .B1(new_n654), .B2(new_n657), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT102), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n739), .A2(new_n740), .A3(new_n666), .A4(new_n726), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n735), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  INV_X1    g557(.A(new_n700), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n586), .A2(new_n593), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n595), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n590), .A2(KEYINPUT45), .A3(new_n592), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT103), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n596), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT46), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n744), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n596), .B1(new_n747), .B2(new_n750), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT46), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n602), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n687), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n616), .A2(new_n621), .ZN(new_n760));
  OAI21_X1  g574(.A(KEYINPUT43), .B1(new_n672), .B2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n539), .A2(new_n762), .A3(new_n622), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n610), .A2(G472), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n651), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n764), .A2(new_n766), .A3(KEYINPUT44), .A4(new_n645), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT44), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n761), .A2(new_n763), .A3(new_n645), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n768), .B1(new_n769), .B2(new_n611), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n669), .A2(new_n355), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n767), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n759), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n223), .ZN(G39));
  INV_X1    g589(.A(KEYINPUT104), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT47), .ZN(new_n777));
  INV_X1    g591(.A(new_n757), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n700), .B1(new_n756), .B2(KEYINPUT46), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n603), .B(new_n777), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NOR4_X1   g594(.A1(new_n290), .A2(new_n353), .A3(new_n695), .A4(new_n771), .ZN(new_n781));
  XNOR2_X1  g595(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n780), .B(new_n781), .C1(new_n758), .C2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G140), .ZN(G42));
  NOR2_X1   g598(.A1(G952), .A2(G953), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT115), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n702), .A2(new_n772), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT112), .ZN(new_n788));
  INV_X1    g602(.A(new_n430), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n764), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n788), .A2(new_n730), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT113), .ZN(new_n792));
  NOR2_X1   g606(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n793));
  AND2_X1   g607(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n794));
  OR3_X1    g608(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n428), .A2(G952), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n713), .A2(new_n714), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n797), .A2(new_n790), .A3(new_n719), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n788), .A2(new_n353), .A3(new_n789), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n681), .A2(new_n683), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI211_X1 g615(.A(new_n796), .B(new_n798), .C1(new_n801), .C2(new_n694), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n795), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(new_n793), .B2(new_n792), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n797), .A2(new_n790), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n670), .A2(new_n702), .A3(new_n671), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT50), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n801), .A2(new_n539), .A3(new_n760), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n713), .A2(new_n645), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n788), .A2(new_n790), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n808), .B(new_n809), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n805), .A2(new_n771), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT111), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n780), .B1(new_n758), .B2(new_n782), .ZN(new_n816));
  INV_X1    g630(.A(new_n699), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n744), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n602), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n815), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  OR3_X1    g634(.A1(new_n812), .A2(new_n813), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n813), .B1(new_n812), .B2(new_n820), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n804), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n654), .A2(new_n680), .ZN(new_n824));
  AND4_X1   g638(.A1(new_n603), .A2(new_n650), .A3(new_n664), .A4(new_n723), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n824), .A2(new_n715), .A3(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n667), .A2(new_n697), .A3(new_n720), .A4(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT109), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n667), .A2(new_n720), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n832), .A2(KEYINPUT52), .A3(new_n697), .A4(new_n826), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT109), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n827), .A2(new_n828), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n606), .B1(new_n354), .B2(new_n646), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n426), .A2(new_n435), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n672), .A2(new_n760), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n839), .B(new_n840), .C1(new_n633), .C2(new_n672), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n609), .A2(new_n612), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n838), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n810), .A2(new_n695), .A3(new_n725), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n735), .B2(new_n741), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n290), .A2(new_n645), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n771), .A2(new_n633), .A3(new_n665), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n848), .B1(new_n604), .B2(new_n605), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT108), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT108), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n658), .A2(new_n662), .A3(new_n851), .A4(new_n848), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n844), .A2(new_n846), .A3(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n706), .A2(new_n703), .A3(new_n709), .A4(new_n717), .ZN(new_n855));
  OR3_X1    g669(.A1(new_n855), .A2(new_n732), .A3(KEYINPUT110), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT110), .B1(new_n855), .B2(new_n732), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n854), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n833), .A2(new_n835), .ZN(new_n859));
  INV_X1    g673(.A(new_n841), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n662), .A2(new_n353), .A3(new_n611), .A4(new_n860), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n647), .B(new_n861), .C1(new_n354), .C2(new_n606), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n706), .A2(new_n709), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n703), .A2(new_n717), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT107), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n855), .A2(KEYINPUT107), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n862), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n732), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n846), .A2(new_n869), .A3(new_n853), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n859), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n837), .A2(new_n858), .B1(new_n871), .B2(new_n843), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n837), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n868), .A2(new_n870), .A3(new_n843), .ZN(new_n876));
  INV_X1    g690(.A(new_n871), .ZN(new_n877));
  OAI22_X1  g691(.A1(new_n875), .A2(new_n876), .B1(new_n877), .B2(new_n843), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n874), .B1(new_n878), .B2(new_n873), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n786), .B1(new_n823), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n714), .A2(new_n724), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT105), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n672), .A2(new_n760), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT49), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n882), .B(new_n883), .C1(new_n884), .C2(new_n818), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT106), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n818), .A2(new_n884), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n886), .A2(new_n800), .A3(new_n670), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n880), .A2(new_n888), .ZN(G75));
  NOR2_X1   g703(.A1(new_n428), .A2(G952), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n834), .B1(new_n833), .B2(new_n835), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n858), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n868), .A2(new_n870), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n827), .B(KEYINPUT52), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n843), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n333), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT56), .B1(new_n898), .B2(G210), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n416), .A2(new_n421), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n419), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT55), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n891), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n899), .A2(new_n902), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT116), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n899), .A2(KEYINPUT116), .A3(new_n902), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(G51));
  NAND2_X1  g722(.A1(new_n597), .A2(new_n598), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n894), .A2(new_n897), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(new_n873), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n596), .B(KEYINPUT57), .Z(new_n912));
  OAI21_X1  g726(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n898), .A2(new_n750), .A3(new_n747), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n890), .B1(new_n913), .B2(new_n914), .ZN(G54));
  AND3_X1   g729(.A1(new_n898), .A2(KEYINPUT58), .A3(G475), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n891), .B1(new_n916), .B2(new_n519), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n917), .B1(new_n519), .B2(new_n916), .ZN(G60));
  AND2_X1   g732(.A1(new_n618), .A2(new_n620), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n615), .B(KEYINPUT59), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n891), .B1(new_n911), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n919), .B1(new_n879), .B2(new_n920), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(G63));
  INV_X1    g738(.A(KEYINPUT121), .ZN(new_n925));
  NAND2_X1  g739(.A1(G217), .A2(G902), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT118), .ZN(new_n927));
  XNOR2_X1  g741(.A(KEYINPUT117), .B(KEYINPUT60), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n927), .B(new_n928), .Z(new_n929));
  NAND3_X1  g743(.A1(new_n910), .A2(new_n643), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT61), .ZN(new_n931));
  INV_X1    g745(.A(new_n929), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n894), .B2(new_n897), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n332), .B(KEYINPUT120), .Z(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n891), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n925), .B1(new_n931), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n933), .B2(new_n643), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n934), .B1(new_n872), .B2(new_n932), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n939), .A2(KEYINPUT121), .A3(new_n891), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  AOI211_X1 g756(.A(new_n644), .B(new_n932), .C1(new_n894), .C2(new_n897), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT119), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n940), .B(new_n891), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n930), .A2(KEYINPUT119), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n938), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n942), .A2(new_n947), .ZN(G66));
  OAI21_X1  g762(.A(G953), .B1(new_n433), .B2(new_n404), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n868), .B2(G953), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n900), .B1(G898), .B2(new_n428), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(G69));
  INV_X1    g766(.A(KEYINPUT122), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n667), .A2(new_n697), .A3(new_n720), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n692), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n953), .B1(new_n955), .B2(KEYINPUT62), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(KEYINPUT62), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT62), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n692), .A2(KEYINPUT122), .A3(new_n958), .A4(new_n954), .ZN(new_n959));
  INV_X1    g773(.A(new_n783), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n840), .B1(new_n633), .B2(new_n672), .ZN(new_n961));
  OR4_X1    g775(.A1(new_n354), .A2(new_n688), .A3(new_n771), .A4(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n759), .B2(new_n773), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n956), .A2(new_n957), .A3(new_n959), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n428), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n481), .B1(KEYINPUT19), .B2(new_n299), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n271), .B(new_n967), .Z(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n954), .A2(new_n869), .A3(new_n742), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT124), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n730), .A2(new_n715), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n773), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n973), .A2(new_n687), .A3(new_n758), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n970), .A2(new_n971), .A3(new_n783), .A4(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n732), .B1(new_n741), .B2(new_n735), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n976), .A2(new_n783), .A3(new_n954), .A4(new_n974), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(KEYINPUT124), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n975), .A2(new_n978), .A3(new_n428), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n968), .B1(G900), .B2(G953), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n428), .B1(G227), .B2(G900), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT123), .Z(new_n983));
  NAND3_X1  g797(.A1(new_n969), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT125), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n979), .A2(KEYINPUT125), .A3(new_n980), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n986), .A2(new_n969), .A3(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT126), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n988), .A2(new_n989), .A3(new_n982), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n989), .B1(new_n988), .B2(new_n982), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n984), .B1(new_n990), .B2(new_n991), .ZN(G72));
  NAND2_X1  g806(.A1(G472), .A2(G902), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT63), .Z(new_n994));
  INV_X1    g808(.A(new_n868), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n994), .B1(new_n965), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n679), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT127), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n678), .A2(new_n286), .A3(new_n994), .ZN(new_n999));
  INV_X1    g813(.A(new_n994), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n975), .A2(new_n978), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1000), .B1(new_n1001), .B2(new_n868), .ZN(new_n1002));
  OAI221_X1 g816(.A(new_n891), .B1(new_n878), .B2(new_n999), .C1(new_n1002), .C2(new_n286), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n998), .A2(new_n1003), .ZN(G57));
endmodule


