//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT3), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(KEYINPUT83), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT83), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(KEYINPUT3), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  OAI22_X1  g006(.A1(new_n189), .A2(new_n191), .B1(new_n192), .B2(G107), .ZN(new_n193));
  INV_X1    g007(.A(G101), .ZN(new_n194));
  INV_X1    g008(.A(G107), .ZN(new_n195));
  OAI211_X1 g009(.A(G104), .B(new_n195), .C1(new_n188), .C2(KEYINPUT83), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(G104), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n193), .A2(new_n194), .A3(new_n196), .A4(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n192), .A2(G107), .ZN(new_n200));
  OAI21_X1  g014(.A(G101), .B1(new_n200), .B2(new_n197), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT2), .B(G113), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n205));
  XNOR2_X1  g019(.A(G116), .B(G119), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G119), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G116), .ZN(new_n209));
  INV_X1    g023(.A(G116), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G119), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT66), .B1(new_n212), .B2(new_n203), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n207), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n209), .A2(new_n211), .A3(KEYINPUT5), .ZN(new_n215));
  OR3_X1    g029(.A1(new_n210), .A2(KEYINPUT5), .A3(G119), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(G113), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n202), .A2(new_n218), .ZN(new_n219));
  XOR2_X1   g033(.A(G110), .B(G122), .Z(new_n220));
  XOR2_X1   g034(.A(new_n220), .B(KEYINPUT8), .Z(new_n221));
  INV_X1    g035(.A(KEYINPUT85), .ZN(new_n222));
  INV_X1    g036(.A(G113), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n223), .B1(new_n206), .B2(KEYINPUT5), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n222), .B1(new_n224), .B2(new_n216), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n215), .A2(new_n216), .A3(new_n222), .A4(G113), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n214), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n219), .B(new_n221), .C1(new_n202), .C2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G143), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G146), .ZN(new_n231));
  INV_X1    g045(.A(G146), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G143), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n231), .A2(new_n233), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  XOR2_X1   g051(.A(KEYINPUT0), .B(G128), .Z(new_n238));
  OAI21_X1  g052(.A(new_n235), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G128), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n230), .B(G146), .C1(new_n240), .C2(KEYINPUT1), .ZN(new_n241));
  OR2_X1    g055(.A1(new_n240), .A2(KEYINPUT1), .ZN(new_n242));
  OAI221_X1 g056(.A(new_n241), .B1(G128), .B2(new_n233), .C1(new_n236), .C2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G125), .ZN(new_n244));
  MUX2_X1   g058(.A(new_n239), .B(new_n243), .S(new_n244), .Z(new_n245));
  INV_X1    g059(.A(G953), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G224), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT7), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n245), .B(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n199), .A2(new_n201), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT86), .B1(new_n228), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n220), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n212), .A2(new_n203), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n214), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT83), .B(KEYINPUT3), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n196), .B(new_n198), .C1(new_n255), .C2(new_n200), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G101), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT4), .A3(new_n199), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n256), .A2(new_n259), .A3(G101), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n254), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n217), .A2(KEYINPUT85), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n262), .A2(new_n226), .B1(new_n207), .B2(new_n213), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT86), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n202), .A3(new_n264), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n251), .A2(new_n252), .A3(new_n261), .A4(new_n265), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n266), .A2(KEYINPUT87), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(KEYINPUT87), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n229), .B(new_n249), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n265), .A2(new_n261), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n252), .B1(new_n270), .B2(new_n251), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(KEYINPUT6), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n251), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n220), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n274), .B1(new_n267), .B2(new_n268), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n272), .B1(new_n275), .B2(KEYINPUT6), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n245), .B(new_n247), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n187), .B(new_n269), .C1(new_n276), .C2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(G210), .B1(G237), .B2(G902), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n274), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT87), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n270), .A2(new_n285), .A3(new_n252), .A4(new_n251), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n266), .A2(KEYINPUT87), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n271), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n284), .B1(new_n288), .B2(new_n283), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n277), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n290), .A2(new_n187), .A3(new_n280), .A4(new_n269), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n282), .A2(KEYINPUT88), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(G902), .B1(new_n289), .B2(new_n277), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n280), .B1(new_n293), .B2(new_n269), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT88), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n202), .A2(KEYINPUT10), .A3(new_n243), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n258), .A2(new_n239), .A3(new_n260), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n199), .A2(new_n243), .A3(new_n201), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT10), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n298), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT11), .ZN(new_n304));
  INV_X1    g118(.A(G134), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n304), .B1(new_n305), .B2(G137), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(G137), .ZN(new_n307));
  INV_X1    g121(.A(G137), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(KEYINPUT11), .A3(G134), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G131), .ZN(new_n311));
  INV_X1    g125(.A(G131), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT64), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT64), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G131), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n316), .A2(new_n307), .A3(new_n309), .A4(new_n306), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n303), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n318), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n298), .A2(new_n299), .A3(new_n320), .A4(new_n302), .ZN(new_n321));
  XNOR2_X1  g135(.A(G110), .B(G140), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(KEYINPUT82), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n246), .A2(G227), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n323), .B(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n319), .A2(new_n321), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n321), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n243), .B1(new_n199), .B2(new_n201), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT84), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n328), .B1(new_n329), .B2(new_n300), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n202), .A2(KEYINPUT84), .A3(new_n243), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n318), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT12), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g148(.A(KEYINPUT12), .B(new_n318), .C1(new_n330), .C2(new_n331), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n327), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OAI211_X1 g150(.A(G469), .B(new_n326), .C1(new_n336), .C2(new_n325), .ZN(new_n337));
  INV_X1    g151(.A(G469), .ZN(new_n338));
  XOR2_X1   g152(.A(KEYINPUT71), .B(G902), .Z(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n321), .A2(new_n325), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n341), .B1(new_n334), .B2(new_n335), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n325), .B1(new_n319), .B2(new_n321), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n338), .B(new_n340), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(G469), .A2(G902), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n337), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G221), .ZN(new_n347));
  XOR2_X1   g161(.A(KEYINPUT9), .B(G234), .Z(new_n348));
  AOI21_X1  g162(.A(new_n347), .B1(new_n348), .B2(new_n187), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(G214), .B1(G237), .B2(G902), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n297), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT74), .B(G140), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT75), .B1(new_n355), .B2(new_n244), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n244), .A2(G140), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT75), .ZN(new_n358));
  INV_X1    g172(.A(G140), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n359), .A2(KEYINPUT74), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n359), .A2(KEYINPUT74), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n358), .B(G125), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n356), .A2(new_n357), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT16), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT16), .B1(new_n359), .B2(G125), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n232), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT76), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n364), .A2(new_n366), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G146), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n364), .A2(KEYINPUT76), .A3(new_n232), .A4(new_n366), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n369), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  XOR2_X1   g187(.A(KEYINPUT24), .B(G110), .Z(new_n374));
  XNOR2_X1  g188(.A(G119), .B(G128), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n208), .A2(KEYINPUT23), .A3(G128), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n377), .B1(new_n375), .B2(KEYINPUT23), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G110), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n373), .A2(new_n376), .A3(new_n379), .ZN(new_n380));
  OAI22_X1  g194(.A1(new_n378), .A2(G110), .B1(new_n375), .B2(new_n374), .ZN(new_n381));
  XNOR2_X1  g195(.A(G125), .B(G140), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(KEYINPUT77), .ZN(new_n383));
  OR2_X1    g197(.A1(new_n383), .A2(G146), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n371), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT78), .B(KEYINPUT22), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n387), .B(G137), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n246), .A2(G221), .A3(G234), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n388), .B(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(KEYINPUT79), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n380), .A2(new_n390), .A3(new_n385), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n340), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT80), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(KEYINPUT25), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(KEYINPUT73), .B(G217), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n400), .B1(new_n340), .B2(G234), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n392), .A2(new_n340), .A3(new_n396), .A4(new_n393), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n398), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT81), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n398), .A2(KEYINPUT81), .A3(new_n401), .A4(new_n402), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n392), .A2(new_n393), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n401), .A2(G902), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n405), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n308), .A2(G134), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n307), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G131), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT65), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT65), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n415), .A3(G131), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n243), .A2(new_n317), .A3(new_n414), .A4(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT67), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n318), .A2(new_n418), .A3(new_n239), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n418), .B1(new_n318), .B2(new_n239), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n417), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n254), .ZN(new_n422));
  INV_X1    g236(.A(new_n254), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n423), .B(new_n417), .C1(new_n419), .C2(new_n420), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n422), .A2(KEYINPUT69), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT69), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n421), .A2(new_n426), .A3(new_n254), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(KEYINPUT28), .A3(new_n427), .ZN(new_n428));
  XOR2_X1   g242(.A(KEYINPUT26), .B(G101), .Z(new_n429));
  INV_X1    g243(.A(G237), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(new_n246), .A3(G210), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n429), .B(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n432), .B(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  OR2_X1    g249(.A1(new_n419), .A2(new_n420), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n436), .A2(KEYINPUT28), .A3(new_n423), .A4(new_n417), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT29), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n318), .A2(new_n239), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n417), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n254), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT28), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(new_n440), .B2(new_n254), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n437), .A2(new_n438), .A3(new_n441), .A4(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n443), .B(KEYINPUT70), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n428), .A2(new_n435), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n340), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n435), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n440), .A2(KEYINPUT30), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n449), .B1(KEYINPUT30), .B2(new_n421), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n434), .B(new_n424), .C1(new_n450), .C2(new_n423), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT29), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(G472), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT72), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g269(.A(KEYINPUT72), .B(G472), .C1(new_n447), .C2(new_n452), .ZN(new_n456));
  INV_X1    g270(.A(new_n424), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n421), .A2(KEYINPUT30), .ZN(new_n458));
  INV_X1    g272(.A(new_n449), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n457), .B1(new_n460), .B2(new_n254), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT31), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n462), .A3(new_n435), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n435), .B(new_n424), .C1(new_n450), .C2(new_n423), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT31), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n437), .A2(new_n441), .A3(new_n443), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n434), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n463), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(G472), .A2(G902), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT32), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT32), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n468), .A2(new_n472), .A3(new_n469), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n455), .A2(new_n456), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n410), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(G475), .A2(G902), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT17), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n430), .A2(new_n246), .A3(G214), .ZN(new_n478));
  OR2_X1    g292(.A1(new_n478), .A2(new_n230), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n230), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n479), .A2(new_n316), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n316), .B1(new_n479), .B2(new_n480), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n477), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OR2_X1    g297(.A1(new_n482), .A2(new_n477), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n369), .A2(new_n371), .A3(new_n485), .A4(new_n372), .ZN(new_n486));
  XNOR2_X1  g300(.A(G113), .B(G122), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(new_n192), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n478), .B(new_n230), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT89), .ZN(new_n490));
  AND2_X1   g304(.A1(KEYINPUT18), .A2(G131), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n363), .A2(G146), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n384), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n492), .B(new_n494), .C1(KEYINPUT89), .C2(new_n489), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n486), .A2(new_n488), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT91), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT91), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n486), .A2(new_n498), .A3(new_n495), .A4(new_n488), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n363), .A2(KEYINPUT19), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n501), .B(new_n232), .C1(KEYINPUT19), .C2(new_n383), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n371), .A2(KEYINPUT90), .A3(new_n502), .ZN(new_n503));
  OR2_X1    g317(.A1(new_n481), .A2(new_n482), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT90), .B1(new_n371), .B2(new_n502), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n495), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n488), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n500), .A2(KEYINPUT92), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(KEYINPUT92), .B1(new_n500), .B2(new_n509), .ZN(new_n511));
  OAI211_X1 g325(.A(KEYINPUT20), .B(new_n476), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n488), .B1(new_n486), .B2(new_n495), .ZN(new_n513));
  OR2_X1    g327(.A1(new_n513), .A2(KEYINPUT93), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(KEYINPUT93), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n500), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(G475), .B1(new_n516), .B2(G902), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n500), .A2(new_n509), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n476), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT20), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g336(.A1(KEYINPUT94), .A2(G122), .ZN(new_n523));
  NOR2_X1   g337(.A1(KEYINPUT94), .A2(G122), .ZN(new_n524));
  OAI21_X1  g338(.A(G116), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n195), .B1(new_n525), .B2(KEYINPUT14), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n210), .A2(G122), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  XOR2_X1   g342(.A(new_n526), .B(new_n528), .Z(new_n529));
  XNOR2_X1  g343(.A(G128), .B(G143), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(new_n305), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n528), .A2(G107), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n195), .B1(new_n525), .B2(new_n527), .ZN(new_n534));
  OR2_X1    g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n530), .A2(KEYINPUT13), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n240), .A2(KEYINPUT13), .A3(G143), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(new_n305), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n536), .A2(new_n538), .B1(new_n305), .B2(new_n530), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT95), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n539), .B(KEYINPUT95), .C1(new_n533), .C2(new_n534), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n532), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n348), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n544), .A2(G953), .A3(new_n400), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n532), .B(new_n545), .C1(new_n540), .C2(new_n542), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(KEYINPUT96), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT96), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n543), .A2(new_n550), .A3(new_n546), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(G478), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(KEYINPUT15), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n552), .A2(new_n340), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n549), .A2(new_n340), .A3(new_n551), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n554), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n246), .A2(G952), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n560), .B1(G234), .B2(G237), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  AOI211_X1 g376(.A(new_n246), .B(new_n340), .C1(G234), .C2(G237), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT21), .B(G898), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(KEYINPUT97), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n562), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n559), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n518), .A2(KEYINPUT98), .A3(new_n522), .A4(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT98), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n512), .A2(new_n517), .A3(new_n522), .ZN(new_n572));
  INV_X1    g386(.A(new_n559), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n567), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n571), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n354), .A2(new_n475), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(G101), .ZN(G3));
  AOI21_X1  g392(.A(new_n353), .B1(new_n282), .B2(new_n291), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n567), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n557), .A2(new_n553), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT33), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n552), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n547), .A2(KEYINPUT33), .A3(new_n548), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n340), .A2(G478), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n581), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n572), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n580), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n468), .A2(new_n340), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(G472), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n470), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n410), .A2(new_n351), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT34), .B(G104), .Z(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(G6));
  INV_X1    g410(.A(KEYINPUT99), .ZN(new_n597));
  INV_X1    g411(.A(new_n291), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n352), .B1(new_n598), .B2(new_n294), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(new_n568), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n476), .B1(new_n510), .B2(new_n511), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n521), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n602), .A2(new_n517), .A3(new_n512), .A4(new_n559), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n597), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n580), .A2(new_n603), .A3(KEYINPUT99), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n593), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT35), .B(G107), .Z(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G9));
  INV_X1    g423(.A(new_n592), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n391), .A2(KEYINPUT36), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n386), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n408), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n405), .A2(new_n406), .A3(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n354), .A2(new_n576), .A3(new_n610), .A4(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT37), .ZN(new_n616));
  XOR2_X1   g430(.A(new_n616), .B(G110), .Z(G12));
  INV_X1    g431(.A(G900), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n561), .B1(new_n563), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n604), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n455), .A2(new_n456), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n471), .A2(new_n473), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n351), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n624), .A2(new_n614), .A3(new_n579), .A4(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(new_n240), .ZN(G30));
  XNOR2_X1  g442(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n297), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n572), .A2(new_n559), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n425), .A2(new_n427), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n187), .B1(new_n632), .B2(new_n435), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n461), .A2(new_n434), .ZN(new_n634));
  OAI21_X1  g448(.A(G472), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n631), .B1(new_n623), .B2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n619), .B(KEYINPUT39), .Z(new_n637));
  NAND2_X1  g451(.A1(new_n625), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n638), .B(KEYINPUT40), .Z(new_n639));
  NAND3_X1  g453(.A1(new_n630), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT101), .ZN(new_n641));
  INV_X1    g455(.A(new_n614), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n352), .ZN(new_n643));
  OR3_X1    g457(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n641), .B1(new_n640), .B2(new_n643), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(new_n230), .ZN(G45));
  NAND3_X1  g461(.A1(new_n572), .A2(new_n587), .A3(new_n620), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n626), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(new_n232), .ZN(G48));
  OAI21_X1  g464(.A(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(G469), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n344), .A2(KEYINPUT102), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n652), .A2(KEYINPUT102), .A3(new_n344), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n350), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n410), .A2(new_n658), .A3(new_n474), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n589), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT41), .B(G113), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G15));
  AOI21_X1  g476(.A(new_n349), .B1(new_n655), .B2(new_n656), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n475), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n600), .A2(new_n604), .A3(new_n597), .ZN(new_n665));
  OAI21_X1  g479(.A(KEYINPUT99), .B1(new_n580), .B2(new_n603), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n210), .ZN(G18));
  NOR2_X1   g482(.A1(new_n642), .A2(new_n474), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n579), .A2(new_n663), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n576), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G119), .ZN(G21));
  NOR2_X1   g487(.A1(new_n670), .A2(new_n631), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n469), .B(KEYINPUT103), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n463), .A2(new_n465), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n435), .B1(new_n428), .B2(new_n445), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT104), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n680), .B(new_n675), .C1(new_n676), .C2(new_n677), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n679), .A2(new_n591), .A3(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n410), .A2(new_n682), .A3(new_n568), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n674), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G122), .ZN(G24));
  AND3_X1   g499(.A1(new_n679), .A2(new_n591), .A3(new_n681), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n614), .A2(new_n579), .A3(new_n663), .A4(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n648), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n572), .A2(new_n587), .A3(KEYINPUT105), .A4(new_n620), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n687), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n244), .ZN(G27));
  AND2_X1   g506(.A1(new_n689), .A2(new_n690), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n353), .B1(new_n292), .B2(new_n296), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n346), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n346), .A2(new_n695), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n349), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n475), .A2(new_n694), .A3(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n693), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n475), .A2(new_n694), .A3(new_n698), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n689), .A2(new_n690), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT42), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n312), .ZN(G33));
  NOR2_X1   g520(.A1(new_n699), .A2(new_n621), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n305), .ZN(G36));
  INV_X1    g522(.A(KEYINPUT46), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n326), .B1(new_n336), .B2(new_n325), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT45), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n709), .B(G469), .C1(new_n711), .C2(G902), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n712), .A2(KEYINPUT107), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(G469), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(KEYINPUT46), .A3(new_n345), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n712), .A2(KEYINPUT107), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n713), .A2(new_n344), .A3(new_n715), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n350), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n719), .A2(new_n637), .ZN(new_n720));
  INV_X1    g534(.A(new_n694), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n614), .A2(new_n592), .ZN(new_n722));
  INV_X1    g536(.A(new_n572), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT43), .B1(new_n723), .B2(KEYINPUT108), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n587), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n724), .A2(new_n725), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n722), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n721), .B1(new_n729), .B2(KEYINPUT44), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n720), .B(new_n730), .C1(KEYINPUT44), .C2(new_n729), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G137), .ZN(G39));
  INV_X1    g546(.A(KEYINPUT109), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(KEYINPUT47), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n733), .A2(KEYINPUT47), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n719), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n648), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n718), .B1(new_n733), .B2(KEYINPUT47), .ZN(new_n738));
  INV_X1    g552(.A(new_n410), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n721), .A2(new_n739), .A3(new_n624), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n736), .A2(new_n737), .A3(new_n738), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G140), .ZN(G42));
  AOI21_X1  g556(.A(new_n562), .B1(new_n727), .B2(new_n728), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n410), .A2(new_n682), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n630), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n745), .A2(new_n353), .A3(new_n746), .A4(new_n663), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n721), .A2(new_n658), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n743), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT114), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n614), .A2(new_n686), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n736), .A2(new_n738), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n350), .B1(new_n655), .B2(new_n656), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n694), .B(new_n745), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n750), .A2(new_n739), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n623), .A2(new_n635), .ZN(new_n761));
  OR3_X1    g575(.A1(new_n760), .A2(new_n562), .A3(new_n761), .ZN(new_n762));
  OR3_X1    g576(.A1(new_n762), .A2(new_n572), .A3(new_n587), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n749), .A2(new_n756), .A3(new_n759), .A4(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT51), .ZN(new_n765));
  INV_X1    g579(.A(new_n707), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n698), .A2(new_n686), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n767), .B1(new_n689), .B2(new_n690), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n559), .B1(new_n601), .B2(new_n521), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n624), .A2(new_n625), .A3(new_n620), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n512), .A2(new_n517), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n614), .B(new_n694), .C1(new_n768), .C2(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n766), .B(new_n773), .C1(new_n701), .C2(new_n704), .ZN(new_n774));
  INV_X1    g588(.A(new_n626), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n603), .A2(new_n619), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n775), .B1(new_n776), .B2(new_n737), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n696), .A2(new_n697), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n350), .ZN(new_n779));
  AND4_X1   g593(.A1(new_n405), .A2(new_n406), .A3(new_n613), .A4(new_n620), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n779), .B1(new_n780), .B2(KEYINPUT113), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n631), .A2(new_n599), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n783), .B1(new_n614), .B2(new_n619), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n781), .A2(new_n761), .A3(new_n782), .A4(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n703), .A2(new_n671), .A3(new_n755), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n777), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n626), .B1(new_n621), .B2(new_n648), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n691), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(KEYINPUT52), .A3(new_n785), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n774), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n297), .A2(new_n353), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n588), .B1(new_n572), .B2(new_n573), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n794), .A2(new_n593), .A3(new_n795), .A4(new_n567), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n615), .A2(new_n577), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n672), .A2(new_n660), .A3(new_n684), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT111), .B1(new_n798), .B2(new_n667), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n659), .B1(new_n605), .B2(new_n606), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n589), .A2(new_n659), .B1(new_n674), .B2(new_n683), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT111), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n800), .A2(new_n801), .A3(new_n802), .A4(new_n672), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n797), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n793), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n789), .A2(new_n792), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT53), .B1(new_n806), .B2(KEYINPUT112), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n805), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT54), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n810));
  INV_X1    g624(.A(new_n774), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n806), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n799), .A2(new_n803), .ZN(new_n813));
  INV_X1    g627(.A(new_n797), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n810), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n798), .A2(new_n667), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n797), .A2(new_n810), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n793), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n816), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n762), .A2(new_n588), .ZN(new_n822));
  AOI211_X1 g636(.A(new_n560), .B(new_n822), .C1(new_n745), .C2(new_n671), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n765), .A2(new_n809), .A3(new_n821), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n753), .A2(new_n475), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(KEYINPUT48), .ZN(new_n827));
  XOR2_X1   g641(.A(new_n825), .B(new_n827), .Z(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(new_n826), .B2(KEYINPUT48), .ZN(new_n829));
  OAI22_X1  g643(.A1(new_n824), .A2(new_n829), .B1(G952), .B2(G953), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT49), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n657), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n623), .A2(new_n350), .A3(new_n635), .ZN(new_n833));
  NOR4_X1   g647(.A1(new_n725), .A2(new_n353), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n746), .A2(new_n834), .A3(new_n739), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n831), .B2(new_n657), .ZN(new_n836));
  XOR2_X1   g650(.A(new_n836), .B(KEYINPUT110), .Z(new_n837));
  NAND2_X1  g651(.A1(new_n830), .A2(new_n837), .ZN(G75));
  AOI21_X1  g652(.A(new_n340), .B1(new_n816), .B2(new_n820), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT56), .B1(new_n839), .B2(new_n281), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n276), .A2(new_n278), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n290), .ZN(new_n842));
  XOR2_X1   g656(.A(new_n842), .B(KEYINPUT55), .Z(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(KEYINPUT116), .B2(KEYINPUT56), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n246), .A2(G952), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n840), .A2(new_n845), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n846), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT117), .ZN(G51));
  INV_X1    g665(.A(new_n714), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n839), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT119), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n839), .A2(new_n855), .A3(new_n852), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT53), .B1(new_n793), .B2(new_n804), .ZN(new_n859));
  AND4_X1   g673(.A1(new_n806), .A2(new_n811), .A3(new_n818), .A4(new_n819), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT54), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n821), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n345), .B(KEYINPUT57), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n858), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  AOI211_X1 g679(.A(KEYINPUT118), .B(new_n863), .C1(new_n861), .C2(new_n821), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n342), .A2(new_n343), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n857), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT120), .B1(new_n869), .B2(new_n847), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n862), .A2(new_n864), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT118), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n862), .A2(new_n858), .A3(new_n864), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(new_n868), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n857), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n877), .A3(new_n848), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n870), .A2(new_n878), .ZN(G54));
  NAND3_X1  g693(.A1(new_n839), .A2(KEYINPUT58), .A3(G475), .ZN(new_n880));
  OR2_X1    g694(.A1(new_n510), .A2(new_n511), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT121), .Z(new_n884));
  OAI21_X1  g698(.A(new_n848), .B1(new_n880), .B2(new_n882), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(G60));
  NAND2_X1  g700(.A1(G478), .A2(G902), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT59), .Z(new_n888));
  INV_X1    g702(.A(new_n585), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n862), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n888), .B1(new_n809), .B2(new_n821), .ZN(new_n891));
  OAI221_X1 g705(.A(new_n848), .B1(new_n888), .B2(new_n890), .C1(new_n891), .C2(new_n889), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(G63));
  NAND2_X1  g707(.A1(G217), .A2(G902), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT60), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n816), .B2(new_n820), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n848), .B1(new_n896), .B2(new_n407), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n612), .B2(new_n896), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT61), .ZN(G66));
  AOI21_X1  g713(.A(new_n246), .B1(new_n566), .B2(G224), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n804), .B(KEYINPUT122), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n900), .B1(new_n902), .B2(new_n246), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n276), .B1(G898), .B2(new_n246), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n903), .B(new_n904), .Z(G69));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n731), .A2(new_n741), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n908));
  INV_X1    g722(.A(new_n791), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n908), .B1(new_n646), .B2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n644), .A2(KEYINPUT62), .A3(new_n645), .A4(new_n791), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n907), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n475), .A2(new_n694), .ZN(new_n913));
  INV_X1    g727(.A(new_n638), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n914), .A3(new_n795), .ZN(new_n915));
  AOI21_X1  g729(.A(G953), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n501), .B1(KEYINPUT19), .B2(new_n383), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n460), .B(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n906), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n915), .ZN(new_n921));
  AOI211_X1 g735(.A(new_n921), .B(new_n907), .C1(new_n910), .C2(new_n911), .ZN(new_n922));
  OAI211_X1 g736(.A(KEYINPUT123), .B(new_n918), .C1(new_n922), .C2(G953), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n246), .B1(G227), .B2(G900), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n907), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n705), .A2(new_n707), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n720), .A2(new_n475), .A3(new_n782), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n928), .A2(new_n791), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n926), .A2(new_n246), .A3(new_n927), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(G900), .A2(G953), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n930), .A2(new_n919), .A3(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n920), .A2(new_n923), .A3(new_n925), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(KEYINPUT124), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT124), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n930), .A2(new_n935), .A3(new_n919), .A4(new_n931), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n920), .A2(new_n923), .A3(new_n934), .A4(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT125), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n937), .A2(new_n938), .A3(new_n924), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n938), .B1(new_n937), .B2(new_n924), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n933), .B1(new_n939), .B2(new_n940), .ZN(G72));
  NAND2_X1  g755(.A1(G472), .A2(G902), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT63), .Z(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT126), .Z(new_n944));
  NAND3_X1  g758(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n944), .B1(new_n945), .B2(new_n902), .ZN(new_n946));
  INV_X1    g760(.A(new_n451), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n847), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n808), .A2(new_n451), .A3(new_n943), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n948), .B1(new_n634), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n922), .A2(new_n901), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n944), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n950), .B1(new_n634), .B2(new_n952), .ZN(G57));
endmodule


