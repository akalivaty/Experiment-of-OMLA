//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 1 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 0 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988,
    new_n989;
  OAI21_X1  g000(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  INV_X1    g003(.A(G176gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT66), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n210));
  AOI22_X1  g009(.A1(new_n202), .A2(new_n206), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT25), .ZN(new_n212));
  NAND3_X1  g011(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND4_X1  g014(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OR3_X1    g016(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT24), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n218), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n211), .B(new_n212), .C1(new_n217), .C2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G183gat), .ZN(new_n225));
  INV_X1    g024(.A(G190gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT67), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(G183gat), .B2(G190gat), .ZN(new_n229));
  AND4_X1   g028(.A1(new_n221), .A2(new_n227), .A3(new_n229), .A4(new_n213), .ZN(new_n230));
  INV_X1    g029(.A(new_n202), .ZN(new_n231));
  NOR3_X1   g030(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n232));
  INV_X1    g031(.A(new_n210), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n234));
  OAI22_X1  g033(.A1(new_n231), .A2(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT25), .B1(new_n230), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n204), .A2(new_n205), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n237), .B1(new_n238), .B2(KEYINPUT26), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n209), .A2(new_n210), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(KEYINPUT26), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT26), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n242), .A2(new_n204), .A3(new_n205), .A4(KEYINPUT68), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n239), .A2(new_n240), .A3(new_n241), .A4(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(new_n219), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT27), .B(G183gat), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT28), .B1(new_n246), .B2(new_n226), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n225), .A2(KEYINPUT27), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT27), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(G183gat), .ZN(new_n250));
  AND4_X1   g049(.A1(KEYINPUT28), .A2(new_n248), .A3(new_n250), .A4(new_n226), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n224), .B(new_n236), .C1(new_n245), .C2(new_n252), .ZN(new_n253));
  OR2_X1    g052(.A1(G127gat), .A2(G134gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n255), .A2(new_n256), .B1(G127gat), .B2(G134gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(G113gat), .B(G120gat), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n254), .B(new_n257), .C1(new_n258), .C2(KEYINPUT1), .ZN(new_n259));
  INV_X1    g058(.A(G120gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G113gat), .ZN(new_n261));
  INV_X1    g060(.A(G113gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G120gat), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT1), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n255), .A2(new_n256), .ZN(new_n265));
  NAND2_X1  g064(.A1(G127gat), .A2(G134gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n254), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n259), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n259), .A2(new_n268), .A3(KEYINPUT70), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OR2_X1    g072(.A1(new_n253), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G227gat), .ZN(new_n275));
  INV_X1    g074(.A(G233gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n253), .A2(new_n273), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n274), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT34), .ZN(new_n281));
  XOR2_X1   g080(.A(G15gat), .B(G43gat), .Z(new_n282));
  XNOR2_X1  g081(.A(G71gat), .B(G99gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n278), .B1(new_n274), .B2(new_n279), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n284), .B1(new_n285), .B2(KEYINPUT33), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT32), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n286), .A2(new_n288), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n281), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n291), .ZN(new_n293));
  INV_X1    g092(.A(new_n281), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n293), .A2(new_n294), .A3(new_n289), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT71), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(KEYINPUT36), .ZN(new_n298));
  XNOR2_X1  g097(.A(G1gat), .B(G29gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(KEYINPUT0), .ZN(new_n300));
  XNOR2_X1  g099(.A(G57gat), .B(G85gat), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n300), .B(new_n301), .Z(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT2), .ZN(new_n307));
  NAND2_X1  g106(.A1(G141gat), .A2(G148gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT79), .ZN(new_n310));
  INV_X1    g109(.A(G155gat), .ZN(new_n311));
  INV_X1    g110(.A(G162gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n310), .B1(new_n313), .B2(new_n306), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n310), .A3(new_n306), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT78), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n307), .A2(new_n317), .ZN(new_n318));
  AND2_X1   g117(.A1(G141gat), .A2(G148gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n319), .A2(new_n304), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n306), .A2(KEYINPUT78), .A3(KEYINPUT2), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n318), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n306), .ZN(new_n323));
  NOR2_X1   g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n315), .A2(new_n316), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(new_n269), .ZN(new_n327));
  NAND2_X1  g126(.A1(G225gat), .A2(G233gat), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT5), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n314), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n330), .A2(new_n307), .A3(new_n320), .A4(new_n316), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n322), .A2(new_n325), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n333), .A2(KEYINPUT4), .A3(new_n269), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT80), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT80), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n271), .A2(new_n326), .A3(new_n272), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n336), .B1(new_n337), .B2(KEYINPUT4), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n335), .B1(new_n338), .B2(new_n334), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n333), .A2(KEYINPUT3), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n342), .A3(new_n269), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n343), .A2(new_n328), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT81), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT81), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n339), .A2(new_n347), .A3(new_n344), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n329), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT4), .B1(new_n333), .B2(new_n269), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n350), .B1(new_n337), .B2(KEYINPUT4), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n343), .ZN(new_n352));
  INV_X1    g151(.A(new_n328), .ZN(new_n353));
  NOR3_X1   g152(.A1(new_n352), .A2(KEYINPUT5), .A3(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n303), .B1(new_n349), .B2(new_n354), .ZN(new_n355));
  XOR2_X1   g154(.A(KEYINPUT82), .B(KEYINPUT6), .Z(new_n356));
  INV_X1    g155(.A(new_n329), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n339), .A2(new_n347), .A3(new_n344), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n347), .B1(new_n339), .B2(new_n344), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n354), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(new_n302), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n355), .A2(new_n356), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n360), .A2(new_n361), .ZN(new_n364));
  INV_X1    g163(.A(new_n356), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n303), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n206), .A2(new_n202), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n227), .A2(new_n229), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n221), .A2(new_n213), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n240), .B(new_n368), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n368), .A2(new_n240), .A3(new_n212), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n225), .A2(new_n226), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n373), .A2(KEYINPUT65), .B1(new_n220), .B2(new_n219), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n215), .A2(new_n216), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(new_n375), .A3(new_n218), .ZN(new_n376));
  AOI22_X1  g175(.A1(KEYINPUT25), .A2(new_n371), .B1(new_n372), .B2(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n244), .B(new_n219), .C1(new_n247), .C2(new_n251), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT29), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G226gat), .A2(G233gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT74), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT29), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n253), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT74), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n385), .A3(new_n380), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n253), .A2(new_n381), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT75), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n380), .B1(new_n377), .B2(new_n378), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT75), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n382), .A2(new_n386), .A3(new_n389), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G211gat), .A2(G218gat), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(G211gat), .A2(G218gat), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT72), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OR2_X1    g195(.A1(G211gat), .A2(G218gat), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT72), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n398), .A3(new_n393), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT22), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n393), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G204gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(G197gat), .ZN(new_n404));
  INV_X1    g203(.A(G197gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(G204gat), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n402), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n400), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n400), .A2(new_n407), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT73), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n400), .A2(KEYINPUT73), .A3(new_n407), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n392), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n381), .B1(new_n253), .B2(new_n383), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n415), .A2(new_n390), .A3(new_n413), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G8gat), .B(G36gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(G64gat), .B(G92gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n414), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT77), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT30), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n416), .B1(new_n392), .B2(new_n413), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT77), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(new_n426), .A3(new_n421), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n423), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n425), .A2(KEYINPUT76), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT76), .ZN(new_n430));
  AOI211_X1 g229(.A(new_n430), .B(new_n416), .C1(new_n392), .C2(new_n413), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n420), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n425), .A2(KEYINPUT30), .A3(new_n421), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n428), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n367), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(G228gat), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n436), .A2(new_n276), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT84), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n400), .A2(KEYINPUT73), .A3(new_n407), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT73), .B1(new_n400), .B2(new_n407), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n411), .A2(KEYINPUT84), .A3(new_n412), .ZN(new_n442));
  INV_X1    g241(.A(new_n408), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n383), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n341), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n333), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT85), .ZN(new_n448));
  INV_X1    g247(.A(new_n413), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT29), .B1(new_n326), .B2(new_n341), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n450), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(KEYINPUT85), .A3(new_n413), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n437), .B1(new_n447), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n341), .B1(new_n413), .B2(KEYINPUT29), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n333), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n437), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n452), .A2(KEYINPUT86), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT86), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n450), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n449), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(G22gat), .B1(new_n456), .B2(new_n464), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n459), .A2(new_n463), .ZN(new_n466));
  INV_X1    g265(.A(new_n437), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n326), .B1(new_n445), .B2(new_n341), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n467), .B1(new_n468), .B2(new_n454), .ZN(new_n469));
  INV_X1    g268(.A(G22gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n466), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  XOR2_X1   g270(.A(G78gat), .B(G106gat), .Z(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(G50gat), .ZN(new_n473));
  XOR2_X1   g272(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n476), .A2(KEYINPUT87), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n465), .A2(new_n471), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n477), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n466), .A2(new_n469), .A3(new_n470), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n466), .A2(new_n469), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(G22gat), .A3(new_n476), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n435), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n298), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n355), .A2(KEYINPUT89), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n346), .A2(new_n348), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n354), .B1(new_n488), .B2(new_n357), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n365), .B1(new_n489), .B2(new_n302), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT89), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n364), .A2(new_n491), .A3(new_n303), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n487), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n423), .A2(new_n427), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT37), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n414), .A2(new_n495), .A3(new_n417), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT90), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT90), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n425), .A2(new_n498), .A3(new_n495), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n421), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n392), .A2(new_n449), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n415), .A2(new_n390), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n495), .B1(new_n502), .B2(new_n413), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT38), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n494), .B1(new_n500), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n493), .A2(new_n366), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT91), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT91), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n493), .A2(new_n508), .A3(new_n366), .A4(new_n505), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n429), .A2(new_n431), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n500), .B1(new_n495), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT38), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n507), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n428), .A2(new_n432), .A3(new_n433), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n328), .B1(new_n351), .B2(new_n343), .ZN(new_n515));
  INV_X1    g314(.A(new_n327), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT39), .B1(new_n516), .B2(new_n353), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n302), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  AOI211_X1 g317(.A(KEYINPUT39), .B(new_n328), .C1(new_n351), .C2(new_n343), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT88), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n520), .A2(KEYINPUT40), .ZN(new_n521));
  OR3_X1    g320(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n521), .B1(new_n518), .B2(new_n519), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n514), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n491), .B1(new_n364), .B2(new_n303), .ZN(new_n525));
  AOI211_X1 g324(.A(KEYINPUT89), .B(new_n302), .C1(new_n360), .C2(new_n361), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n484), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n486), .B1(new_n513), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n366), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n530), .B1(new_n527), .B2(new_n490), .ZN(new_n531));
  INV_X1    g330(.A(new_n296), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT35), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n434), .A2(new_n532), .A3(new_n483), .A4(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n514), .B1(new_n366), .B2(new_n363), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n479), .B1(new_n481), .B2(G22gat), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n470), .B1(new_n466), .B2(new_n469), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n537), .A2(new_n471), .B1(new_n538), .B2(new_n476), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n296), .B1(new_n539), .B2(new_n480), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n533), .B1(new_n536), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n529), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G43gat), .B(G50gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT92), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NOR3_X1   g347(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n549));
  INV_X1    g348(.A(G29gat), .ZN(new_n550));
  INV_X1    g349(.A(G36gat), .ZN(new_n551));
  OAI22_X1  g350(.A1(new_n548), .A2(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n546), .A2(KEYINPUT15), .A3(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT93), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n546), .A2(KEYINPUT15), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n549), .B1(KEYINPUT94), .B2(new_n547), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n556), .B1(KEYINPUT94), .B2(new_n549), .ZN(new_n557));
  OAI22_X1  g356(.A1(new_n544), .A2(KEYINPUT15), .B1(new_n550), .B2(new_n551), .ZN(new_n558));
  OR3_X1    g357(.A1(new_n555), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT17), .ZN(new_n561));
  XNOR2_X1  g360(.A(G15gat), .B(G22gat), .ZN(new_n562));
  INV_X1    g361(.A(G1gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(KEYINPUT16), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n564), .B1(new_n563), .B2(new_n562), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(G8gat), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n561), .B1(new_n566), .B2(KEYINPUT95), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n560), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n554), .A2(new_n559), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT95), .B1(new_n569), .B2(new_n561), .ZN(new_n570));
  INV_X1    g369(.A(new_n566), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n568), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G229gat), .A2(G233gat), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n574), .A2(KEYINPUT18), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(KEYINPUT18), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT96), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n577), .B1(new_n569), .B2(new_n571), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n569), .A2(new_n571), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n569), .A2(new_n577), .A3(new_n571), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n573), .B(KEYINPUT13), .Z(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n575), .A2(new_n576), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G113gat), .B(G141gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT11), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(new_n204), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(G197gat), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n589), .B(KEYINPUT12), .Z(new_n590));
  NAND2_X1  g389(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n590), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n575), .A2(new_n576), .A3(new_n584), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n543), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT21), .ZN(new_n597));
  OR2_X1    g396(.A1(G57gat), .A2(G64gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(G57gat), .A2(G64gat), .ZN(new_n599));
  AND2_X1   g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n598), .B(new_n599), .C1(new_n600), .C2(KEYINPUT9), .ZN(new_n601));
  NOR2_X1   g400(.A1(G71gat), .A2(G78gat), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n601), .B(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n566), .B1(new_n597), .B2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(new_n605), .B(KEYINPUT98), .Z(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n604), .A2(new_n597), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n608), .B(KEYINPUT97), .Z(new_n609));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G127gat), .B(G155gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n611), .A2(new_n612), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n611), .A2(new_n612), .ZN(new_n617));
  INV_X1    g416(.A(new_n614), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G183gat), .B(G211gat), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n615), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n620), .B1(new_n615), .B2(new_n619), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n607), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n623), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(new_n606), .A3(new_n621), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(G99gat), .A2(G106gat), .ZN(new_n628));
  INV_X1    g427(.A(G85gat), .ZN(new_n629));
  INV_X1    g428(.A(G92gat), .ZN(new_n630));
  AOI22_X1  g429(.A1(KEYINPUT8), .A2(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n632), .B1(new_n629), .B2(new_n630), .ZN(new_n633));
  NAND4_X1  g432(.A1(KEYINPUT99), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n631), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(G99gat), .B(G106gat), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n561), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n569), .A2(new_n638), .ZN(new_n639));
  AND2_X1   g438(.A1(G232gat), .A2(G233gat), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n569), .A2(new_n638), .B1(KEYINPUT41), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G190gat), .B(G218gat), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n640), .A2(KEYINPUT41), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n644), .B(new_n645), .C1(KEYINPUT41), .C2(new_n640), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(G134gat), .B(G162gat), .Z(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n651), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n648), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT101), .ZN(new_n656));
  XNOR2_X1  g455(.A(G120gat), .B(G148gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(G230gat), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n660), .A2(new_n276), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n604), .B1(KEYINPUT100), .B2(new_n636), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(new_n637), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT10), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OR3_X1    g464(.A1(new_n637), .A2(new_n604), .A3(new_n664), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n661), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n663), .A2(new_n660), .A3(new_n276), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n659), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n667), .A2(new_n668), .A3(new_n659), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n656), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n671), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n673), .A2(KEYINPUT101), .A3(new_n669), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n627), .A2(new_n655), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n596), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n677), .A2(new_n367), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(new_n563), .ZN(G1324gat));
  NAND3_X1  g478(.A1(new_n596), .A2(new_n514), .A3(new_n676), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT16), .B(G8gat), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n682), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n680), .ZN(new_n683));
  INV_X1    g482(.A(new_n682), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n685), .B1(new_n684), .B2(new_n686), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n683), .B1(new_n688), .B2(new_n689), .ZN(G1325gat));
  OAI21_X1  g489(.A(G15gat), .B1(new_n677), .B2(new_n298), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n296), .A2(G15gat), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n691), .B1(new_n677), .B2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT103), .ZN(G1326gat));
  NOR2_X1   g493(.A1(new_n677), .A2(new_n483), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT43), .B(G22gat), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1327gat));
  AOI21_X1  g496(.A(new_n508), .B1(new_n531), .B2(new_n505), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n509), .A2(new_n512), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n528), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n486), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(new_n541), .B2(new_n535), .ZN(new_n703));
  INV_X1    g502(.A(new_n675), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n627), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n655), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n703), .A2(new_n594), .A3(new_n707), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n708), .A2(G29gat), .A3(new_n367), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT45), .Z(new_n710));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(new_n529), .B2(new_n542), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n705), .A2(new_n595), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n715), .B1(new_n535), .B2(new_n541), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n493), .A2(new_n366), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n717), .A2(new_n533), .A3(new_n434), .A4(new_n540), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n532), .A2(new_n483), .ZN(new_n719));
  OAI21_X1  g518(.A(KEYINPUT35), .B1(new_n435), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n718), .A2(new_n720), .A3(KEYINPUT104), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n706), .B1(new_n702), .B2(new_n722), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n713), .B(new_n714), .C1(new_n723), .C2(KEYINPUT44), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n700), .A2(new_n701), .B1(new_n716), .B2(new_n721), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n711), .B1(new_n727), .B2(new_n706), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n728), .A2(KEYINPUT105), .A3(new_n713), .A4(new_n714), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(G29gat), .B1(new_n730), .B2(new_n367), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n710), .A2(new_n731), .ZN(G1328gat));
  NOR3_X1   g531(.A1(new_n708), .A2(G36gat), .A3(new_n434), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT46), .ZN(new_n734));
  OAI21_X1  g533(.A(G36gat), .B1(new_n730), .B2(new_n434), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(G1329gat));
  NOR2_X1   g535(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n702), .A2(new_n722), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n655), .ZN(new_n739));
  AOI22_X1  g538(.A1(new_n739), .A2(new_n711), .B1(new_n703), .B2(new_n712), .ZN(new_n740));
  INV_X1    g539(.A(new_n298), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n740), .A2(new_n741), .A3(new_n714), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G43gat), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n737), .B1(new_n743), .B2(KEYINPUT47), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n708), .A2(G43gat), .A3(new_n296), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n726), .A2(new_n741), .A3(new_n729), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n746), .A2(G43gat), .B1(KEYINPUT106), .B2(new_n745), .ZN(new_n747));
  OAI22_X1  g546(.A1(new_n744), .A2(new_n745), .B1(new_n747), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g547(.A(G50gat), .B1(new_n724), .B2(new_n483), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n483), .A2(G50gat), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n708), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(KEYINPUT108), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n708), .A2(new_n754), .A3(new_n751), .ZN(new_n755));
  OAI211_X1 g554(.A(KEYINPUT48), .B(new_n749), .C1(new_n753), .C2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n726), .A2(new_n484), .A3(new_n729), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n752), .B1(new_n757), .B2(G50gat), .ZN(new_n758));
  XOR2_X1   g557(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n759));
  OAI21_X1  g558(.A(new_n756), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT109), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n762), .B(new_n756), .C1(new_n758), .C2(new_n759), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(G1331gat));
  NOR2_X1   g563(.A1(new_n627), .A2(new_n655), .ZN(new_n765));
  AND4_X1   g564(.A1(new_n595), .A2(new_n738), .A3(new_n765), .A4(new_n675), .ZN(new_n766));
  INV_X1    g565(.A(new_n367), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g568(.A(new_n434), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n771), .B(new_n772), .Z(G1333gat));
  NAND3_X1  g572(.A1(new_n766), .A2(G71gat), .A3(new_n741), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n766), .A2(new_n532), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n775), .B2(G71gat), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g576(.A1(new_n766), .A2(new_n484), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(G78gat), .ZN(G1335gat));
  INV_X1    g578(.A(new_n627), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n780), .A2(new_n594), .A3(new_n704), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n728), .A2(new_n713), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n767), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n629), .B1(new_n784), .B2(KEYINPUT110), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(KEYINPUT110), .B2(new_n784), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n780), .A2(new_n594), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n738), .A2(KEYINPUT51), .A3(new_n655), .A4(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n723), .A2(KEYINPUT111), .A3(KEYINPUT51), .A4(new_n787), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n535), .A2(new_n541), .A3(new_n715), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT104), .B1(new_n718), .B2(new_n720), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n655), .B(new_n787), .C1(new_n796), .C2(new_n529), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n792), .B1(new_n793), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n767), .A2(new_n629), .A3(new_n675), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n786), .B1(new_n798), .B2(new_n799), .ZN(G1336gat));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801));
  OAI21_X1  g600(.A(G92gat), .B1(new_n782), .B2(new_n434), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n704), .A2(G92gat), .A3(new_n434), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n801), .B(new_n802), .C1(new_n798), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n797), .A2(KEYINPUT112), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n723), .A2(new_n807), .A3(new_n787), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT51), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n803), .B1(new_n792), .B2(new_n809), .ZN(new_n810));
  AOI211_X1 g609(.A(KEYINPUT113), .B(new_n801), .C1(new_n810), .C2(new_n802), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n806), .A2(new_n808), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n813), .A2(new_n793), .B1(new_n790), .B2(new_n791), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n802), .B1(new_n814), .B2(new_n804), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n812), .B1(new_n815), .B2(KEYINPUT52), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n805), .B1(new_n811), .B2(new_n816), .ZN(G1337gat));
  OAI21_X1  g616(.A(G99gat), .B1(new_n782), .B2(new_n298), .ZN(new_n818));
  OR3_X1    g617(.A1(new_n704), .A2(G99gat), .A3(new_n296), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n818), .B1(new_n798), .B2(new_n819), .ZN(G1338gat));
  NAND2_X1  g619(.A1(new_n783), .A2(new_n484), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT53), .B1(new_n821), .B2(G106gat), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n704), .A2(G106gat), .A3(new_n483), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n798), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n814), .A2(new_n824), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n826), .B1(G106gat), .B2(new_n821), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(G1339gat));
  INV_X1    g628(.A(new_n667), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n665), .A2(new_n666), .A3(new_n661), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(KEYINPUT54), .A3(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833));
  INV_X1    g632(.A(new_n659), .ZN(new_n834));
  XOR2_X1   g633(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n835));
  AOI21_X1  g634(.A(new_n834), .B1(new_n667), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n832), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n833), .B1(new_n832), .B2(new_n836), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n673), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n840), .B1(new_n591), .B2(new_n593), .ZN(new_n841));
  INV_X1    g640(.A(new_n583), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n580), .A2(new_n581), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT115), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n844), .B1(new_n573), .B2(new_n572), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n843), .A2(KEYINPUT115), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n589), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n593), .A2(new_n847), .A3(new_n675), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n706), .B1(new_n841), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n840), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n655), .A2(new_n593), .A3(new_n851), .A4(new_n847), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n780), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  NOR4_X1   g652(.A1(new_n627), .A2(new_n594), .A3(new_n655), .A4(new_n675), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT116), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n850), .A2(new_n852), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n627), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n765), .A2(new_n595), .A3(new_n704), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n861), .A2(new_n367), .A3(new_n719), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n862), .A2(new_n434), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n594), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n675), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g666(.A1(new_n863), .A2(new_n780), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g668(.A1(new_n706), .A2(new_n514), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n862), .A2(new_n870), .ZN(new_n871));
  OR3_X1    g670(.A1(new_n871), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT56), .B1(new_n871), .B2(G134gat), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(G134gat), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(G1343gat));
  INV_X1    g674(.A(G141gat), .ZN(new_n876));
  OAI21_X1  g675(.A(KEYINPUT119), .B1(new_n861), .B2(new_n367), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n855), .A2(new_n860), .A3(new_n878), .A4(new_n767), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n741), .A2(new_n483), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n877), .A2(new_n434), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n876), .B1(new_n881), .B2(new_n595), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT117), .B1(new_n832), .B2(new_n836), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n883), .A2(new_n833), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n671), .B1(new_n883), .B2(new_n833), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n594), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n887), .A3(new_n848), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n706), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n887), .B1(new_n886), .B2(new_n848), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n852), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n854), .B1(new_n891), .B2(new_n627), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT57), .B1(new_n892), .B2(new_n483), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n855), .A2(new_n860), .A3(new_n894), .A4(new_n484), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n741), .A2(new_n367), .A3(new_n514), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n595), .A2(new_n876), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n893), .A2(new_n895), .A3(new_n896), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT58), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n882), .A2(KEYINPUT58), .A3(new_n898), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1344gat));
  NAND4_X1  g702(.A1(new_n893), .A2(new_n675), .A3(new_n895), .A4(new_n896), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(new_n905), .A3(G148gat), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT120), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n886), .A2(new_n848), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT118), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n706), .A3(new_n888), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n780), .B1(new_n910), .B2(new_n852), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n894), .B(new_n484), .C1(new_n911), .C2(new_n854), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n861), .A2(new_n483), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n913), .B2(new_n894), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n896), .A2(new_n675), .ZN(new_n915));
  OAI21_X1  g714(.A(G148gat), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT59), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n904), .A2(new_n918), .A3(new_n905), .A4(G148gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n907), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  OR3_X1    g719(.A1(new_n881), .A2(G148gat), .A3(new_n704), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1345gat));
  NAND3_X1  g721(.A1(new_n893), .A2(new_n895), .A3(new_n896), .ZN(new_n923));
  OAI21_X1  g722(.A(G155gat), .B1(new_n923), .B2(new_n627), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n780), .A2(new_n311), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n881), .B2(new_n925), .ZN(G1346gat));
  OAI21_X1  g725(.A(G162gat), .B1(new_n923), .B2(new_n706), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n879), .A2(new_n880), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n877), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n870), .A2(new_n312), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(G1347gat));
  AND2_X1   g730(.A1(new_n855), .A2(new_n860), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n367), .A2(new_n514), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n933), .A2(new_n719), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n935), .A2(new_n204), .A3(new_n595), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n855), .A2(new_n860), .A3(new_n367), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT121), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n855), .A2(new_n860), .A3(KEYINPUT121), .A4(new_n367), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n434), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n941), .A2(new_n540), .A3(new_n594), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n936), .B1(new_n942), .B2(new_n204), .ZN(G1348gat));
  NOR3_X1   g742(.A1(new_n935), .A2(new_n205), .A3(new_n704), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n939), .A2(new_n940), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n945), .A2(new_n514), .A3(new_n540), .A4(new_n675), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n944), .B1(new_n946), .B2(new_n205), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n947), .A2(KEYINPUT122), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT122), .ZN(new_n949));
  AOI211_X1 g748(.A(new_n949), .B(new_n944), .C1(new_n946), .C2(new_n205), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n948), .A2(new_n950), .ZN(G1349gat));
  AND2_X1   g750(.A1(new_n780), .A2(new_n246), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n941), .A2(new_n540), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(G183gat), .B1(new_n935), .B2(new_n627), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g755(.A(G190gat), .B1(new_n935), .B2(new_n706), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT61), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n941), .A2(new_n226), .A3(new_n540), .A4(new_n655), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1351gat));
  NAND4_X1  g759(.A1(new_n941), .A2(new_n405), .A3(new_n594), .A4(new_n880), .ZN(new_n961));
  OR2_X1    g760(.A1(new_n961), .A2(KEYINPUT123), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(KEYINPUT123), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n914), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n912), .B(KEYINPUT124), .C1(new_n913), .C2(new_n894), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n741), .A2(new_n933), .ZN(new_n967));
  AND4_X1   g766(.A1(new_n594), .A2(new_n965), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n962), .B(new_n963), .C1(new_n968), .C2(new_n405), .ZN(G1352gat));
  XOR2_X1   g768(.A(KEYINPUT125), .B(G204gat), .Z(new_n970));
  NAND3_X1  g769(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n970), .B1(new_n971), .B2(new_n704), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n704), .A2(new_n970), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n945), .A2(new_n514), .A3(new_n880), .A4(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n972), .A2(new_n976), .ZN(G1353gat));
  NOR2_X1   g776(.A1(new_n627), .A2(G211gat), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n941), .A2(new_n880), .A3(new_n978), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n979), .B(KEYINPUT126), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n741), .A2(new_n627), .A3(new_n933), .ZN(new_n981));
  OAI211_X1 g780(.A(new_n912), .B(new_n981), .C1(new_n913), .C2(new_n894), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(G211gat), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT63), .ZN(new_n984));
  XNOR2_X1  g783(.A(new_n983), .B(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n980), .A2(new_n985), .ZN(G1354gat));
  OAI21_X1  g785(.A(G218gat), .B1(new_n971), .B2(new_n706), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n706), .A2(G218gat), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n941), .A2(new_n880), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n987), .A2(new_n989), .ZN(G1355gat));
endmodule


