//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 1 0 1 0 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1034, new_n1035,
    new_n1036, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  OAI21_X1  g001(.A(G210), .B1(G237), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G116), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT2), .B(G113), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT71), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT2), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G113), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(G116), .B(G119), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT71), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n190), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT5), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n196), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n201), .A2(KEYINPUT5), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n195), .A2(new_n203), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G104), .ZN(new_n209));
  NOR3_X1   g023(.A1(new_n209), .A2(KEYINPUT3), .A3(G107), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G104), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT3), .B1(new_n209), .B2(G107), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n213), .A2(KEYINPUT83), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(new_n211), .A3(G104), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n209), .A2(G107), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n215), .A2(new_n218), .A3(new_n214), .A4(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT83), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n216), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n211), .A2(G104), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n224), .A2(new_n219), .A3(KEYINPUT85), .ZN(new_n225));
  OAI21_X1  g039(.A(G101), .B1(new_n224), .B2(KEYINPUT85), .ZN(new_n226));
  OR2_X1    g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n208), .A2(new_n223), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n215), .A2(new_n218), .A3(new_n219), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G101), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT4), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n231), .B1(new_n222), .B2(new_n216), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n193), .A2(new_n194), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n200), .A2(new_n201), .A3(new_n202), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n202), .B1(new_n200), .B2(new_n201), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n229), .A2(new_n237), .A3(G101), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n228), .B1(new_n232), .B2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G110), .B(G122), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT89), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT6), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n240), .A2(new_n242), .A3(new_n245), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n229), .A2(new_n237), .A3(G101), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n195), .A2(new_n203), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n247), .B1(new_n248), .B2(new_n233), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n237), .B1(new_n229), .B2(G101), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n220), .A2(new_n221), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n220), .A2(new_n221), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n225), .A2(new_n226), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n254), .B1(new_n216), .B2(new_n222), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n249), .A2(new_n253), .B1(new_n255), .B2(new_n208), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n244), .B1(new_n256), .B2(new_n241), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(new_n241), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n246), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G146), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G143), .ZN(new_n261));
  INV_X1    g075(.A(G143), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G146), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(KEYINPUT0), .A2(G128), .ZN(new_n265));
  OR2_X1    g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(G143), .B(G146), .ZN(new_n268));
  AND2_X1   g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT64), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AND4_X1   g084(.A1(KEYINPUT64), .A2(new_n261), .A3(new_n263), .A4(new_n269), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n267), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT1), .B1(new_n262), .B2(G146), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n262), .A2(G146), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n260), .A2(G143), .ZN(new_n275));
  OAI211_X1 g089(.A(G128), .B(new_n273), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G128), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n261), .B(new_n263), .C1(KEYINPUT1), .C2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(G125), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT90), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n272), .A2(G125), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(KEYINPUT91), .B(G224), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n282), .A2(G953), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  OR2_X1    g098(.A1(new_n279), .A2(new_n280), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n281), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n284), .B1(new_n281), .B2(new_n285), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n259), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT92), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT92), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n259), .A2(new_n292), .A3(new_n289), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n281), .A2(new_n285), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT7), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n296), .B1(new_n297), .B2(new_n283), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n228), .B(new_n241), .C1(new_n232), .C2(new_n239), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n281), .A2(new_n285), .A3(KEYINPUT7), .A4(new_n284), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  XOR2_X1   g115(.A(new_n241), .B(KEYINPUT8), .Z(new_n302));
  INV_X1    g116(.A(new_n208), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n227), .B1(new_n251), .B2(new_n252), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n302), .B1(new_n305), .B2(new_n228), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n295), .B1(new_n301), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n188), .B1(new_n294), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n299), .A2(new_n245), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n240), .A2(new_n242), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI211_X1 g126(.A(KEYINPUT92), .B(new_n288), .C1(new_n312), .C2(new_n246), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n292), .B1(new_n259), .B2(new_n289), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n188), .B(new_n308), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n187), .B1(new_n309), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G221), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT9), .B(G234), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n318), .B1(new_n320), .B2(new_n295), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(G110), .B(G140), .ZN(new_n323));
  INV_X1    g137(.A(G953), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n324), .A2(G227), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n323), .B(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT11), .ZN(new_n327));
  INV_X1    g141(.A(G134), .ZN(new_n328));
  OAI211_X1 g142(.A(KEYINPUT65), .B(new_n327), .C1(new_n328), .C2(G137), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n328), .A2(KEYINPUT67), .A3(G137), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT67), .B1(new_n328), .B2(G137), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT65), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(KEYINPUT11), .ZN(new_n334));
  INV_X1    g148(.A(G137), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G134), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(KEYINPUT11), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(G131), .B1(new_n332), .B2(new_n338), .ZN(new_n339));
  OAI22_X1  g153(.A1(KEYINPUT65), .A2(new_n327), .B1(new_n328), .B2(G137), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n327), .A2(KEYINPUT65), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(KEYINPUT66), .A2(G131), .ZN(new_n343));
  NOR2_X1   g157(.A1(KEYINPUT66), .A2(G131), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT67), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(new_n335), .B2(G134), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n328), .A2(KEYINPUT67), .A3(G137), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n342), .A2(new_n345), .A3(new_n349), .A4(new_n329), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n339), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n261), .A2(new_n263), .A3(new_n269), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT64), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n268), .A2(KEYINPUT64), .A3(new_n269), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n266), .A2(new_n265), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n355), .A2(new_n356), .B1(new_n264), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n238), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT84), .B1(new_n232), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n272), .A2(new_n247), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT84), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n253), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n276), .A2(KEYINPUT72), .A3(new_n278), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT72), .B1(new_n276), .B2(new_n278), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT10), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT87), .B1(new_n367), .B2(new_n304), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n276), .A2(new_n278), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT72), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n276), .A2(KEYINPUT72), .A3(new_n278), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT87), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n373), .A2(new_n374), .A3(new_n255), .A4(KEYINPUT10), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n368), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT86), .B(KEYINPUT10), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n369), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n378), .B1(new_n255), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  AND4_X1   g195(.A1(new_n352), .A2(new_n364), .A3(new_n376), .A4(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n380), .B1(new_n360), .B2(new_n363), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n352), .B1(new_n383), .B2(new_n376), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n326), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT12), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n304), .A2(new_n369), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n255), .A2(new_n379), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n386), .B1(new_n389), .B2(new_n351), .ZN(new_n390));
  AOI211_X1 g204(.A(KEYINPUT12), .B(new_n352), .C1(new_n387), .C2(new_n388), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n364), .A2(new_n376), .A3(new_n352), .A4(new_n381), .ZN(new_n393));
  INV_X1    g207(.A(new_n326), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  AOI211_X1 g209(.A(G469), .B(G902), .C1(new_n385), .C2(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n304), .A2(new_n369), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n255), .A2(new_n379), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n351), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT12), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n389), .A2(new_n386), .A3(new_n351), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n326), .B1(new_n382), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n376), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n361), .A2(new_n253), .A3(new_n362), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n362), .B1(new_n361), .B2(new_n253), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n381), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n351), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n393), .A3(new_n394), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n403), .A2(G469), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G469), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(new_n295), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n322), .B1(new_n396), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT88), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g231(.A(KEYINPUT88), .B(new_n322), .C1(new_n396), .C2(new_n414), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n317), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT28), .ZN(new_n420));
  OR3_X1    g234(.A1(new_n335), .A2(KEYINPUT69), .A3(G134), .ZN(new_n421));
  INV_X1    g235(.A(new_n336), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT69), .B1(new_n335), .B2(G134), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n421), .B(G131), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n350), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n373), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n236), .ZN(new_n427));
  INV_X1    g241(.A(new_n345), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n332), .A2(new_n338), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G131), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n347), .A2(new_n348), .B1(new_n334), .B2(new_n336), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n430), .B1(new_n431), .B2(new_n342), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n358), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n426), .A2(new_n427), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT74), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n373), .A2(new_n425), .B1(new_n351), .B2(new_n358), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(KEYINPUT74), .A3(new_n427), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT68), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n358), .B(new_n441), .C1(new_n429), .C2(new_n432), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n441), .B1(new_n351), .B2(new_n358), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n350), .A2(new_n278), .A3(new_n276), .A4(new_n424), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT70), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n379), .A2(KEYINPUT70), .A3(new_n350), .A4(new_n424), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n236), .B1(new_n445), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n420), .B1(new_n440), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n434), .A2(new_n420), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(G237), .A2(G953), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G210), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(KEYINPUT27), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT26), .B(G101), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n457), .B(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n452), .A2(new_n454), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT73), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n433), .A2(KEYINPUT68), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n442), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n448), .A2(new_n449), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT30), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n437), .A2(KEYINPUT30), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n236), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n462), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n427), .B1(new_n437), .B2(KEYINPUT30), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n450), .B1(new_n463), .B2(new_n442), .ZN(new_n471));
  OAI211_X1 g285(.A(KEYINPUT73), .B(new_n470), .C1(new_n471), .C2(KEYINPUT30), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n459), .B1(new_n473), .B2(new_n440), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n461), .A2(new_n474), .A3(KEYINPUT29), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n436), .B(new_n438), .C1(new_n427), .C2(new_n437), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT28), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n459), .A2(KEYINPUT29), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n453), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT75), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n477), .A2(KEYINPUT75), .A3(new_n453), .A4(new_n478), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n295), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(G472), .B1(new_n475), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n460), .B1(new_n452), .B2(new_n454), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n436), .A2(new_n438), .A3(new_n459), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT31), .B1(new_n473), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT31), .ZN(new_n489));
  AOI211_X1 g303(.A(new_n489), .B(new_n486), .C1(new_n469), .C2(new_n472), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n485), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT32), .ZN(new_n492));
  NOR2_X1   g306(.A1(G472), .A2(G902), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n492), .B1(new_n491), .B2(new_n493), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n484), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT25), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT22), .B(G137), .ZN(new_n498));
  INV_X1    g312(.A(G234), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n318), .A2(new_n499), .A3(G953), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n498), .B(new_n500), .Z(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n189), .A2(G128), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n277), .A2(G119), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT77), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n277), .A2(G119), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n189), .A2(G128), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT77), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  XOR2_X1   g323(.A(KEYINPUT24), .B(G110), .Z(new_n510));
  NAND3_X1  g324(.A1(new_n505), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(G140), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G125), .ZN(new_n513));
  INV_X1    g327(.A(G125), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(G140), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(new_n515), .A3(KEYINPUT16), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n514), .A2(G140), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT16), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n516), .A2(new_n519), .A3(G146), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(G146), .B1(new_n516), .B2(new_n519), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n277), .A2(KEYINPUT23), .A3(G119), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n523), .B(new_n507), .C1(new_n503), .C2(KEYINPUT23), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G110), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(KEYINPUT78), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT78), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n527), .B1(new_n524), .B2(G110), .ZN(new_n528));
  OAI221_X1 g342(.A(new_n511), .B1(new_n521), .B2(new_n522), .C1(new_n526), .C2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n513), .A2(new_n515), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT79), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n513), .A2(new_n515), .A3(KEYINPUT79), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(new_n260), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n510), .B1(new_n505), .B2(new_n509), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n524), .A2(G110), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n520), .B(new_n534), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT80), .B1(new_n529), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n526), .A2(new_n528), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n511), .B1(new_n521), .B2(new_n522), .ZN(new_n540));
  OAI211_X1 g354(.A(KEYINPUT80), .B(new_n537), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n502), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n501), .ZN(new_n545));
  AOI21_X1  g359(.A(G902), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g360(.A(KEYINPUT82), .B(new_n497), .C1(new_n546), .C2(KEYINPUT81), .ZN(new_n547));
  OAI21_X1  g361(.A(G217), .B1(new_n499), .B2(G902), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(KEYINPUT76), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT80), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n501), .B1(new_n551), .B2(new_n541), .ZN(new_n552));
  INV_X1    g366(.A(new_n545), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n295), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT82), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT25), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT81), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n555), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n547), .B(new_n549), .C1(new_n557), .C2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n549), .A2(G902), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(new_n552), .B2(new_n553), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT94), .ZN(new_n565));
  INV_X1    g379(.A(G237), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(new_n324), .A3(G214), .ZN(new_n567));
  NOR2_X1   g381(.A1(KEYINPUT93), .A2(G143), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n455), .B(G214), .C1(KEYINPUT93), .C2(G143), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n428), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n570), .A3(new_n345), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n521), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT19), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n532), .A2(new_n575), .A3(new_n533), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n530), .A2(KEYINPUT19), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(new_n260), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(KEYINPUT18), .A2(G131), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n569), .A2(new_n570), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n579), .B1(new_n569), .B2(new_n570), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n530), .A2(G146), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n534), .A2(new_n584), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n574), .A2(new_n578), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(G113), .B(G122), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(new_n209), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n565), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n583), .A2(new_n585), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT17), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n572), .A2(KEYINPUT95), .A3(new_n591), .A4(new_n573), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n521), .A2(new_n522), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n345), .B1(new_n569), .B2(new_n570), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT17), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n569), .A2(new_n570), .A3(new_n345), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(new_n594), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT95), .B1(new_n598), .B2(new_n591), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n588), .B(new_n590), .C1(new_n596), .C2(new_n599), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n576), .A2(new_n260), .A3(new_n577), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n520), .B1(new_n597), .B2(new_n594), .ZN(new_n602));
  INV_X1    g416(.A(new_n584), .ZN(new_n603));
  INV_X1    g417(.A(new_n533), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT79), .B1(new_n513), .B2(new_n515), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n603), .B1(new_n606), .B2(new_n260), .ZN(new_n607));
  INV_X1    g421(.A(new_n579), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n571), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n580), .ZN(new_n610));
  OAI22_X1  g424(.A1(new_n601), .A2(new_n602), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n588), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(KEYINPUT94), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n589), .A2(new_n600), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT96), .ZN(new_n615));
  NOR2_X1   g429(.A1(G475), .A2(G902), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT96), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n589), .A2(new_n613), .A3(new_n600), .A4(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n615), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT20), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT20), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n614), .A2(new_n621), .A3(new_n616), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n590), .B1(new_n596), .B2(new_n599), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n612), .ZN(new_n625));
  AOI21_X1  g439(.A(G902), .B1(new_n625), .B2(new_n600), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n627));
  OAI21_X1  g441(.A(G475), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI211_X1 g442(.A(KEYINPUT97), .B(G902), .C1(new_n625), .C2(new_n600), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n623), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n262), .A2(G128), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n277), .A2(G143), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n633), .A2(new_n634), .A3(new_n328), .ZN(new_n635));
  INV_X1    g449(.A(G122), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G116), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n191), .A2(G122), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(G107), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n637), .A2(new_n638), .A3(new_n211), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n635), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT13), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n633), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n634), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n633), .A2(new_n643), .ZN(new_n646));
  OAI21_X1  g460(.A(G134), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n191), .A2(KEYINPUT14), .A3(G122), .ZN(new_n649));
  OAI211_X1 g463(.A(G107), .B(new_n649), .C1(new_n639), .C2(KEYINPUT14), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n328), .B1(new_n633), .B2(new_n634), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n650), .B(new_n641), .C1(new_n635), .C2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n320), .A2(G217), .A3(new_n324), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT98), .ZN(new_n656));
  INV_X1    g470(.A(new_n654), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n648), .A2(new_n652), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n653), .A2(KEYINPUT98), .A3(new_n654), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n295), .A3(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(G478), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(KEYINPUT15), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n661), .B(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT99), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n324), .A2(G952), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n668), .B1(new_n499), .B2(new_n566), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  AOI211_X1 g484(.A(new_n295), .B(new_n324), .C1(G234), .C2(G237), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT21), .B(G898), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n666), .A2(new_n667), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n632), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n419), .A2(new_n496), .A3(new_n564), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G101), .ZN(G3));
  OAI21_X1  g492(.A(new_n308), .B1(new_n313), .B2(new_n314), .ZN(new_n679));
  INV_X1    g493(.A(new_n188), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(KEYINPUT100), .A3(new_n315), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT100), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n679), .A2(new_n683), .A3(new_n680), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n682), .A2(new_n674), .A3(new_n187), .A4(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n686));
  AOI21_X1  g500(.A(KEYINPUT33), .B1(new_n659), .B2(new_n660), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT33), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n657), .B1(new_n648), .B2(new_n652), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT101), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n658), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n648), .A2(new_n652), .A3(KEYINPUT101), .A4(new_n657), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n688), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n295), .B1(new_n687), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(G478), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n661), .A2(G478), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n686), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  AOI211_X1 g512(.A(KEYINPUT102), .B(new_n696), .C1(new_n694), .C2(G478), .ZN(new_n699));
  INV_X1    g513(.A(new_n622), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n619), .B2(KEYINPUT20), .ZN(new_n701));
  OAI22_X1  g515(.A1(new_n698), .A2(new_n699), .B1(new_n701), .B2(new_n630), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n685), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n417), .A2(new_n418), .ZN(new_n704));
  INV_X1    g518(.A(G472), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n705), .B1(new_n491), .B2(new_n295), .ZN(new_n706));
  INV_X1    g520(.A(new_n493), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n466), .A2(new_n468), .A3(new_n462), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT30), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n709), .B1(new_n445), .B2(new_n450), .ZN(new_n710));
  AOI21_X1  g524(.A(KEYINPUT73), .B1(new_n710), .B2(new_n470), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n487), .B1(new_n708), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n489), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n473), .A2(KEYINPUT31), .A3(new_n487), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n707), .B1(new_n715), .B2(new_n485), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n706), .A2(new_n716), .A3(new_n563), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n703), .A2(new_n704), .A3(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT34), .B(G104), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G6));
  NAND4_X1  g534(.A1(new_n615), .A2(new_n621), .A3(new_n616), .A4(new_n618), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n620), .A2(KEYINPUT103), .A3(new_n721), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n722), .A2(new_n631), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n666), .A2(new_n667), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n620), .A2(new_n721), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT103), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n723), .A2(new_n724), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n685), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n704), .A3(new_n717), .ZN(new_n730));
  XOR2_X1   g544(.A(KEYINPUT35), .B(G107), .Z(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G9));
  INV_X1    g546(.A(new_n317), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n706), .A2(new_n716), .ZN(new_n734));
  OAI21_X1  g548(.A(KEYINPUT82), .B1(new_n546), .B2(KEYINPUT81), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n556), .A3(KEYINPUT25), .ZN(new_n736));
  INV_X1    g550(.A(new_n549), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n737), .B1(new_n559), .B2(new_n497), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n551), .A2(new_n541), .ZN(new_n739));
  OR2_X1    g553(.A1(new_n502), .A2(KEYINPUT36), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n736), .A2(new_n738), .B1(new_n561), .B2(new_n741), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n742), .A2(new_n632), .A3(new_n675), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n704), .A2(new_n733), .A3(new_n734), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT104), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT37), .B(G110), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G12));
  AND3_X1   g561(.A1(new_n681), .A2(KEYINPUT100), .A3(new_n315), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n684), .A2(new_n187), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n742), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n496), .A2(new_n704), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(G900), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n671), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n669), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n728), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n752), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n277), .ZN(G30));
  XNOR2_X1  g574(.A(new_n755), .B(KEYINPUT39), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n704), .A2(new_n761), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n762), .A2(KEYINPUT40), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(KEYINPUT40), .ZN(new_n764));
  INV_X1    g578(.A(new_n451), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT28), .B1(new_n765), .B2(new_n439), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n459), .B1(new_n766), .B2(new_n453), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n767), .B1(new_n713), .B2(new_n714), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT32), .B1(new_n768), .B2(new_n707), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n476), .A2(new_n460), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT105), .ZN(new_n773));
  INV_X1    g587(.A(new_n712), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n295), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(G472), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n751), .B1(new_n771), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n309), .A2(new_n316), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT38), .ZN(new_n779));
  AOI22_X1  g593(.A1(new_n623), .A2(new_n631), .B1(new_n666), .B2(new_n667), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n187), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n763), .A2(new_n764), .A3(new_n777), .A4(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT106), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(new_n262), .ZN(G45));
  INV_X1    g602(.A(new_n698), .ZN(new_n789));
  INV_X1    g603(.A(new_n699), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n632), .A3(new_n755), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n752), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(KEYINPUT107), .B(G146), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n793), .B(new_n794), .ZN(G48));
  INV_X1    g609(.A(new_n395), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n394), .B1(new_n408), .B2(new_n393), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n295), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(G469), .ZN(new_n799));
  AOI21_X1  g613(.A(G902), .B1(new_n385), .B2(new_n395), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n411), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n799), .A2(new_n801), .A3(new_n322), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n703), .A2(new_n496), .A3(new_n564), .A4(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(KEYINPUT41), .B(G113), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n804), .B(new_n805), .ZN(G15));
  NAND4_X1  g620(.A1(new_n729), .A2(new_n496), .A3(new_n564), .A4(new_n803), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G116), .ZN(G18));
  NOR3_X1   g622(.A1(new_n748), .A2(new_n802), .A3(new_n749), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n496), .A2(new_n809), .A3(new_n676), .A4(new_n751), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G119), .ZN(G21));
  NAND2_X1  g625(.A1(new_n477), .A2(new_n453), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n460), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n707), .B1(new_n715), .B2(new_n813), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n706), .A2(new_n814), .A3(new_n563), .ZN(new_n815));
  INV_X1    g629(.A(new_n187), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n816), .B1(new_n309), .B2(new_n683), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n817), .A2(new_n682), .A3(new_n780), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n802), .A2(new_n673), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n815), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G122), .ZN(G24));
  NOR3_X1   g635(.A1(new_n706), .A2(new_n814), .A3(new_n742), .ZN(new_n822));
  INV_X1    g636(.A(new_n792), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(new_n809), .A3(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G125), .ZN(G27));
  AND3_X1   g639(.A1(new_n681), .A2(new_n187), .A3(new_n315), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n392), .A2(new_n393), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT108), .B1(new_n827), .B2(new_n326), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT108), .ZN(new_n829));
  AOI211_X1 g643(.A(new_n829), .B(new_n394), .C1(new_n392), .C2(new_n393), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n409), .A2(KEYINPUT109), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT109), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n408), .A2(new_n833), .A3(new_n393), .A4(new_n394), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n831), .A2(new_n835), .A3(G469), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n412), .B1(new_n800), .B2(new_n411), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n826), .A2(new_n838), .A3(new_n322), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT110), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(KEYINPUT42), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n792), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n496), .A2(new_n839), .A3(new_n564), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n840), .A2(KEYINPUT42), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n563), .B1(new_n771), .B2(new_n484), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n847), .A2(new_n839), .A3(new_n842), .A4(new_n844), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(new_n430), .ZN(G33));
  NAND3_X1  g664(.A1(new_n847), .A2(new_n757), .A3(new_n839), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(G134), .ZN(G36));
  INV_X1    g666(.A(new_n826), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n701), .A2(new_n630), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n791), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT112), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT43), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n855), .B(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n734), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n858), .A2(new_n859), .A3(new_n751), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT44), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n853), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n862), .B1(new_n861), .B2(new_n860), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT113), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n831), .A2(new_n835), .A3(KEYINPUT45), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT45), .B1(new_n403), .B2(new_n409), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n411), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n865), .A2(KEYINPUT111), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT111), .B1(new_n865), .B2(new_n867), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n413), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT46), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n396), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(KEYINPUT46), .B(new_n413), .C1(new_n868), .C2(new_n869), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n321), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n874), .A2(new_n761), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n864), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(G137), .ZN(G39));
  OR2_X1    g691(.A1(new_n874), .A2(KEYINPUT47), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n874), .A2(KEYINPUT47), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR4_X1   g694(.A1(new_n496), .A2(new_n564), .A3(new_n792), .A4(new_n853), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(G140), .ZN(G42));
  AND2_X1   g697(.A1(new_n858), .A2(new_n670), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n815), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n803), .A2(new_n816), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n886), .A2(KEYINPUT118), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(KEYINPUT118), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n887), .A2(new_n779), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT50), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n853), .A2(new_n802), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n884), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n814), .ZN(new_n894));
  OAI21_X1  g708(.A(G472), .B1(new_n768), .B2(G902), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n895), .A3(new_n751), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n776), .B1(new_n494), .B2(new_n495), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  AND4_X1   g713(.A1(new_n564), .A2(new_n899), .A3(new_n670), .A4(new_n892), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n791), .A2(new_n632), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n891), .A2(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n799), .A2(new_n801), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n321), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n878), .A2(new_n879), .A3(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n885), .A2(new_n853), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT117), .Z(new_n908));
  AOI21_X1  g722(.A(new_n903), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  XOR2_X1   g723(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n910));
  OAI21_X1  g724(.A(KEYINPUT119), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n884), .A2(new_n847), .A3(new_n892), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT48), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n884), .A2(new_n809), .A3(new_n815), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n900), .A2(new_n632), .A3(new_n791), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n913), .A2(new_n668), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n909), .B2(KEYINPUT51), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT119), .ZN(new_n918));
  INV_X1    g732(.A(new_n910), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n908), .A2(new_n906), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n918), .B(new_n919), .C1(new_n920), .C2(new_n903), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n911), .A2(new_n917), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT115), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n846), .A2(new_n848), .A3(new_n851), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n822), .A2(new_n839), .A3(new_n823), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n496), .A2(new_n704), .A3(new_n751), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n664), .A2(new_n756), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n723), .A2(new_n727), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT114), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT114), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n723), .A2(new_n727), .A3(new_n930), .A4(new_n927), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n826), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n925), .B1(new_n926), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n924), .A2(new_n933), .ZN(new_n934));
  AND4_X1   g748(.A1(new_n496), .A2(new_n704), .A3(new_n750), .A4(new_n751), .ZN(new_n935));
  AOI211_X1 g749(.A(new_n321), .B(new_n756), .C1(new_n836), .C2(new_n837), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n818), .A2(new_n936), .ZN(new_n937));
  AOI22_X1  g751(.A1(new_n935), .A2(new_n823), .B1(new_n777), .B2(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n904), .A2(new_n817), .A3(new_n322), .A4(new_n682), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n896), .A2(new_n939), .A3(new_n792), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n935), .B2(new_n757), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT52), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n938), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n677), .A2(new_n807), .A3(new_n804), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n623), .A2(new_n631), .A3(new_n664), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n702), .A2(new_n945), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n674), .B(new_n187), .C1(new_n309), .C2(new_n316), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n948), .A2(new_n717), .A3(new_n704), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n810), .A2(new_n949), .A3(new_n744), .A4(new_n820), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n944), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n824), .B1(new_n752), .B2(new_n758), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n898), .A2(new_n818), .A3(new_n936), .A4(new_n742), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n752), .B2(new_n792), .ZN(new_n954));
  OAI21_X1  g768(.A(KEYINPUT52), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n934), .A2(new_n943), .A3(new_n951), .A4(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT53), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n923), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n942), .B1(new_n938), .B2(new_n941), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n952), .A2(new_n954), .A3(KEYINPUT52), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NOR4_X1   g775(.A1(new_n924), .A2(new_n944), .A3(new_n950), .A4(new_n933), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n961), .A2(KEYINPUT115), .A3(KEYINPUT53), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n956), .A2(new_n957), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n958), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(KEYINPUT54), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n961), .A2(KEYINPUT53), .A3(new_n962), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT54), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n967), .A2(new_n964), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  OAI22_X1  g784(.A1(new_n922), .A2(new_n970), .B1(G952), .B2(G953), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n904), .B(KEYINPUT49), .ZN(new_n972));
  NOR4_X1   g786(.A1(new_n855), .A2(new_n563), .A3(new_n321), .A4(new_n816), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n899), .A2(new_n972), .A3(new_n779), .A4(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n971), .A2(new_n974), .ZN(G75));
  NOR2_X1   g789(.A1(new_n324), .A2(G952), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n295), .B1(new_n967), .B2(new_n964), .ZN(new_n978));
  AOI21_X1  g792(.A(KEYINPUT56), .B1(new_n978), .B2(G210), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n259), .B(new_n288), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT55), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n977), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n982), .B1(new_n979), .B2(new_n981), .ZN(G51));
  AOI21_X1  g797(.A(KEYINPUT53), .B1(new_n961), .B2(new_n962), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n943), .A2(new_n955), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n846), .A2(new_n848), .A3(new_n851), .ZN(new_n986));
  INV_X1    g800(.A(new_n933), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n951), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n985), .A2(new_n988), .A3(new_n957), .ZN(new_n989));
  OAI21_X1  g803(.A(KEYINPUT54), .B1(new_n984), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n990), .A2(KEYINPUT120), .A3(new_n969), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n967), .A2(new_n964), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT120), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n992), .A2(new_n993), .A3(KEYINPUT54), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n412), .B(KEYINPUT57), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n991), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(new_n797), .B2(new_n796), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n868), .A2(new_n869), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n978), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n976), .B1(new_n997), .B2(new_n999), .ZN(G54));
  NAND2_X1  g814(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT121), .Z(new_n1002));
  NAND2_X1  g816(.A1(new_n978), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n615), .A2(new_n618), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n1005), .A2(new_n1006), .A3(new_n976), .ZN(G60));
  OR2_X1    g821(.A1(new_n687), .A2(new_n693), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g823(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n662), .A2(new_n295), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1010), .B(new_n1011), .Z(new_n1012));
  INV_X1    g826(.A(new_n1012), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1009), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n991), .A2(new_n994), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n977), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1008), .B1(new_n970), .B2(new_n1012), .ZN(new_n1017));
  OAI21_X1  g831(.A(KEYINPUT123), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AND3_X1   g832(.A1(new_n967), .A2(new_n964), .A3(new_n968), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1019), .B1(KEYINPUT54), .B2(new_n965), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1009), .B1(new_n1020), .B2(new_n1013), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT123), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1021), .A2(new_n1022), .A3(new_n977), .A4(new_n1015), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1018), .A2(new_n1023), .ZN(G63));
  NAND2_X1  g838(.A1(G217), .A2(G902), .ZN(new_n1025));
  XOR2_X1   g839(.A(new_n1025), .B(KEYINPUT60), .Z(new_n1026));
  NAND2_X1  g840(.A1(new_n992), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n552), .A2(new_n553), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n976), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(new_n741), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1029), .B1(new_n1030), .B2(new_n1027), .ZN(new_n1031));
  INV_X1    g845(.A(KEYINPUT61), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1031), .B(new_n1032), .ZN(G66));
  OAI21_X1  g847(.A(G953), .B1(new_n672), .B2(new_n282), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1034), .B1(new_n951), .B2(G953), .ZN(new_n1035));
  OAI211_X1 g849(.A(new_n312), .B(new_n246), .C1(G898), .C2(new_n324), .ZN(new_n1036));
  XNOR2_X1  g850(.A(new_n1035), .B(new_n1036), .ZN(G69));
  AND2_X1   g851(.A1(new_n710), .A2(new_n467), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n576), .A2(new_n577), .ZN(new_n1039));
  XOR2_X1   g853(.A(new_n1038), .B(new_n1039), .Z(new_n1040));
  OAI211_X1 g854(.A(G900), .B(G953), .C1(new_n1040), .C2(G227), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1041), .B1(G227), .B2(new_n1040), .ZN(new_n1042));
  AOI22_X1  g856(.A1(new_n864), .A2(new_n875), .B1(new_n880), .B2(new_n881), .ZN(new_n1043));
  INV_X1    g857(.A(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g858(.A(new_n924), .B(KEYINPUT125), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n952), .A2(new_n793), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n875), .A2(new_n847), .A3(new_n818), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g862(.A(KEYINPUT126), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g863(.A(KEYINPUT126), .ZN(new_n1050));
  INV_X1    g864(.A(new_n1048), .ZN(new_n1051));
  NAND3_X1  g865(.A1(new_n1043), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  NAND3_X1  g866(.A1(new_n1049), .A2(new_n1052), .A3(new_n1040), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n785), .A2(new_n786), .A3(new_n1046), .ZN(new_n1054));
  INV_X1    g868(.A(KEYINPUT62), .ZN(new_n1055));
  XNOR2_X1  g869(.A(new_n1054), .B(new_n1055), .ZN(new_n1056));
  INV_X1    g870(.A(new_n946), .ZN(new_n1057));
  AND2_X1   g871(.A1(new_n1057), .A2(KEYINPUT124), .ZN(new_n1058));
  NOR2_X1   g872(.A1(new_n1057), .A2(KEYINPUT124), .ZN(new_n1059));
  NOR3_X1   g873(.A1(new_n1058), .A2(new_n1059), .A3(new_n853), .ZN(new_n1060));
  NAND4_X1  g874(.A1(new_n1060), .A2(new_n847), .A3(new_n704), .A4(new_n761), .ZN(new_n1061));
  NAND3_X1  g875(.A1(new_n1056), .A2(new_n1043), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g876(.A(new_n1040), .ZN(new_n1063));
  AOI21_X1  g877(.A(G953), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g878(.A(new_n1042), .B1(new_n1053), .B2(new_n1064), .ZN(G72));
  NAND2_X1  g879(.A1(G472), .A2(G902), .ZN(new_n1066));
  XOR2_X1   g880(.A(new_n1066), .B(KEYINPUT63), .Z(new_n1067));
  INV_X1    g881(.A(new_n1067), .ZN(new_n1068));
  INV_X1    g882(.A(new_n474), .ZN(new_n1069));
  OR2_X1    g883(.A1(new_n1069), .A2(KEYINPUT127), .ZN(new_n1070));
  AOI21_X1  g884(.A(new_n774), .B1(new_n1069), .B2(KEYINPUT127), .ZN(new_n1071));
  AOI21_X1  g885(.A(new_n1068), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g886(.A(new_n976), .B1(new_n965), .B2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g887(.A1(new_n1056), .A2(new_n1043), .A3(new_n951), .A4(new_n1061), .ZN(new_n1074));
  AND2_X1   g888(.A1(new_n1074), .A2(new_n1067), .ZN(new_n1075));
  INV_X1    g889(.A(new_n473), .ZN(new_n1076));
  OAI21_X1  g890(.A(new_n459), .B1(new_n1076), .B2(new_n439), .ZN(new_n1077));
  OAI21_X1  g891(.A(new_n1073), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g892(.A1(new_n473), .A2(new_n440), .A3(new_n460), .ZN(new_n1079));
  NAND3_X1  g893(.A1(new_n1049), .A2(new_n1052), .A3(new_n951), .ZN(new_n1080));
  AOI21_X1  g894(.A(new_n1079), .B1(new_n1080), .B2(new_n1067), .ZN(new_n1081));
  NOR2_X1   g895(.A1(new_n1078), .A2(new_n1081), .ZN(G57));
endmodule


