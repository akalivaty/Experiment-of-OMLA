//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n555, new_n556, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n615, new_n617, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1124,
    new_n1125, new_n1126, new_n1128;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT67), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OR2_X1    g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n463), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n469), .A2(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n463), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n472), .A2(new_n475), .ZN(G160));
  NOR2_X1   g051(.A1(new_n467), .A2(new_n468), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(new_n463), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n477), .A2(G2105), .ZN(new_n479));
  AOI22_X1  g054(.A1(G124), .A2(new_n478), .B1(new_n479), .B2(G136), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G112), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT68), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n487), .B1(new_n470), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n479), .A2(KEYINPUT4), .A3(G138), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n478), .A2(G126), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n489), .A2(new_n490), .A3(new_n491), .A4(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  NAND2_X1  g070(.A1(KEYINPUT70), .A2(G543), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n504), .B1(new_n502), .B2(KEYINPUT69), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT6), .A3(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(G50), .A3(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n500), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n503), .A2(new_n512), .ZN(G303));
  INV_X1    g088(.A(G303), .ZN(G166));
  AND3_X1   g089(.A1(new_n506), .A2(KEYINPUT6), .A3(G651), .ZN(new_n515));
  AOI21_X1  g090(.A(KEYINPUT6), .B1(new_n506), .B2(G651), .ZN(new_n516));
  OAI21_X1  g091(.A(KEYINPUT71), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n505), .A2(new_n518), .A3(new_n507), .ZN(new_n519));
  AND3_X1   g094(.A1(new_n517), .A2(G543), .A3(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n520), .A2(G51), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n500), .ZN(new_n526));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI221_X1 g103(.A(new_n525), .B1(new_n526), .B2(new_n527), .C1(new_n510), .C2(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(KEYINPUT72), .B1(new_n521), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  NOR3_X1   g106(.A1(new_n521), .A2(KEYINPUT72), .A3(new_n529), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND2_X1  g109(.A1(new_n520), .A2(G52), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n500), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(new_n502), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n508), .A2(new_n500), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G90), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n535), .A2(new_n537), .A3(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n526), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(KEYINPUT73), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n546), .B(new_n542), .C1(new_n526), .C2(new_n543), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n545), .A2(new_n547), .A3(G651), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n520), .A2(G43), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n538), .A2(G81), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  AND3_X1   g132(.A1(new_n508), .A2(new_n500), .A3(G91), .ZN(new_n558));
  AND3_X1   g133(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n559));
  AOI21_X1  g134(.A(KEYINPUT5), .B1(KEYINPUT70), .B2(G543), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n561));
  NOR3_X1   g136(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(KEYINPUT74), .B1(new_n498), .B2(new_n499), .ZN(new_n563));
  OAI21_X1  g138(.A(G65), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n558), .B1(new_n566), .B2(G651), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n517), .A2(G53), .A3(G543), .A4(new_n519), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n570));
  INV_X1    g145(.A(G543), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(new_n508), .B2(KEYINPUT71), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT9), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n572), .A2(new_n573), .A3(G53), .A4(new_n519), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  AND3_X1   g150(.A1(new_n567), .A2(new_n568), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n568), .B1(new_n567), .B2(new_n575), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(G299));
  NAND2_X1  g153(.A1(new_n520), .A2(G49), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT76), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n500), .A2(G74), .ZN(new_n581));
  AOI22_X1  g156(.A1(G651), .A2(new_n581), .B1(new_n538), .B2(G87), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(G288));
  AOI22_X1  g158(.A1(new_n500), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n502), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n508), .A2(G48), .A3(G543), .ZN(new_n586));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n510), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(new_n520), .A2(G47), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n538), .A2(G85), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n591), .B(new_n592), .C1(new_n502), .C2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n538), .A2(G92), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n561), .B1(new_n559), .B2(new_n560), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n498), .A2(KEYINPUT74), .A3(new_n499), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(G651), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n572), .A2(G54), .A3(new_n519), .ZN(new_n606));
  AND3_X1   g181(.A1(new_n605), .A2(KEYINPUT77), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(KEYINPUT77), .B1(new_n605), .B2(new_n606), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n598), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n595), .B1(new_n610), .B2(G868), .ZN(G284));
  OAI21_X1  g186(.A(new_n595), .B1(new_n610), .B2(G868), .ZN(G321));
  MUX2_X1   g187(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g188(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n610), .B1(new_n615), .B2(G860), .ZN(G148));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n551), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n609), .A2(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n617), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n479), .A2(G135), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n478), .A2(G123), .ZN(new_n623));
  OR2_X1    g198(.A1(G99), .A2(G2105), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n624), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n622), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2096), .Z(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT78), .B(KEYINPUT12), .ZN(new_n628));
  NOR3_X1   g203(.A1(new_n465), .A2(new_n466), .A3(G2105), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n627), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT79), .ZN(G156));
  XOR2_X1   g211(.A(KEYINPUT15), .B(G2435), .Z(new_n637));
  XOR2_X1   g212(.A(KEYINPUT81), .B(G2438), .Z(new_n638));
  XOR2_X1   g213(.A(new_n637), .B(new_n638), .Z(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2430), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND3_X1   g216(.A1(new_n641), .A2(KEYINPUT82), .A3(KEYINPUT14), .ZN(new_n642));
  AOI21_X1  g217(.A(KEYINPUT82), .B1(new_n641), .B2(KEYINPUT14), .ZN(new_n643));
  OAI22_X1  g218(.A1(new_n642), .A2(new_n643), .B1(new_n640), .B2(new_n639), .ZN(new_n644));
  XOR2_X1   g219(.A(G1341), .B(G1348), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2451), .B(G2454), .Z(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  AND2_X1   g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(G14), .B1(new_n650), .B2(new_n652), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT17), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n660), .B2(new_n657), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n661), .B1(KEYINPUT83), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(KEYINPUT83), .B2(new_n663), .ZN(new_n665));
  INV_X1    g240(.A(new_n657), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n666), .A2(new_n662), .A3(new_n659), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT18), .Z(new_n668));
  NAND3_X1  g243(.A1(new_n658), .A2(new_n662), .A3(new_n660), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n665), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2096), .B(G2100), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(KEYINPUT84), .B(KEYINPUT19), .Z(new_n673));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(new_n678), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT20), .Z(new_n682));
  NAND2_X1  g257(.A1(new_n675), .A2(new_n679), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(KEYINPUT85), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(KEYINPUT85), .ZN(new_n685));
  AOI211_X1 g260(.A(new_n680), .B(new_n682), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT86), .ZN(new_n687));
  XOR2_X1   g262(.A(G1981), .B(G1986), .Z(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n687), .B(new_n692), .ZN(G229));
  INV_X1    g268(.A(G29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G25), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n478), .A2(G119), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT87), .ZN(new_n697));
  OAI21_X1  g272(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n698));
  INV_X1    g273(.A(G107), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(G2105), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n479), .A2(G131), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NOR3_X1   g277(.A1(new_n697), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n695), .B1(new_n703), .B2(new_n694), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT88), .Z(new_n705));
  XOR2_X1   g280(.A(KEYINPUT35), .B(G1991), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G23), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n580), .A2(new_n582), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n708), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT33), .B(G1976), .Z(new_n712));
  OR2_X1    g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n708), .A2(G22), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G166), .B2(new_n708), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(G1971), .Z(new_n717));
  NOR2_X1   g292(.A1(G6), .A2(G16), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n589), .B2(G16), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT32), .B(G1981), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n713), .A2(new_n714), .A3(new_n717), .A4(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n722), .A2(KEYINPUT34), .ZN(new_n723));
  AND3_X1   g298(.A1(new_n708), .A2(KEYINPUT89), .A3(G24), .ZN(new_n724));
  AOI21_X1  g299(.A(KEYINPUT89), .B1(new_n708), .B2(G24), .ZN(new_n725));
  AOI211_X1 g300(.A(new_n724), .B(new_n725), .C1(G290), .C2(G16), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n727), .A2(G1986), .B1(KEYINPUT90), .B2(KEYINPUT36), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G1986), .B2(new_n727), .ZN(new_n729));
  NOR3_X1   g304(.A1(new_n707), .A2(new_n723), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n722), .A2(KEYINPUT34), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n694), .A2(G35), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G162), .B2(new_n694), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G2090), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT100), .B(KEYINPUT29), .Z(new_n738));
  XOR2_X1   g313(.A(new_n737), .B(new_n738), .Z(new_n739));
  NOR2_X1   g314(.A1(G16), .A2(G19), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n552), .B2(G16), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G1341), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G16), .A2(G21), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G168), .B2(G16), .ZN(new_n745));
  INV_X1    g320(.A(G1966), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT92), .Z(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(KEYINPUT91), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(KEYINPUT91), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT25), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n750), .A2(KEYINPUT25), .A3(new_n751), .ZN(new_n755));
  NAND2_X1  g330(.A1(G115), .A2(G2104), .ZN(new_n756));
  INV_X1    g331(.A(G127), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n477), .B2(new_n757), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n758), .A2(G2105), .B1(new_n479), .B2(G139), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n754), .A2(new_n755), .A3(new_n759), .ZN(new_n760));
  MUX2_X1   g335(.A(G33), .B(new_n760), .S(G29), .Z(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT93), .Z(new_n762));
  OAI211_X1 g337(.A(new_n743), .B(new_n747), .C1(G2072), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n708), .A2(G5), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G171), .B2(new_n708), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT98), .Z(new_n766));
  NOR2_X1   g341(.A1(new_n766), .A2(G1961), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT24), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n694), .B1(new_n768), .B2(G34), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n768), .B2(G34), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G160), .B2(G29), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(G2084), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT31), .B(G11), .Z(new_n773));
  INV_X1    g348(.A(G28), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n774), .A2(KEYINPUT30), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT97), .ZN(new_n776));
  AOI21_X1  g351(.A(G29), .B1(new_n774), .B2(KEYINPUT30), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n773), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n772), .B(new_n778), .C1(new_n694), .C2(new_n626), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n694), .A2(G26), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT28), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n479), .A2(G140), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n478), .A2(G128), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n463), .A2(G116), .ZN(new_n784));
  OAI21_X1  g359(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n782), .B(new_n783), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n781), .B1(new_n786), .B2(G29), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G2067), .ZN(new_n788));
  NAND3_X1  g363(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT96), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT26), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n478), .A2(G129), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT95), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n479), .A2(G141), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND3_X1   g372(.A1(new_n791), .A2(new_n792), .A3(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(new_n694), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n694), .B2(G32), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT27), .B(G1996), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n788), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AOI211_X1 g377(.A(new_n779), .B(new_n802), .C1(new_n800), .C2(new_n801), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n766), .A2(G1961), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n771), .A2(G2084), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT99), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n694), .A2(G27), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G164), .B2(new_n694), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G2078), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n803), .A2(new_n804), .A3(new_n810), .ZN(new_n811));
  OR3_X1    g386(.A1(new_n763), .A2(new_n767), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n762), .A2(G2072), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT94), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n708), .A2(G4), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n610), .B2(new_n708), .ZN(new_n816));
  INV_X1    g391(.A(G1348), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n708), .A2(G20), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT23), .ZN(new_n820));
  INV_X1    g395(.A(G299), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(new_n708), .ZN(new_n822));
  INV_X1    g397(.A(G1956), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n814), .A2(new_n818), .A3(new_n824), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n734), .A2(new_n812), .A3(new_n825), .ZN(G311));
  INV_X1    g401(.A(new_n734), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n825), .A2(new_n812), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(G150));
  NOR2_X1   g404(.A1(new_n609), .A2(new_n615), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT38), .ZN(new_n831));
  NAND2_X1  g406(.A1(G80), .A2(G543), .ZN(new_n832));
  INV_X1    g407(.A(G67), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n526), .B2(new_n833), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n834), .A2(G651), .B1(new_n538), .B2(G93), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n520), .A2(G55), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n551), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n551), .A2(new_n837), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n831), .B(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT101), .B(G860), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n844), .B1(new_n835), .B2(new_n836), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT37), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(G145));
  XNOR2_X1  g423(.A(new_n494), .B(new_n786), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n760), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(new_n798), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n478), .A2(G130), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n463), .A2(G118), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(G142), .B2(new_n479), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(new_n630), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n703), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT103), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n851), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(G160), .B(KEYINPUT102), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n485), .B(new_n626), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G37), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n851), .A2(new_n858), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(new_n864), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n851), .A2(new_n858), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT40), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(G395));
  XNOR2_X1  g448(.A(G288), .B(G305), .ZN(new_n874));
  XNOR2_X1  g449(.A(G290), .B(G303), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT42), .ZN(new_n877));
  INV_X1    g452(.A(new_n875), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n874), .B(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT42), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n840), .B(new_n619), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n609), .B1(new_n576), .B2(new_n577), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(G299), .A2(new_n610), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n609), .B(KEYINPUT104), .C1(new_n576), .C2(new_n577), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n883), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n892), .B1(G299), .B2(new_n610), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(new_n886), .A3(new_n888), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT105), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n889), .A2(new_n892), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n893), .A2(new_n886), .A3(KEYINPUT105), .A4(new_n888), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n883), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n882), .A2(new_n891), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n882), .B1(new_n891), .B2(new_n900), .ZN(new_n902));
  OAI21_X1  g477(.A(G868), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n837), .A2(new_n617), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(G295));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n903), .A2(new_n906), .A3(new_n904), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n906), .B1(new_n903), .B2(new_n904), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(G331));
  XOR2_X1   g484(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n910));
  NOR3_X1   g485(.A1(new_n531), .A2(G171), .A3(new_n532), .ZN(new_n911));
  INV_X1    g486(.A(new_n532), .ZN(new_n912));
  AOI21_X1  g487(.A(G301), .B1(new_n912), .B2(new_n530), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n840), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(G171), .B1(new_n531), .B2(new_n532), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n912), .A2(new_n530), .A3(G301), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n915), .A2(new_n916), .A3(new_n839), .A4(new_n838), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n894), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n920), .B1(new_n897), .B2(KEYINPUT109), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n889), .A2(new_n922), .A3(new_n892), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n919), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n890), .A2(new_n918), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n879), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n925), .B1(new_n899), .B2(new_n918), .ZN(new_n927));
  AOI21_X1  g502(.A(G37), .B1(new_n927), .B2(new_n876), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI22_X1  g505(.A1(new_n895), .A2(new_n894), .B1(new_n889), .B2(new_n892), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n919), .B1(new_n931), .B2(new_n898), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n879), .B1(new_n932), .B2(new_n925), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n929), .B1(new_n928), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n930), .B1(new_n934), .B2(KEYINPUT108), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n936));
  AOI211_X1 g511(.A(new_n936), .B(new_n929), .C1(new_n928), .C2(new_n933), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n910), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n928), .A2(new_n929), .A3(new_n933), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n926), .A2(new_n928), .ZN(new_n940));
  OAI211_X1 g515(.A(KEYINPUT44), .B(new_n939), .C1(new_n940), .C2(new_n929), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(new_n941), .ZN(G397));
  INV_X1    g517(.A(G1384), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n494), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT45), .B1(new_n944), .B2(KEYINPUT110), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(KEYINPUT110), .B2(new_n944), .ZN(new_n946));
  NAND2_X1  g521(.A1(G160), .A2(G40), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G2067), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n786), .B(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n798), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g527(.A(new_n952), .B(KEYINPUT126), .Z(new_n953));
  INV_X1    g528(.A(G1996), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n948), .A2(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n955), .B(KEYINPUT46), .Z(new_n956));
  NOR2_X1   g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT47), .ZN(new_n958));
  INV_X1    g533(.A(new_n948), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n703), .B(new_n706), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n798), .B(G1996), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n950), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  OR3_X1    g539(.A1(new_n959), .A2(G1986), .A3(G290), .ZN(new_n965));
  XNOR2_X1  g540(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(new_n965), .B2(new_n966), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n703), .A2(new_n706), .ZN(new_n969));
  OAI22_X1  g544(.A1(new_n962), .A2(new_n969), .B1(G2067), .B2(new_n786), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n948), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n958), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n947), .B1(new_n974), .B2(new_n944), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n494), .A2(new_n943), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT45), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n944), .A2(KEYINPUT50), .ZN(new_n980));
  INV_X1    g555(.A(new_n947), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n494), .A2(new_n982), .A3(new_n943), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n980), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  OAI22_X1  g559(.A1(new_n979), .A2(G1971), .B1(G2090), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(G8), .ZN(new_n986));
  NAND2_X1  g561(.A1(G303), .A2(G8), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT55), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n944), .A2(new_n947), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n991), .A2(KEYINPUT111), .A3(G8), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n993));
  INV_X1    g568(.A(G8), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n993), .B1(new_n990), .B2(new_n994), .ZN(new_n995));
  AOI22_X1  g570(.A1(new_n992), .A2(new_n995), .B1(G1976), .B2(new_n710), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT52), .ZN(new_n998));
  INV_X1    g573(.A(G1976), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT52), .B1(G288), .B2(new_n999), .ZN(new_n1000));
  OR2_X1    g575(.A1(G305), .A2(G1981), .ZN(new_n1001));
  NAND2_X1  g576(.A1(G305), .A2(G1981), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n1003), .B(KEYINPUT49), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n992), .A2(new_n995), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n996), .A2(new_n1000), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n988), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n985), .A2(G8), .A3(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n989), .A2(new_n998), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n978), .A2(KEYINPUT112), .A3(new_n746), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n980), .A2(new_n981), .A3(new_n983), .ZN(new_n1011));
  INV_X1    g586(.A(G2084), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1966), .B1(new_n975), .B2(new_n977), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(KEYINPUT112), .ZN(new_n1016));
  OAI21_X1  g591(.A(G8), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(G286), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1009), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(KEYINPUT113), .A2(KEYINPUT63), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n998), .A2(new_n1006), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1008), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n710), .A2(new_n999), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1001), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n1023), .A2(new_n1024), .B1(new_n1005), .B2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g603(.A(KEYINPUT113), .B(KEYINPUT63), .Z(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(new_n1009), .B2(new_n1019), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1022), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(G286), .A2(G8), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1017), .A2(KEYINPUT51), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n979), .B2(G1966), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1015), .A2(KEYINPUT112), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1034), .B(G8), .C1(new_n1038), .C2(G286), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT122), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1032), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1040), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1042));
  AOI211_X1 g617(.A(KEYINPUT122), .B(new_n1032), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1033), .B(new_n1039), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G2078), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n979), .A2(KEYINPUT53), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(new_n978), .B2(G2078), .ZN(new_n1048));
  INV_X1    g623(.A(G1961), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n984), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1046), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(G171), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1052), .A2(KEYINPUT62), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1044), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n984), .A2(new_n823), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n567), .A2(new_n575), .ZN(new_n1056));
  XOR2_X1   g631(.A(new_n1056), .B(KEYINPUT57), .Z(new_n1057));
  XOR2_X1   g632(.A(KEYINPUT56), .B(G2072), .Z(new_n1058));
  XNOR2_X1  g633(.A(new_n1058), .B(KEYINPUT114), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n975), .A2(new_n977), .A3(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1055), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n984), .A2(new_n817), .B1(new_n949), .B2(new_n990), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(new_n609), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1057), .B1(new_n1055), .B2(new_n1060), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1061), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1065), .B(new_n1066), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n610), .A2(KEYINPUT121), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n610), .A2(KEYINPUT121), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1062), .A2(KEYINPUT60), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1062), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT60), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1070), .B(new_n1073), .C1(new_n1074), .C2(new_n1068), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT61), .B1(new_n1064), .B2(KEYINPUT120), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1055), .A2(new_n1060), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1057), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n1061), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1076), .A2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1079), .A2(new_n1061), .A3(KEYINPUT120), .A4(KEYINPUT61), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1075), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n979), .A2(new_n1084), .A3(new_n954), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT116), .B1(new_n978), .B2(G1996), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT58), .B(G1341), .Z(new_n1087));
  NAND2_X1  g662(.A1(new_n991), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT117), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n991), .A2(new_n1090), .A3(new_n1087), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1085), .A2(new_n1086), .A3(new_n1089), .A4(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT119), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n551), .B1(new_n1095), .B2(KEYINPUT59), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1092), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1094), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1067), .B1(new_n1083), .B2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT123), .B(G2078), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n947), .A2(new_n1047), .A3(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n946), .A2(new_n977), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1048), .A2(new_n1103), .A3(new_n1050), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT125), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1104), .A2(new_n1105), .A3(G171), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1105), .B1(new_n1104), .B2(G171), .ZN(new_n1107));
  OAI221_X1 g682(.A(KEYINPUT54), .B1(G171), .B2(new_n1051), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT124), .B1(new_n1104), .B2(G171), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n1052), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1104), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1109), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1108), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1054), .B1(new_n1100), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1044), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1051), .A2(KEYINPUT62), .A3(G171), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1009), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1031), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  XOR2_X1   g694(.A(G290), .B(G1986), .Z(new_n1120));
  AOI21_X1  g695(.A(new_n959), .B1(new_n963), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n973), .B1(new_n1119), .B2(new_n1121), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g697(.A1(new_n935), .A2(new_n937), .ZN(new_n1124));
  NOR3_X1   g698(.A1(G229), .A2(new_n461), .A3(G227), .ZN(new_n1125));
  OAI211_X1 g699(.A(new_n655), .B(new_n1125), .C1(new_n865), .C2(new_n870), .ZN(new_n1126));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1126), .ZN(G308));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1128));
  OAI21_X1  g702(.A(new_n1128), .B1(new_n937), .B2(new_n935), .ZN(G225));
endmodule


