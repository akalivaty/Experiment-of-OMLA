//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 1 0 1 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n215));
  XNOR2_X1  g0015(.A(new_n214), .B(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G97), .ZN(new_n219));
  INV_X1    g0019(.A(G257), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n217), .B1(new_n201), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n212), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(new_n210), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n206), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n216), .B(new_n226), .C1(new_n228), .C2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(new_n218), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G68), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT66), .B(G50), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  XNOR2_X1  g0047(.A(KEYINPUT3), .B(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n248), .A2(G232), .A3(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G107), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n248), .A2(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(G238), .ZN(new_n253));
  OAI221_X1 g0053(.A(new_n250), .B1(new_n251), .B2(new_n248), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G41), .ZN(new_n257));
  INV_X1    g0057(.A(G45), .ZN(new_n258));
  AOI21_X1  g0058(.A(G1), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G1), .A3(G13), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n259), .A2(new_n261), .A3(G274), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n263), .B1(G244), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n256), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G169), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n227), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT15), .B(G87), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n274), .B(KEYINPUT69), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(new_n210), .A3(G33), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n278), .A2(new_n279), .B1(G20), .B2(G77), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n273), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(new_n272), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT68), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n285), .B1(new_n210), .B2(G1), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n209), .A2(KEYINPUT68), .A3(G20), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n284), .A2(G77), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n289), .B1(G77), .B2(new_n282), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n270), .B1(G179), .B2(new_n268), .C1(new_n281), .C2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G200), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n292), .B1(new_n256), .B2(new_n267), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n281), .A2(new_n290), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n294), .B1(new_n295), .B2(new_n268), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n291), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT70), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT17), .ZN(new_n299));
  AND2_X1   g0099(.A1(KEYINPUT3), .A2(G33), .ZN(new_n300));
  NOR2_X1   g0100(.A1(KEYINPUT3), .A2(G33), .ZN(new_n301));
  OAI211_X1 g0101(.A(G226), .B(G1698), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G223), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(G1698), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(new_n300), .B2(new_n301), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G87), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT78), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(KEYINPUT78), .A2(G33), .A3(G87), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n302), .A2(new_n305), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n255), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT79), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n311), .A2(KEYINPUT79), .A3(new_n255), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n262), .B(new_n295), .C1(new_n218), .C2(new_n265), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n314), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT80), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n311), .A2(new_n255), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n262), .B1(new_n218), .B2(new_n265), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n292), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n318), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n319), .B1(new_n318), .B2(new_n322), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n284), .A2(new_n278), .A3(new_n288), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n277), .A2(new_n283), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n326), .A2(KEYINPUT77), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT77), .B1(new_n326), .B2(new_n327), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT3), .ZN(new_n331));
  INV_X1    g0131(.A(G33), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(KEYINPUT3), .A2(G33), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(new_n210), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT76), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n300), .A2(new_n301), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n339), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n336), .B1(new_n335), .B2(new_n337), .ZN(new_n342));
  OAI21_X1  g0142(.A(G68), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n203), .B(new_n205), .C1(new_n201), .C2(new_n202), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(G20), .B1(G159), .B2(new_n279), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT16), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  XOR2_X1   g0146(.A(KEYINPUT75), .B(KEYINPUT7), .Z(new_n347));
  NOR2_X1   g0147(.A1(new_n347), .A2(new_n335), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n300), .A2(new_n301), .A3(G20), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT7), .ZN(new_n350));
  OAI21_X1  g0150(.A(G68), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n345), .B(KEYINPUT16), .C1(new_n348), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n272), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n330), .B1(new_n346), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n299), .B1(new_n325), .B2(new_n354), .ZN(new_n355));
  AND3_X1   g0155(.A1(new_n311), .A2(KEYINPUT79), .A3(new_n255), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT79), .B1(new_n311), .B2(new_n255), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n321), .A2(G179), .ZN(new_n359));
  INV_X1    g0159(.A(new_n321), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n312), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n358), .A2(new_n359), .B1(new_n361), .B2(new_n269), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n354), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT18), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT18), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n354), .A2(new_n365), .A3(new_n362), .ZN(new_n366));
  NOR3_X1   g0166(.A1(new_n356), .A2(new_n357), .A3(new_n316), .ZN(new_n367));
  AOI21_X1  g0167(.A(G200), .B1(new_n360), .B2(new_n312), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT80), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n318), .A2(new_n322), .A3(new_n319), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n354), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT17), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n355), .A2(new_n364), .A3(new_n366), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n283), .A2(new_n202), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT12), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n284), .A2(G68), .A3(new_n288), .ZN(new_n377));
  INV_X1    g0177(.A(new_n279), .ZN(new_n378));
  INV_X1    g0178(.A(G50), .ZN(new_n379));
  OAI22_X1  g0179(.A1(new_n378), .A2(new_n379), .B1(new_n210), .B2(G68), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n210), .A2(G33), .ZN(new_n381));
  INV_X1    g0181(.A(G77), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n272), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT11), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n376), .B(new_n377), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n384), .A2(new_n385), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT14), .ZN(new_n390));
  OAI211_X1 g0190(.A(G232), .B(G1698), .C1(new_n300), .C2(new_n301), .ZN(new_n391));
  OAI211_X1 g0191(.A(G226), .B(new_n249), .C1(new_n300), .C2(new_n301), .ZN(new_n392));
  AND3_X1   g0192(.A1(KEYINPUT74), .A2(G33), .A3(G97), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT74), .B1(G33), .B2(G97), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n391), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n255), .ZN(new_n397));
  INV_X1    g0197(.A(G274), .ZN(new_n398));
  INV_X1    g0198(.A(new_n227), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n398), .B1(new_n399), .B2(new_n260), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n266), .A2(G238), .B1(new_n400), .B2(new_n259), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT13), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n397), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n402), .B1(new_n397), .B2(new_n401), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n390), .B(G169), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(G179), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n397), .A2(new_n401), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT13), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n397), .A2(new_n401), .A3(new_n402), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n405), .B1(new_n406), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n390), .B1(new_n410), .B2(G169), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n389), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n410), .A2(G200), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n414), .B(new_n388), .C1(new_n295), .C2(new_n410), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OR3_X1    g0216(.A1(new_n298), .A2(new_n374), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT72), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n248), .A2(G222), .A3(new_n249), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n419), .B1(new_n382), .B2(new_n248), .C1(new_n252), .C2(new_n303), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n255), .ZN(new_n421));
  XNOR2_X1  g0221(.A(KEYINPUT67), .B(G226), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n263), .B1(new_n266), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n418), .B1(new_n425), .B2(new_n292), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(KEYINPUT72), .A3(G200), .ZN(new_n427));
  OR3_X1    g0227(.A1(new_n424), .A2(KEYINPUT73), .A3(new_n295), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT73), .B1(new_n424), .B2(new_n295), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n426), .A2(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT10), .B1(new_n430), .B2(KEYINPUT71), .ZN(new_n431));
  OAI21_X1  g0231(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n432));
  INV_X1    g0232(.A(G150), .ZN(new_n433));
  OAI221_X1 g0233(.A(new_n432), .B1(new_n433), .B2(new_n378), .C1(new_n381), .C2(new_n277), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n272), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n379), .B1(new_n286), .B2(new_n287), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n284), .A2(new_n436), .B1(new_n379), .B2(new_n283), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n438), .B(KEYINPUT9), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n430), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n431), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n430), .B(new_n439), .C1(KEYINPUT71), .C2(KEYINPUT10), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n435), .A2(new_n437), .B1(new_n424), .B2(new_n269), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(G179), .B2(new_n424), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n417), .A2(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(G264), .B(G1698), .C1(new_n300), .C2(new_n301), .ZN(new_n447));
  OAI211_X1 g0247(.A(G257), .B(new_n249), .C1(new_n300), .C2(new_n301), .ZN(new_n448));
  INV_X1    g0248(.A(G303), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n447), .B(new_n448), .C1(new_n449), .C2(new_n248), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n255), .ZN(new_n451));
  XNOR2_X1  g0251(.A(KEYINPUT5), .B(G41), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n258), .A2(G1), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n452), .A2(new_n453), .B1(new_n399), .B2(new_n260), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n209), .A2(G45), .ZN(new_n455));
  NOR2_X1   g0255(.A1(KEYINPUT5), .A2(G41), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(KEYINPUT5), .A2(G41), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n455), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n454), .A2(G270), .B1(new_n400), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n451), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT20), .ZN(new_n462));
  AOI21_X1  g0262(.A(G20), .B1(G33), .B2(G283), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n332), .A2(G97), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT86), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(G116), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n271), .A2(new_n227), .B1(G20), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n465), .B1(new_n463), .B2(new_n464), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n462), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n463), .A2(new_n464), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT86), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n473), .A2(KEYINPUT20), .A3(new_n466), .A4(new_n468), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT87), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n332), .A2(G1), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n283), .A2(new_n272), .A3(new_n477), .ZN(new_n478));
  OR3_X1    g0278(.A1(new_n282), .A2(KEYINPUT85), .A3(G116), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT85), .B1(new_n282), .B2(G116), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n478), .A2(G116), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n475), .A2(new_n476), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n476), .B1(new_n475), .B2(new_n481), .ZN(new_n483));
  OAI211_X1 g0283(.A(G169), .B(new_n461), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT88), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT21), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n461), .A2(G169), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n475), .A2(new_n481), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT87), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n475), .A2(new_n476), .A3(new_n481), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(KEYINPUT21), .B1(new_n492), .B2(KEYINPUT88), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n482), .A2(new_n483), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n451), .A2(new_n460), .A3(G179), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n461), .A2(G200), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n494), .B(new_n498), .C1(new_n295), .C2(new_n461), .ZN(new_n499));
  AND4_X1   g0299(.A1(new_n487), .A2(new_n493), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n282), .A2(G97), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n501), .B1(new_n478), .B2(G97), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(G107), .B1(new_n341), .B2(new_n342), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n279), .A2(KEYINPUT81), .A3(G77), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT81), .B1(new_n279), .B2(G77), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT6), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n508), .A2(new_n219), .A3(G107), .ZN(new_n509));
  XNOR2_X1  g0309(.A(G97), .B(G107), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n509), .B1(new_n510), .B2(new_n508), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n507), .B1(new_n511), .B2(new_n210), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n504), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n503), .B1(new_n514), .B2(new_n272), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n459), .A2(new_n220), .A3(new_n255), .ZN(new_n516));
  OAI211_X1 g0316(.A(G244), .B(new_n249), .C1(new_n300), .C2(new_n301), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT4), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n248), .A2(KEYINPUT4), .A3(G244), .A4(new_n249), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G283), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n248), .A2(G250), .A3(G1698), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n519), .A2(new_n520), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n516), .B1(new_n523), .B2(new_n255), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n459), .A2(new_n400), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n524), .A2(new_n295), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(G200), .B1(new_n524), .B2(new_n525), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n515), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT76), .B1(new_n349), .B2(new_n347), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(new_n340), .A3(new_n338), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n512), .B1(new_n530), .B2(G107), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n502), .B1(new_n531), .B2(new_n273), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n523), .A2(new_n255), .ZN(new_n533));
  INV_X1    g0333(.A(new_n516), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n533), .A2(new_n525), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n269), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n524), .A2(new_n406), .A3(new_n525), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n532), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n528), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT83), .ZN(new_n540));
  NOR3_X1   g0340(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n541));
  OAI21_X1  g0341(.A(KEYINPUT19), .B1(new_n393), .B2(new_n394), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n541), .B1(new_n542), .B2(new_n210), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n210), .B(G68), .C1(new_n300), .C2(new_n301), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n210), .A2(G33), .A3(G97), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT19), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n540), .B1(new_n543), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n541), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G97), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT74), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(KEYINPUT74), .A2(G33), .A3(G97), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n546), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n550), .B1(new_n555), .B2(G20), .ZN(new_n556));
  AOI21_X1  g0356(.A(G20), .B1(new_n333), .B2(new_n334), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n557), .A2(G68), .B1(new_n546), .B2(new_n545), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n558), .A3(KEYINPUT83), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n549), .A2(new_n559), .A3(new_n272), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n275), .A2(new_n478), .ZN(new_n561));
  INV_X1    g0361(.A(new_n275), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n283), .ZN(new_n563));
  AND3_X1   g0363(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n261), .A2(G250), .A3(new_n455), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n261), .A2(G274), .A3(new_n453), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT82), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n261), .A2(KEYINPUT82), .A3(G274), .A4(new_n453), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n565), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(G244), .B(G1698), .C1(new_n300), .C2(new_n301), .ZN(new_n571));
  OAI211_X1 g0371(.A(G238), .B(new_n249), .C1(new_n300), .C2(new_n301), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G33), .A2(G116), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n255), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n570), .A2(new_n406), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n570), .A2(new_n575), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n576), .B1(new_n578), .B2(G169), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n570), .A2(new_n295), .A3(new_n575), .ZN(new_n580));
  AOI21_X1  g0380(.A(G200), .B1(new_n570), .B2(new_n575), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n478), .A2(G87), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n560), .A2(new_n563), .A3(new_n583), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n564), .A2(new_n579), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  OR3_X1    g0385(.A1(new_n539), .A2(KEYINPUT84), .A3(new_n585), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n454), .A2(G264), .B1(new_n400), .B2(new_n459), .ZN(new_n587));
  OAI211_X1 g0387(.A(G257), .B(G1698), .C1(new_n300), .C2(new_n301), .ZN(new_n588));
  OAI211_X1 g0388(.A(G250), .B(new_n249), .C1(new_n300), .C2(new_n301), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G33), .A2(G294), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n255), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n587), .A2(KEYINPUT89), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT89), .B1(new_n587), .B2(new_n592), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n295), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n587), .A2(new_n592), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n292), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n251), .A2(KEYINPUT23), .A3(G20), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT23), .B1(new_n251), .B2(G20), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n599), .A2(new_n600), .B1(G20), .B2(new_n573), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n210), .B(G87), .C1(new_n300), .C2(new_n301), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT22), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT22), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n248), .A2(new_n604), .A3(new_n210), .A4(G87), .ZN(new_n605));
  AOI211_X1 g0405(.A(KEYINPUT24), .B(new_n601), .C1(new_n603), .C2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT24), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n603), .A2(new_n605), .ZN(new_n608));
  INV_X1    g0408(.A(new_n601), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n272), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n282), .A2(G107), .ZN(new_n612));
  XOR2_X1   g0412(.A(new_n612), .B(KEYINPUT25), .Z(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(G107), .B2(new_n478), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n598), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n611), .A2(new_n614), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n593), .A2(new_n594), .A3(new_n269), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n587), .A2(new_n592), .A3(G179), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT90), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT90), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n587), .A2(new_n592), .A3(new_n621), .A4(G179), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n617), .B1(new_n618), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n616), .A2(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n560), .A2(new_n563), .A3(new_n583), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n577), .A2(new_n292), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(G190), .B2(new_n577), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n570), .A2(new_n406), .A3(new_n575), .ZN(new_n629));
  AOI21_X1  g0429(.A(G169), .B1(new_n570), .B2(new_n575), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n626), .A2(new_n628), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n633), .A2(new_n528), .A3(new_n538), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n625), .B1(new_n634), .B2(KEYINPUT84), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n446), .A2(new_n500), .A3(new_n586), .A4(new_n635), .ZN(new_n636));
  XOR2_X1   g0436(.A(new_n636), .B(KEYINPUT91), .Z(G372));
  INV_X1    g0437(.A(KEYINPUT94), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n617), .B(KEYINPUT93), .C1(new_n618), .C2(new_n623), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT89), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n591), .A2(new_n255), .ZN(new_n642));
  INV_X1    g0442(.A(new_n458), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n453), .B1(new_n643), .B2(new_n456), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n644), .A2(G264), .A3(new_n261), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n525), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n641), .B1(new_n642), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n587), .A2(new_n592), .A3(KEYINPUT89), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(G169), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n649), .A2(new_n620), .A3(new_n622), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT93), .B1(new_n650), .B2(new_n617), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n640), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n493), .A2(new_n487), .A3(new_n497), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n638), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT93), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n624), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n639), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n484), .A2(new_n485), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n658), .A2(KEYINPUT21), .B1(new_n495), .B2(new_n496), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n657), .A2(new_n659), .A3(KEYINPUT94), .A4(new_n487), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n617), .B1(new_n595), .B2(new_n597), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT92), .B1(new_n634), .B2(new_n661), .ZN(new_n662));
  NOR3_X1   g0462(.A1(new_n539), .A2(new_n661), .A3(new_n585), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT92), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n654), .A2(new_n660), .A3(new_n662), .A4(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n564), .A2(new_n579), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n585), .B2(new_n538), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n532), .A2(new_n536), .A3(new_n537), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n633), .A2(new_n670), .A3(KEYINPUT26), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n667), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n446), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n444), .ZN(new_n675));
  INV_X1    g0475(.A(new_n413), .ZN(new_n676));
  INV_X1    g0476(.A(new_n291), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n676), .B1(new_n415), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n355), .A2(new_n373), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n364), .B(new_n366), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n441), .A2(new_n442), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n675), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n674), .A2(new_n682), .ZN(G369));
  NAND3_X1  g0483(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G213), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n495), .A2(new_n689), .ZN(new_n690));
  MUX2_X1   g0490(.A(new_n653), .B(new_n500), .S(new_n690), .Z(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G330), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n625), .ZN(new_n694));
  INV_X1    g0494(.A(new_n689), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n694), .B1(new_n615), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n624), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n689), .B1(new_n659), .B2(new_n487), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n699), .A2(new_n694), .B1(new_n652), .B2(new_n695), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(G399));
  INV_X1    g0501(.A(new_n213), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G41), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n550), .A2(G116), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(G1), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n229), .B2(new_n704), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT95), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n673), .A2(new_n695), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n493), .A2(new_n487), .A3(new_n497), .A4(new_n624), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n663), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n672), .ZN(new_n715));
  AOI21_X1  g0515(.A(KEYINPUT98), .B1(new_n715), .B2(new_n695), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT98), .ZN(new_n717));
  AOI211_X1 g0517(.A(new_n717), .B(new_n689), .C1(new_n714), .C2(new_n672), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n712), .B1(new_n719), .B2(new_n711), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT97), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n635), .A2(new_n586), .A3(new_n500), .A4(new_n695), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n461), .A2(new_n577), .A3(new_n406), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n644), .A2(new_n255), .A3(new_n398), .ZN(new_n725));
  AOI211_X1 g0525(.A(new_n725), .B(new_n516), .C1(new_n523), .C2(new_n255), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n642), .A2(new_n646), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n726), .A2(KEYINPUT96), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT96), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n535), .B2(new_n596), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n724), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n496), .A2(new_n578), .A3(new_n727), .A4(new_n524), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n577), .A2(new_n596), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(KEYINPUT30), .A3(new_n496), .A4(new_n524), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n731), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT31), .B1(new_n737), .B2(new_n689), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n734), .A2(new_n736), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT96), .B1(new_n726), .B2(new_n727), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n535), .A2(new_n729), .A3(new_n596), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n723), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI211_X1 g0542(.A(KEYINPUT31), .B(new_n689), .C1(new_n739), .C2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n738), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n722), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n721), .B1(new_n746), .B2(G330), .ZN(new_n747));
  INV_X1    g0547(.A(G330), .ZN(new_n748));
  AOI211_X1 g0548(.A(KEYINPUT97), .B(new_n748), .C1(new_n722), .C2(new_n745), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n720), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n709), .B1(new_n753), .B2(G1), .ZN(G364));
  INV_X1    g0554(.A(G13), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n209), .B1(new_n756), .B2(G45), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n703), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n693), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(G330), .B2(new_n691), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n759), .B(KEYINPUT99), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n213), .A2(new_n248), .ZN(new_n763));
  INV_X1    g0563(.A(G355), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n763), .A2(new_n764), .B1(G116), .B2(new_n213), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n243), .A2(G45), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n702), .A2(new_n248), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n768), .B1(new_n230), .B2(new_n258), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n765), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n227), .B1(G20), .B2(new_n269), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n762), .B1(new_n770), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n406), .A2(new_n292), .A3(KEYINPUT101), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT101), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(G179), .B2(G200), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n295), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n210), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G294), .ZN(new_n784));
  NAND3_X1  g0584(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G190), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(KEYINPUT33), .B(G317), .Z(new_n788));
  NOR2_X1   g0588(.A1(new_n210), .A2(G179), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n789), .A2(G190), .A3(G200), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n787), .A2(new_n788), .B1(new_n790), .B2(new_n449), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n785), .A2(new_n295), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G326), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n789), .A2(new_n295), .A3(G200), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n793), .A2(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n791), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n406), .A2(G200), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n799), .A2(G20), .A3(G190), .ZN(new_n800));
  INV_X1    g0600(.A(G322), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n339), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n210), .A2(G190), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n799), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n802), .B1(G311), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n778), .A2(new_n780), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n803), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G329), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n784), .A2(new_n798), .A3(new_n806), .A4(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G159), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT32), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n783), .A2(G97), .ZN(new_n815));
  INV_X1    g0615(.A(G87), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n793), .A2(new_n379), .B1(new_n790), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G68), .B2(new_n786), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n814), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n800), .A2(new_n201), .B1(new_n804), .B2(new_n382), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n820), .A2(KEYINPUT100), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(KEYINPUT100), .ZN(new_n822));
  INV_X1    g0622(.A(new_n795), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n339), .B1(new_n823), .B2(G107), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n811), .B1(new_n819), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n777), .B1(new_n774), .B2(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT102), .Z(new_n828));
  XOR2_X1   g0628(.A(new_n773), .B(KEYINPUT103), .Z(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n691), .B2(new_n829), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n761), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(G396));
  NOR2_X1   g0632(.A1(new_n291), .A2(new_n689), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n296), .A2(new_n293), .B1(new_n294), .B2(new_n695), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n833), .B1(new_n291), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n710), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n689), .B1(new_n666), .B2(new_n672), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n835), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n751), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n841), .A2(KEYINPUT106), .ZN(new_n842));
  INV_X1    g0642(.A(new_n759), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(KEYINPUT106), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n750), .A2(new_n837), .A3(new_n839), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n842), .A2(new_n843), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n774), .A2(new_n771), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n762), .B1(G77), .B2(new_n848), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n793), .A2(new_n449), .B1(new_n795), .B2(new_n816), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n787), .A2(new_n796), .B1(new_n790), .B2(new_n251), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n809), .A2(G311), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n339), .B1(new_n804), .B2(new_n467), .ZN(new_n854));
  INV_X1    g0654(.A(new_n800), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n854), .B1(G294), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n815), .A2(new_n852), .A3(new_n853), .A4(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n855), .A2(G143), .B1(new_n805), .B2(G159), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n433), .B2(new_n787), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(G137), .B2(new_n792), .ZN(new_n860));
  XNOR2_X1  g0660(.A(KEYINPUT104), .B(KEYINPUT34), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT105), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n860), .B(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n248), .B1(new_n795), .B2(new_n202), .ZN(new_n864));
  INV_X1    g0664(.A(new_n790), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n864), .B1(G50), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(G132), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n866), .B1(new_n201), .B2(new_n782), .C1(new_n867), .C2(new_n808), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n857), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n849), .B1(new_n869), .B2(new_n774), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n835), .B2(new_n772), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n846), .A2(new_n871), .ZN(G384));
  NAND2_X1  g0672(.A1(new_n228), .A2(G116), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n510), .A2(new_n508), .ZN(new_n874));
  INV_X1    g0674(.A(new_n509), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n873), .B1(new_n876), .B2(KEYINPUT35), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(KEYINPUT35), .B2(new_n876), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT36), .ZN(new_n879));
  OAI21_X1  g0679(.A(G77), .B1(new_n201), .B2(new_n202), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n229), .A2(new_n880), .B1(G50), .B2(new_n202), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(G1), .A3(new_n755), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT107), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n364), .A2(new_n366), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n687), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT39), .ZN(new_n887));
  INV_X1    g0687(.A(new_n687), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n354), .A2(new_n888), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n363), .B(new_n889), .C1(new_n325), .C2(new_n354), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT37), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n889), .B2(KEYINPUT109), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n890), .B(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n889), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n374), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT38), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n354), .B1(new_n369), .B2(new_n370), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n358), .A2(new_n359), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n361), .A2(new_n269), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n345), .B1(new_n348), .B2(new_n351), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT16), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n904), .A2(new_n272), .A3(new_n352), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n901), .A2(new_n687), .B1(new_n330), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT37), .B1(new_n898), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n371), .A2(new_n372), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT37), .B1(new_n354), .B2(new_n888), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n908), .A2(new_n363), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n687), .B1(new_n905), .B2(new_n330), .ZN(new_n911));
  AOI221_X4 g0711(.A(new_n897), .B1(new_n907), .B2(new_n910), .C1(new_n374), .C2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n887), .B1(new_n896), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n374), .A2(new_n911), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n907), .A2(new_n910), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT38), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n913), .B1(new_n918), .B2(new_n887), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n676), .A2(new_n695), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n886), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n833), .B1(new_n838), .B2(new_n835), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n389), .A2(new_n689), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n416), .B2(KEYINPUT108), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n413), .A2(KEYINPUT108), .A3(new_n415), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n923), .A2(new_n411), .A3(new_n412), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n922), .A2(new_n917), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n921), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n712), .B(new_n446), .C1(new_n719), .C2(new_n711), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n682), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n930), .B(new_n932), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n924), .A2(new_n927), .A3(new_n835), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n746), .A2(new_n934), .A3(KEYINPUT40), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT110), .B1(new_n896), .B2(new_n912), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n374), .A2(new_n894), .ZN(new_n937));
  INV_X1    g0737(.A(new_n892), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n890), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n892), .A2(new_n363), .A3(new_n908), .A4(new_n889), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n897), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT110), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n914), .A2(KEYINPUT38), .A3(new_n915), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n935), .A2(new_n936), .A3(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT40), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n746), .A2(new_n934), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n947), .B1(new_n917), .B2(new_n948), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n446), .A2(new_n746), .ZN(new_n952));
  OAI21_X1  g0752(.A(G330), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n951), .B2(new_n952), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n933), .A2(new_n954), .B1(new_n209), .B2(new_n756), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n933), .A2(new_n954), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n884), .B1(new_n955), .B2(new_n956), .ZN(G367));
  OAI221_X1 g0757(.A(new_n775), .B1(new_n213), .B2(new_n562), .C1(new_n768), .C2(new_n238), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n762), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n584), .A2(new_n689), .ZN(new_n960));
  MUX2_X1   g0760(.A(new_n667), .B(new_n633), .S(new_n960), .Z(new_n961));
  NOR2_X1   g0761(.A1(new_n795), .A2(new_n382), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n787), .A2(new_n812), .B1(new_n790), .B2(new_n201), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n962), .B(new_n963), .C1(G143), .C2(new_n792), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n783), .A2(G68), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n809), .A2(G137), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n248), .B1(new_n804), .B2(new_n379), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(G150), .B2(new_n855), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n964), .A2(new_n965), .A3(new_n966), .A4(new_n968), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n339), .B1(new_n804), .B2(new_n796), .C1(new_n449), .C2(new_n800), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT46), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n865), .A2(G116), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n809), .A2(G317), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n973), .B(new_n974), .C1(new_n971), .C2(new_n972), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n795), .A2(new_n219), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(G294), .B2(new_n786), .ZN(new_n977));
  INV_X1    g0777(.A(G311), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n977), .B1(new_n251), .B2(new_n782), .C1(new_n978), .C2(new_n793), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n969), .B1(new_n975), .B2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT47), .Z(new_n981));
  INV_X1    g0781(.A(new_n774), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n959), .B1(new_n961), .B2(new_n829), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n528), .B(new_n538), .C1(new_n515), .C2(new_n695), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n670), .A2(new_n689), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n700), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT45), .Z(new_n988));
  NOR2_X1   g0788(.A1(new_n700), .A2(new_n986), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT44), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(new_n698), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n699), .A2(new_n694), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n697), .B2(new_n699), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(new_n692), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n752), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n753), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n703), .B(KEYINPUT41), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n758), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n986), .ZN(new_n1001));
  OR3_X1    g0801(.A1(new_n698), .A2(KEYINPUT111), .A3(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(KEYINPUT111), .B1(new_n698), .B2(new_n1001), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(KEYINPUT43), .B2(new_n961), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1002), .A2(new_n1006), .A3(new_n1003), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n699), .A2(new_n694), .A3(new_n986), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1009), .A2(KEYINPUT42), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n538), .B1(new_n984), .B2(new_n624), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n1009), .A2(KEYINPUT42), .B1(new_n695), .B2(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n1010), .A2(new_n1012), .B1(KEYINPUT43), .B2(new_n961), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1008), .B(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n983), .B1(new_n1000), .B2(new_n1015), .ZN(G387));
  NOR2_X1   g0816(.A1(new_n996), .A2(new_n704), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n1018), .A2(KEYINPUT115), .B1(new_n752), .B2(new_n995), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT115), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n995), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n697), .A2(new_n829), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n763), .A2(new_n705), .B1(G107), .B2(new_n213), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n235), .A2(new_n258), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n705), .ZN(new_n1027));
  AOI211_X1 g0827(.A(G45), .B(new_n1027), .C1(G68), .C2(G77), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n277), .A2(G50), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n768), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1025), .B1(new_n1026), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n762), .B1(new_n1033), .B2(new_n776), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT113), .Z(new_n1035));
  OAI22_X1  g0835(.A1(new_n787), .A2(new_n277), .B1(new_n790), .B2(new_n382), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n976), .B(new_n1036), .C1(G159), .C2(new_n792), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n783), .A2(new_n275), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n809), .A2(G150), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n248), .B1(new_n800), .B2(new_n379), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G68), .B2(new_n805), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n248), .B1(new_n823), .B2(G116), .ZN(new_n1043));
  INV_X1    g0843(.A(G294), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n782), .A2(new_n796), .B1(new_n1044), .B2(new_n790), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n855), .A2(G317), .B1(new_n805), .B2(G303), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n787), .B2(new_n978), .C1(new_n801), .C2(new_n793), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT48), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1045), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n1048), .B2(new_n1047), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT49), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1043), .B1(new_n794), .B2(new_n808), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1042), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1054), .A2(KEYINPUT114), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n982), .B1(new_n1054), .B2(KEYINPUT114), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1035), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1023), .A2(new_n758), .B1(new_n1024), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1022), .A2(new_n1058), .ZN(G393));
  AOI21_X1  g0859(.A(new_n704), .B1(new_n992), .B2(new_n996), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n996), .B2(new_n992), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n992), .A2(new_n758), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n767), .A2(new_n246), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1063), .B(new_n775), .C1(new_n219), .C2(new_n213), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT116), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n762), .A2(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n787), .A2(new_n449), .B1(new_n790), .B2(new_n796), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n339), .B1(new_n804), .B2(new_n1044), .C1(new_n251), .C2(new_n795), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(G322), .C2(new_n809), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n855), .A2(G311), .B1(G317), .B2(new_n792), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT52), .Z(new_n1073));
  OAI211_X1 g0873(.A(new_n1071), .B(new_n1073), .C1(new_n467), .C2(new_n782), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT117), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n787), .A2(new_n379), .B1(new_n790), .B2(new_n202), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n248), .B1(new_n804), .B2(new_n277), .C1(new_n816), .C2(new_n795), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(G143), .C2(new_n809), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n793), .A2(new_n433), .B1(new_n800), .B2(new_n812), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT51), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n783), .A2(G77), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1080), .A2(new_n1083), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1076), .A2(new_n1077), .A3(new_n1086), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1066), .B(new_n1068), .C1(new_n1087), .C2(new_n774), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n773), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1088), .B1(new_n1089), .B2(new_n986), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1061), .A2(new_n1062), .A3(new_n1090), .ZN(G390));
  INV_X1    g0891(.A(new_n922), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n928), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n750), .B2(new_n835), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n746), .A2(G330), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n1095), .A2(new_n836), .A3(new_n928), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1092), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n750), .A2(new_n835), .A3(new_n1093), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n928), .B1(new_n1095), .B2(new_n836), .ZN(new_n1099));
  NOR3_X1   g0899(.A1(new_n716), .A2(new_n718), .A3(new_n833), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT118), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n834), .A2(new_n291), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n1100), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n715), .A2(new_n695), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n717), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n715), .A2(KEYINPUT98), .A3(new_n695), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n833), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(KEYINPUT118), .B1(new_n1109), .B2(new_n1102), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1098), .B(new_n1099), .C1(new_n1104), .C2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1097), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1095), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n446), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n931), .A2(new_n682), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1117));
  NOR4_X1   g0917(.A1(new_n747), .A2(new_n749), .A3(new_n836), .A4(new_n928), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n920), .B1(new_n922), .B2(new_n928), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1101), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1109), .A2(KEYINPUT118), .A3(new_n1102), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1120), .A2(new_n1093), .A3(new_n1121), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n936), .A2(new_n945), .A3(new_n920), .ZN(new_n1123));
  AOI221_X4 g0923(.A(new_n1118), .B1(new_n1119), .B2(new_n919), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1096), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1119), .A2(new_n919), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1117), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1115), .B1(new_n1097), .B2(new_n1111), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1126), .A2(new_n1127), .A3(new_n1098), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1122), .A2(new_n1123), .B1(new_n919), .B2(new_n1119), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1130), .B(new_n1131), .C1(new_n1132), .C2(new_n1125), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1129), .A2(new_n1133), .A3(new_n703), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT54), .B(G143), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n248), .B1(new_n804), .B2(new_n1135), .C1(new_n867), .C2(new_n800), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n865), .A2(G150), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT53), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1136), .B(new_n1138), .C1(G125), .C2(new_n809), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n823), .A2(G50), .B1(G137), .B2(new_n786), .ZN(new_n1140));
  INV_X1    g0940(.A(G128), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1140), .B1(new_n1141), .B2(new_n793), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G159), .B2(new_n783), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n339), .B1(new_n804), .B2(new_n219), .C1(new_n467), .C2(new_n800), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n786), .A2(G107), .B1(new_n792), .B2(G283), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1145), .B1(new_n202), .B2(new_n795), .C1(new_n816), .C2(new_n790), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1144), .B(new_n1146), .C1(G294), .C2(new_n809), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1139), .A2(new_n1143), .B1(new_n1084), .B2(new_n1147), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n762), .B1(new_n278), .B2(new_n848), .C1(new_n1148), .C2(new_n982), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n919), .B2(new_n771), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1150), .B1(new_n1151), .B2(new_n758), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1134), .A2(new_n1152), .ZN(G378));
  NOR2_X1   g0953(.A1(new_n248), .A2(G41), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1154), .B1(new_n790), .B2(new_n382), .C1(new_n251), .C2(new_n800), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G283), .B2(new_n809), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n275), .A2(new_n805), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n219), .A2(new_n787), .B1(new_n793), .B2(new_n467), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G58), .B2(new_n823), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1156), .A2(new_n965), .A3(new_n1157), .A4(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT58), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1154), .ZN(new_n1162));
  AOI21_X1  g0962(.A(G50), .B1(new_n332), .B2(new_n257), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1160), .A2(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n805), .A2(G137), .B1(G132), .B2(new_n786), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT119), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n792), .A2(G125), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1141), .B2(new_n800), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1135), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n865), .B2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1166), .B(new_n1170), .C1(new_n433), .C2(new_n782), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(KEYINPUT59), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n332), .B(new_n257), .C1(new_n795), .C2(new_n812), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G124), .B2(new_n809), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1171), .A2(KEYINPUT59), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1164), .B1(new_n1161), .B2(new_n1160), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n774), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n847), .A2(new_n379), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1178), .A2(new_n759), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n438), .A2(new_n888), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT120), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n445), .A2(new_n1183), .ZN(new_n1184));
  XOR2_X1   g0984(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1185));
  NAND4_X1  g0985(.A1(new_n441), .A2(new_n442), .A3(new_n444), .A4(new_n1182), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1185), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1180), .B1(new_n1189), .B2(new_n771), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n946), .A2(G330), .A3(new_n949), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT121), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n946), .A2(KEYINPUT121), .A3(G330), .A4(new_n949), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1189), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n950), .A2(new_n1189), .A3(KEYINPUT121), .A4(G330), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n1196), .A2(new_n930), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n930), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1190), .B1(new_n1200), .B2(new_n758), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1115), .B1(new_n1151), .B2(new_n1130), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n930), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1196), .A2(new_n930), .A3(new_n1197), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(KEYINPUT57), .A3(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n703), .B1(new_n1202), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1133), .A2(new_n1116), .ZN(new_n1209));
  AOI21_X1  g1009(.A(KEYINPUT57), .B1(new_n1209), .B2(new_n1200), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1201), .B1(new_n1208), .B2(new_n1210), .ZN(G375));
  INV_X1    g1011(.A(new_n1112), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1115), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1213), .A2(new_n999), .A3(new_n1117), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n762), .B1(G68), .B2(new_n848), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n793), .A2(new_n1044), .B1(new_n790), .B2(new_n219), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n339), .B1(new_n800), .B2(new_n796), .C1(new_n382), .C2(new_n795), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(G303), .C2(new_n809), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n805), .A2(G107), .B1(G116), .B2(new_n786), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT122), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1218), .A2(new_n1038), .A3(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT123), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n248), .B1(new_n804), .B2(new_n433), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n793), .A2(new_n867), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1225), .A2(KEYINPUT124), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1224), .B(new_n1226), .C1(G137), .C2(new_n855), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n809), .A2(G128), .B1(new_n1225), .B2(KEYINPUT124), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n783), .A2(G50), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n201), .A2(new_n795), .B1(new_n790), .B2(new_n812), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n786), .B2(new_n1169), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .A4(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1223), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1215), .B1(new_n1234), .B2(new_n774), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n1093), .B2(new_n772), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1212), .B2(new_n757), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1214), .A2(new_n1238), .ZN(G381));
  NAND2_X1  g1039(.A1(G378), .A2(KEYINPUT125), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT125), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1134), .A2(new_n1152), .A3(new_n1241), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1243), .B(new_n1201), .C1(new_n1210), .C2(new_n1208), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1058), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n831), .ZN(new_n1247));
  OR4_X1    g1047(.A1(G384), .A2(new_n1247), .A3(G387), .A4(G390), .ZN(new_n1248));
  OR3_X1    g1048(.A1(new_n1244), .A2(new_n1248), .A3(G381), .ZN(G407));
  OAI211_X1 g1049(.A(G407), .B(G213), .C1(G343), .C2(new_n1244), .ZN(G409));
  XNOR2_X1  g1050(.A(G387), .B(KEYINPUT126), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1247), .ZN(new_n1252));
  INV_X1    g1052(.A(G390), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1246), .A2(new_n831), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(G393), .A2(G396), .ZN(new_n1256));
  AOI21_X1  g1056(.A(G390), .B1(new_n1256), .B2(new_n1247), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1251), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT126), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(G387), .B(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1253), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1256), .A2(G390), .A3(new_n1247), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1258), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1209), .A2(new_n999), .A3(new_n1200), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1201), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1240), .A2(new_n1266), .A3(new_n1242), .ZN(new_n1267));
  OAI211_X1 g1067(.A(G378), .B(new_n1201), .C1(new_n1208), .C2(new_n1210), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n688), .A2(G213), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1270), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(G2897), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(G384), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1097), .A2(new_n1111), .A3(new_n1115), .A4(KEYINPUT60), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n703), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1117), .A2(KEYINPUT60), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1277), .B1(new_n1278), .B2(new_n1213), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1275), .B1(new_n1279), .B2(new_n1237), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NOR3_X1   g1081(.A1(new_n1279), .A2(new_n1275), .A3(new_n1237), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1274), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  OR3_X1    g1083(.A1(new_n1279), .A2(new_n1275), .A3(new_n1237), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1284), .A2(new_n1280), .A3(new_n1273), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT61), .B1(new_n1271), .B2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1272), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT63), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1288), .A2(KEYINPUT63), .A3(new_n1289), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1264), .A2(new_n1287), .A3(new_n1292), .A4(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT62), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1288), .A2(new_n1295), .A3(new_n1289), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT61), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1297), .B1(new_n1288), .B2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1295), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1300));
  NOR3_X1   g1100(.A1(new_n1296), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1294), .B1(new_n1301), .B2(new_n1264), .ZN(G405));
  NAND2_X1  g1102(.A1(new_n1243), .A2(G375), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1268), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT127), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1289), .A2(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(KEYINPUT127), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1304), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1303), .A2(new_n1305), .A3(new_n1289), .A4(new_n1268), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n1264), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1308), .A2(new_n1263), .A3(new_n1258), .A4(new_n1309), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(G402));
endmodule


