

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(n631), .A2(n537), .ZN(n634) );
  XOR2_X1 U549 ( .A(KEYINPUT65), .B(n539), .Z(n639) );
  OR2_X1 U550 ( .A1(n781), .A2(n793), .ZN(n513) );
  OR2_X1 U551 ( .A1(n745), .A2(KEYINPUT33), .ZN(n514) );
  OR2_X1 U552 ( .A1(n978), .A2(n687), .ZN(n515) );
  INV_X1 U553 ( .A(n701), .ZN(n720) );
  NAND2_X1 U554 ( .A1(G8), .A2(n720), .ZN(n793) );
  NOR2_X1 U555 ( .A1(n671), .A2(G1384), .ZN(n747) );
  NOR2_X2 U556 ( .A1(G2104), .A2(n521), .ZN(n885) );
  AND2_X1 U557 ( .A1(n782), .A2(n513), .ZN(n783) );
  NOR2_X1 U558 ( .A1(G543), .A2(G651), .ZN(n635) );
  XNOR2_X1 U559 ( .A(KEYINPUT15), .B(n580), .ZN(n978) );
  BUF_X1 U560 ( .A(n671), .Z(G164) );
  INV_X1 U561 ( .A(G2105), .ZN(n521) );
  AND2_X1 U562 ( .A1(n521), .A2(G2104), .ZN(n881) );
  NAND2_X1 U563 ( .A1(G102), .A2(n881), .ZN(n518) );
  NOR2_X1 U564 ( .A1(G2104), .A2(G2105), .ZN(n516) );
  XOR2_X2 U565 ( .A(KEYINPUT17), .B(n516), .Z(n882) );
  NAND2_X1 U566 ( .A1(G138), .A2(n882), .ZN(n517) );
  NAND2_X1 U567 ( .A1(n518), .A2(n517), .ZN(n526) );
  NAND2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  XNOR2_X2 U569 ( .A(n519), .B(KEYINPUT67), .ZN(n886) );
  NAND2_X1 U570 ( .A1(n886), .A2(G114), .ZN(n520) );
  XOR2_X1 U571 ( .A(KEYINPUT83), .B(n520), .Z(n524) );
  NAND2_X1 U572 ( .A1(G126), .A2(n885), .ZN(n522) );
  XNOR2_X1 U573 ( .A(n522), .B(KEYINPUT82), .ZN(n523) );
  NAND2_X1 U574 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U575 ( .A1(n526), .A2(n525), .ZN(n671) );
  NAND2_X1 U576 ( .A1(G125), .A2(n885), .ZN(n527) );
  XNOR2_X1 U577 ( .A(n527), .B(KEYINPUT66), .ZN(n530) );
  NAND2_X1 U578 ( .A1(G101), .A2(n881), .ZN(n528) );
  XOR2_X1 U579 ( .A(KEYINPUT23), .B(n528), .Z(n529) );
  NAND2_X1 U580 ( .A1(n530), .A2(n529), .ZN(n534) );
  NAND2_X1 U581 ( .A1(G137), .A2(n882), .ZN(n532) );
  NAND2_X1 U582 ( .A1(G113), .A2(n886), .ZN(n531) );
  NAND2_X1 U583 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X2 U584 ( .A1(n534), .A2(n533), .ZN(G160) );
  XOR2_X1 U585 ( .A(KEYINPUT0), .B(G543), .Z(n631) );
  INV_X1 U586 ( .A(G651), .ZN(n537) );
  NAND2_X1 U587 ( .A1(G78), .A2(n634), .ZN(n536) );
  NAND2_X1 U588 ( .A1(G91), .A2(n635), .ZN(n535) );
  NAND2_X1 U589 ( .A1(n536), .A2(n535), .ZN(n543) );
  NOR2_X1 U590 ( .A1(G543), .A2(n537), .ZN(n538) );
  XOR2_X1 U591 ( .A(KEYINPUT1), .B(n538), .Z(n638) );
  NAND2_X1 U592 ( .A1(G65), .A2(n638), .ZN(n541) );
  NOR2_X1 U593 ( .A1(n631), .A2(G651), .ZN(n539) );
  NAND2_X1 U594 ( .A1(G53), .A2(n639), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n541), .A2(n540), .ZN(n542) );
  OR2_X1 U596 ( .A1(n543), .A2(n542), .ZN(G299) );
  AND2_X1 U597 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U598 ( .A(G132), .ZN(G219) );
  INV_X1 U599 ( .A(G82), .ZN(G220) );
  INV_X1 U600 ( .A(G57), .ZN(G237) );
  NAND2_X1 U601 ( .A1(G77), .A2(n634), .ZN(n545) );
  NAND2_X1 U602 ( .A1(G90), .A2(n635), .ZN(n544) );
  NAND2_X1 U603 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U604 ( .A(KEYINPUT9), .B(n546), .ZN(n550) );
  NAND2_X1 U605 ( .A1(G64), .A2(n638), .ZN(n548) );
  NAND2_X1 U606 ( .A1(G52), .A2(n639), .ZN(n547) );
  AND2_X1 U607 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U608 ( .A1(n550), .A2(n549), .ZN(G301) );
  NAND2_X1 U609 ( .A1(n635), .A2(G89), .ZN(n551) );
  XNOR2_X1 U610 ( .A(n551), .B(KEYINPUT4), .ZN(n553) );
  NAND2_X1 U611 ( .A1(G76), .A2(n634), .ZN(n552) );
  NAND2_X1 U612 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U613 ( .A(n554), .B(KEYINPUT5), .ZN(n559) );
  NAND2_X1 U614 ( .A1(G63), .A2(n638), .ZN(n556) );
  NAND2_X1 U615 ( .A1(G51), .A2(n639), .ZN(n555) );
  NAND2_X1 U616 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U617 ( .A(KEYINPUT6), .B(n557), .Z(n558) );
  NAND2_X1 U618 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U619 ( .A(n560), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U620 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U621 ( .A1(G7), .A2(G661), .ZN(n561) );
  XOR2_X1 U622 ( .A(n561), .B(KEYINPUT10), .Z(n913) );
  NAND2_X1 U623 ( .A1(n913), .A2(G567), .ZN(n562) );
  XOR2_X1 U624 ( .A(KEYINPUT11), .B(n562), .Z(G234) );
  NAND2_X1 U625 ( .A1(n638), .A2(G56), .ZN(n563) );
  XNOR2_X1 U626 ( .A(n563), .B(KEYINPUT14), .ZN(n565) );
  NAND2_X1 U627 ( .A1(G43), .A2(n639), .ZN(n564) );
  NAND2_X1 U628 ( .A1(n565), .A2(n564), .ZN(n572) );
  NAND2_X1 U629 ( .A1(n635), .A2(G81), .ZN(n566) );
  XNOR2_X1 U630 ( .A(n566), .B(KEYINPUT12), .ZN(n568) );
  NAND2_X1 U631 ( .A1(G68), .A2(n634), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT70), .B(n569), .Z(n570) );
  XNOR2_X1 U634 ( .A(KEYINPUT13), .B(n570), .ZN(n571) );
  NOR2_X1 U635 ( .A1(n572), .A2(n571), .ZN(n965) );
  NAND2_X1 U636 ( .A1(n965), .A2(G860), .ZN(G153) );
  NAND2_X1 U637 ( .A1(G868), .A2(G301), .ZN(n582) );
  NAND2_X1 U638 ( .A1(n639), .A2(G54), .ZN(n579) );
  NAND2_X1 U639 ( .A1(G92), .A2(n635), .ZN(n574) );
  NAND2_X1 U640 ( .A1(G66), .A2(n638), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U642 ( .A1(G79), .A2(n634), .ZN(n575) );
  XNOR2_X1 U643 ( .A(KEYINPUT71), .B(n575), .ZN(n576) );
  NOR2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  OR2_X1 U646 ( .A1(n978), .A2(G868), .ZN(n581) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(G284) );
  XOR2_X1 U648 ( .A(KEYINPUT72), .B(G868), .Z(n583) );
  NOR2_X1 U649 ( .A1(G286), .A2(n583), .ZN(n585) );
  NOR2_X1 U650 ( .A1(G868), .A2(G299), .ZN(n584) );
  NOR2_X1 U651 ( .A1(n585), .A2(n584), .ZN(G297) );
  INV_X1 U652 ( .A(G860), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n586), .A2(G559), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n587), .A2(n978), .ZN(n588) );
  XNOR2_X1 U655 ( .A(n588), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U656 ( .A1(n978), .A2(G868), .ZN(n589) );
  NOR2_X1 U657 ( .A1(G559), .A2(n589), .ZN(n591) );
  INV_X1 U658 ( .A(G868), .ZN(n653) );
  AND2_X1 U659 ( .A1(n653), .A2(n965), .ZN(n590) );
  NOR2_X1 U660 ( .A1(n591), .A2(n590), .ZN(G282) );
  NAND2_X1 U661 ( .A1(G99), .A2(n881), .ZN(n593) );
  NAND2_X1 U662 ( .A1(G135), .A2(n882), .ZN(n592) );
  NAND2_X1 U663 ( .A1(n593), .A2(n592), .ZN(n599) );
  NAND2_X1 U664 ( .A1(G123), .A2(n885), .ZN(n594) );
  XNOR2_X1 U665 ( .A(n594), .B(KEYINPUT18), .ZN(n597) );
  NAND2_X1 U666 ( .A1(G111), .A2(n886), .ZN(n595) );
  XOR2_X1 U667 ( .A(KEYINPUT73), .B(n595), .Z(n596) );
  NAND2_X1 U668 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U669 ( .A1(n599), .A2(n598), .ZN(n928) );
  XNOR2_X1 U670 ( .A(G2096), .B(n928), .ZN(n600) );
  INV_X1 U671 ( .A(G2100), .ZN(n840) );
  NAND2_X1 U672 ( .A1(n600), .A2(n840), .ZN(G156) );
  NAND2_X1 U673 ( .A1(G559), .A2(n978), .ZN(n601) );
  XOR2_X1 U674 ( .A(n965), .B(n601), .Z(n650) );
  XNOR2_X1 U675 ( .A(KEYINPUT74), .B(n650), .ZN(n602) );
  NOR2_X1 U676 ( .A1(G860), .A2(n602), .ZN(n603) );
  XNOR2_X1 U677 ( .A(n603), .B(KEYINPUT77), .ZN(n612) );
  NAND2_X1 U678 ( .A1(G55), .A2(n639), .ZN(n604) );
  XNOR2_X1 U679 ( .A(n604), .B(KEYINPUT76), .ZN(n611) );
  NAND2_X1 U680 ( .A1(G93), .A2(n635), .ZN(n606) );
  NAND2_X1 U681 ( .A1(G67), .A2(n638), .ZN(n605) );
  NAND2_X1 U682 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U683 ( .A1(G80), .A2(n634), .ZN(n607) );
  XNOR2_X1 U684 ( .A(KEYINPUT75), .B(n607), .ZN(n608) );
  NOR2_X1 U685 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n611), .A2(n610), .ZN(n652) );
  XNOR2_X1 U687 ( .A(n612), .B(n652), .ZN(G145) );
  NAND2_X1 U688 ( .A1(n634), .A2(G72), .ZN(n613) );
  XNOR2_X1 U689 ( .A(n613), .B(KEYINPUT68), .ZN(n615) );
  NAND2_X1 U690 ( .A1(G85), .A2(n635), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U692 ( .A(KEYINPUT69), .B(n616), .ZN(n620) );
  NAND2_X1 U693 ( .A1(G60), .A2(n638), .ZN(n618) );
  NAND2_X1 U694 ( .A1(G47), .A2(n639), .ZN(n617) );
  AND2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n620), .A2(n619), .ZN(G290) );
  NAND2_X1 U697 ( .A1(G86), .A2(n635), .ZN(n622) );
  NAND2_X1 U698 ( .A1(G61), .A2(n638), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U700 ( .A1(n634), .A2(G73), .ZN(n623) );
  XOR2_X1 U701 ( .A(KEYINPUT2), .B(n623), .Z(n624) );
  NOR2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n639), .A2(G48), .ZN(n626) );
  NAND2_X1 U704 ( .A1(n627), .A2(n626), .ZN(G305) );
  NAND2_X1 U705 ( .A1(G49), .A2(n639), .ZN(n629) );
  NAND2_X1 U706 ( .A1(G74), .A2(G651), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U708 ( .A1(n638), .A2(n630), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n631), .A2(G87), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(G288) );
  NAND2_X1 U711 ( .A1(G75), .A2(n634), .ZN(n637) );
  NAND2_X1 U712 ( .A1(G88), .A2(n635), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n637), .A2(n636), .ZN(n643) );
  NAND2_X1 U714 ( .A1(G62), .A2(n638), .ZN(n641) );
  NAND2_X1 U715 ( .A1(G50), .A2(n639), .ZN(n640) );
  NAND2_X1 U716 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U717 ( .A1(n643), .A2(n642), .ZN(G166) );
  XOR2_X1 U718 ( .A(G290), .B(G305), .Z(n644) );
  XNOR2_X1 U719 ( .A(n652), .B(n644), .ZN(n645) );
  XNOR2_X1 U720 ( .A(KEYINPUT19), .B(n645), .ZN(n647) );
  XNOR2_X1 U721 ( .A(G288), .B(KEYINPUT78), .ZN(n646) );
  XNOR2_X1 U722 ( .A(n647), .B(n646), .ZN(n648) );
  XOR2_X1 U723 ( .A(n648), .B(G166), .Z(n649) );
  XNOR2_X1 U724 ( .A(n649), .B(G299), .ZN(n900) );
  XNOR2_X1 U725 ( .A(n650), .B(n900), .ZN(n651) );
  NAND2_X1 U726 ( .A1(n651), .A2(G868), .ZN(n655) );
  NAND2_X1 U727 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U728 ( .A1(n655), .A2(n654), .ZN(G295) );
  NAND2_X1 U729 ( .A1(G2078), .A2(G2084), .ZN(n656) );
  XOR2_X1 U730 ( .A(KEYINPUT20), .B(n656), .Z(n657) );
  NAND2_X1 U731 ( .A1(G2090), .A2(n657), .ZN(n658) );
  XNOR2_X1 U732 ( .A(KEYINPUT21), .B(n658), .ZN(n659) );
  NAND2_X1 U733 ( .A1(n659), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U734 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U735 ( .A1(G120), .A2(G69), .ZN(n660) );
  NOR2_X1 U736 ( .A1(G237), .A2(n660), .ZN(n661) );
  XNOR2_X1 U737 ( .A(KEYINPUT80), .B(n661), .ZN(n662) );
  NAND2_X1 U738 ( .A1(n662), .A2(G108), .ZN(n833) );
  NAND2_X1 U739 ( .A1(G567), .A2(n833), .ZN(n668) );
  NOR2_X1 U740 ( .A1(G220), .A2(G219), .ZN(n663) );
  XNOR2_X1 U741 ( .A(KEYINPUT22), .B(n663), .ZN(n664) );
  NAND2_X1 U742 ( .A1(n664), .A2(G96), .ZN(n665) );
  NOR2_X1 U743 ( .A1(n665), .A2(G218), .ZN(n666) );
  XNOR2_X1 U744 ( .A(n666), .B(KEYINPUT79), .ZN(n834) );
  NAND2_X1 U745 ( .A1(G2106), .A2(n834), .ZN(n667) );
  NAND2_X1 U746 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U747 ( .A(KEYINPUT81), .B(n669), .Z(n856) );
  NAND2_X1 U748 ( .A1(G661), .A2(G483), .ZN(n670) );
  NOR2_X1 U749 ( .A1(n856), .A2(n670), .ZN(n831) );
  NAND2_X1 U750 ( .A1(n831), .A2(G36), .ZN(G176) );
  INV_X1 U751 ( .A(G166), .ZN(G303) );
  INV_X1 U752 ( .A(n747), .ZN(n672) );
  NAND2_X1 U753 ( .A1(G160), .A2(G40), .ZN(n746) );
  NOR2_X4 U754 ( .A1(n672), .A2(n746), .ZN(n701) );
  NOR2_X1 U755 ( .A1(G1966), .A2(n793), .ZN(n735) );
  NOR2_X1 U756 ( .A1(G2084), .A2(n720), .ZN(n731) );
  NOR2_X1 U757 ( .A1(n735), .A2(n731), .ZN(n673) );
  XNOR2_X1 U758 ( .A(n673), .B(KEYINPUT96), .ZN(n674) );
  NAND2_X1 U759 ( .A1(n674), .A2(G8), .ZN(n675) );
  XNOR2_X1 U760 ( .A(KEYINPUT30), .B(n675), .ZN(n676) );
  NOR2_X1 U761 ( .A1(G168), .A2(n676), .ZN(n677) );
  XNOR2_X1 U762 ( .A(n677), .B(KEYINPUT97), .ZN(n681) );
  XOR2_X1 U763 ( .A(KEYINPUT25), .B(G2078), .Z(n942) );
  NOR2_X1 U764 ( .A1(n942), .A2(n720), .ZN(n679) );
  NOR2_X1 U765 ( .A1(n701), .A2(G1961), .ZN(n678) );
  NOR2_X1 U766 ( .A1(n679), .A2(n678), .ZN(n713) );
  NAND2_X1 U767 ( .A1(n713), .A2(G301), .ZN(n680) );
  NAND2_X1 U768 ( .A1(n681), .A2(n680), .ZN(n683) );
  XOR2_X1 U769 ( .A(KEYINPUT98), .B(KEYINPUT31), .Z(n682) );
  XNOR2_X1 U770 ( .A(n683), .B(n682), .ZN(n717) );
  NAND2_X1 U771 ( .A1(G1348), .A2(n720), .ZN(n685) );
  NAND2_X1 U772 ( .A1(G2067), .A2(n701), .ZN(n684) );
  NAND2_X1 U773 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U774 ( .A(KEYINPUT93), .B(n686), .ZN(n687) );
  AND2_X1 U775 ( .A1(n978), .A2(n687), .ZN(n699) );
  XNOR2_X1 U776 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n689) );
  NOR2_X1 U777 ( .A1(G1996), .A2(n689), .ZN(n697) );
  INV_X1 U778 ( .A(G1341), .ZN(n966) );
  NAND2_X1 U779 ( .A1(n966), .A2(n689), .ZN(n688) );
  NAND2_X1 U780 ( .A1(n688), .A2(n720), .ZN(n692) );
  AND2_X1 U781 ( .A1(G1996), .A2(n701), .ZN(n690) );
  NAND2_X1 U782 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U783 ( .A1(n692), .A2(n691), .ZN(n694) );
  INV_X1 U784 ( .A(n965), .ZN(n693) );
  NOR2_X1 U785 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U786 ( .A1(n515), .A2(n695), .ZN(n696) );
  NOR2_X1 U787 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U788 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U789 ( .A(n700), .B(KEYINPUT94), .ZN(n707) );
  NAND2_X1 U790 ( .A1(n701), .A2(G2072), .ZN(n702) );
  XOR2_X1 U791 ( .A(KEYINPUT27), .B(n702), .Z(n704) );
  NAND2_X1 U792 ( .A1(G1956), .A2(n720), .ZN(n703) );
  NAND2_X1 U793 ( .A1(n704), .A2(n703), .ZN(n708) );
  NOR2_X1 U794 ( .A1(G299), .A2(n708), .ZN(n705) );
  XNOR2_X1 U795 ( .A(KEYINPUT95), .B(n705), .ZN(n706) );
  NAND2_X1 U796 ( .A1(n707), .A2(n706), .ZN(n711) );
  NAND2_X1 U797 ( .A1(G299), .A2(n708), .ZN(n709) );
  XNOR2_X1 U798 ( .A(n709), .B(KEYINPUT28), .ZN(n710) );
  NAND2_X1 U799 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U800 ( .A(n712), .B(KEYINPUT29), .ZN(n715) );
  NOR2_X1 U801 ( .A1(G301), .A2(n713), .ZN(n714) );
  NOR2_X1 U802 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U803 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U804 ( .A(n718), .B(KEYINPUT99), .ZN(n732) );
  AND2_X1 U805 ( .A1(G286), .A2(G8), .ZN(n719) );
  AND2_X1 U806 ( .A1(n732), .A2(n719), .ZN(n728) );
  INV_X1 U807 ( .A(G8), .ZN(n726) );
  NOR2_X1 U808 ( .A1(G1971), .A2(n793), .ZN(n722) );
  NOR2_X1 U809 ( .A1(G2090), .A2(n720), .ZN(n721) );
  NOR2_X1 U810 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U811 ( .A1(n723), .A2(G303), .ZN(n724) );
  XOR2_X1 U812 ( .A(KEYINPUT101), .B(n724), .Z(n725) );
  NOR2_X1 U813 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U814 ( .A1(n728), .A2(n727), .ZN(n730) );
  XNOR2_X1 U815 ( .A(KEYINPUT32), .B(KEYINPUT102), .ZN(n729) );
  XNOR2_X1 U816 ( .A(n730), .B(n729), .ZN(n739) );
  NAND2_X1 U817 ( .A1(n731), .A2(G8), .ZN(n737) );
  INV_X1 U818 ( .A(KEYINPUT100), .ZN(n733) );
  XNOR2_X1 U819 ( .A(n733), .B(n732), .ZN(n734) );
  NOR2_X1 U820 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U821 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U822 ( .A1(n739), .A2(n738), .ZN(n787) );
  NOR2_X1 U823 ( .A1(G1976), .A2(G288), .ZN(n780) );
  NOR2_X1 U824 ( .A1(G1971), .A2(G303), .ZN(n740) );
  NOR2_X1 U825 ( .A1(n780), .A2(n740), .ZN(n972) );
  NAND2_X1 U826 ( .A1(n787), .A2(n972), .ZN(n741) );
  XNOR2_X1 U827 ( .A(n741), .B(KEYINPUT103), .ZN(n744) );
  NAND2_X1 U828 ( .A1(G1976), .A2(G288), .ZN(n964) );
  INV_X1 U829 ( .A(n964), .ZN(n742) );
  OR2_X1 U830 ( .A1(n793), .A2(n742), .ZN(n743) );
  NOR2_X1 U831 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U832 ( .A(G1981), .B(G305), .Z(n974) );
  NOR2_X1 U833 ( .A1(n747), .A2(n746), .ZN(n812) );
  XNOR2_X1 U834 ( .A(G2067), .B(KEYINPUT37), .ZN(n810) );
  NAND2_X1 U835 ( .A1(G104), .A2(n881), .ZN(n749) );
  NAND2_X1 U836 ( .A1(G140), .A2(n882), .ZN(n748) );
  NAND2_X1 U837 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U838 ( .A(KEYINPUT34), .B(n750), .ZN(n756) );
  NAND2_X1 U839 ( .A1(n885), .A2(G128), .ZN(n751) );
  XNOR2_X1 U840 ( .A(n751), .B(KEYINPUT84), .ZN(n753) );
  NAND2_X1 U841 ( .A1(G116), .A2(n886), .ZN(n752) );
  NAND2_X1 U842 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U843 ( .A(KEYINPUT35), .B(n754), .Z(n755) );
  NOR2_X1 U844 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U845 ( .A(KEYINPUT36), .B(n757), .ZN(n897) );
  NOR2_X1 U846 ( .A1(n810), .A2(n897), .ZN(n927) );
  NAND2_X1 U847 ( .A1(n812), .A2(n927), .ZN(n758) );
  XNOR2_X1 U848 ( .A(KEYINPUT85), .B(n758), .ZN(n807) );
  NAND2_X1 U849 ( .A1(G119), .A2(n885), .ZN(n760) );
  NAND2_X1 U850 ( .A1(G95), .A2(n881), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n763) );
  NAND2_X1 U852 ( .A1(n886), .A2(G107), .ZN(n761) );
  XOR2_X1 U853 ( .A(KEYINPUT86), .B(n761), .Z(n762) );
  NOR2_X1 U854 ( .A1(n763), .A2(n762), .ZN(n765) );
  NAND2_X1 U855 ( .A1(n882), .A2(G131), .ZN(n764) );
  AND2_X1 U856 ( .A1(n765), .A2(n764), .ZN(n873) );
  XNOR2_X1 U857 ( .A(KEYINPUT87), .B(G1991), .ZN(n946) );
  NOR2_X1 U858 ( .A1(n873), .A2(n946), .ZN(n775) );
  XOR2_X1 U859 ( .A(KEYINPUT38), .B(KEYINPUT88), .Z(n767) );
  NAND2_X1 U860 ( .A1(G105), .A2(n881), .ZN(n766) );
  XNOR2_X1 U861 ( .A(n767), .B(n766), .ZN(n771) );
  NAND2_X1 U862 ( .A1(G129), .A2(n885), .ZN(n769) );
  NAND2_X1 U863 ( .A1(G141), .A2(n882), .ZN(n768) );
  NAND2_X1 U864 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U865 ( .A1(n771), .A2(n770), .ZN(n773) );
  NAND2_X1 U866 ( .A1(n886), .A2(G117), .ZN(n772) );
  NAND2_X1 U867 ( .A1(n773), .A2(n772), .ZN(n876) );
  AND2_X1 U868 ( .A1(n876), .A2(G1996), .ZN(n774) );
  NOR2_X1 U869 ( .A1(n775), .A2(n774), .ZN(n925) );
  XNOR2_X1 U870 ( .A(KEYINPUT89), .B(n812), .ZN(n776) );
  NOR2_X1 U871 ( .A1(n925), .A2(n776), .ZN(n804) );
  XNOR2_X1 U872 ( .A(KEYINPUT90), .B(n804), .ZN(n777) );
  NOR2_X1 U873 ( .A1(n807), .A2(n777), .ZN(n778) );
  XOR2_X1 U874 ( .A(n778), .B(KEYINPUT91), .Z(n796) );
  AND2_X1 U875 ( .A1(n974), .A2(n796), .ZN(n779) );
  XNOR2_X1 U876 ( .A(G1986), .B(G290), .ZN(n983) );
  NAND2_X1 U877 ( .A1(n983), .A2(n812), .ZN(n784) );
  AND2_X1 U878 ( .A1(n779), .A2(n784), .ZN(n782) );
  NAND2_X1 U879 ( .A1(n780), .A2(KEYINPUT33), .ZN(n781) );
  NAND2_X1 U880 ( .A1(n514), .A2(n783), .ZN(n817) );
  INV_X1 U881 ( .A(n784), .ZN(n800) );
  NOR2_X1 U882 ( .A1(G2090), .A2(G303), .ZN(n785) );
  XNOR2_X1 U883 ( .A(n785), .B(KEYINPUT104), .ZN(n786) );
  NAND2_X1 U884 ( .A1(n786), .A2(G8), .ZN(n788) );
  NAND2_X1 U885 ( .A1(n788), .A2(n787), .ZN(n790) );
  AND2_X1 U886 ( .A1(n793), .A2(n796), .ZN(n789) );
  AND2_X1 U887 ( .A1(n790), .A2(n789), .ZN(n798) );
  NOR2_X1 U888 ( .A1(G1981), .A2(G305), .ZN(n791) );
  XOR2_X1 U889 ( .A(n791), .B(KEYINPUT24), .Z(n792) );
  NOR2_X1 U890 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U891 ( .A(n794), .B(KEYINPUT92), .ZN(n795) );
  AND2_X1 U892 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U893 ( .A1(n798), .A2(n797), .ZN(n799) );
  OR2_X1 U894 ( .A1(n800), .A2(n799), .ZN(n815) );
  NOR2_X1 U895 ( .A1(G1996), .A2(n876), .ZN(n801) );
  XOR2_X1 U896 ( .A(KEYINPUT105), .B(n801), .Z(n919) );
  NOR2_X1 U897 ( .A1(G1986), .A2(G290), .ZN(n802) );
  AND2_X1 U898 ( .A1(n946), .A2(n873), .ZN(n929) );
  NOR2_X1 U899 ( .A1(n802), .A2(n929), .ZN(n803) );
  NOR2_X1 U900 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U901 ( .A1(n919), .A2(n805), .ZN(n806) );
  XNOR2_X1 U902 ( .A(KEYINPUT39), .B(n806), .ZN(n809) );
  INV_X1 U903 ( .A(n807), .ZN(n808) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n810), .A2(n897), .ZN(n933) );
  NAND2_X1 U906 ( .A1(n811), .A2(n933), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n814) );
  AND2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U909 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U910 ( .A(KEYINPUT40), .B(n818), .ZN(G329) );
  XNOR2_X1 U911 ( .A(G2454), .B(G2451), .ZN(n827) );
  XNOR2_X1 U912 ( .A(G2430), .B(G2446), .ZN(n825) );
  XOR2_X1 U913 ( .A(G2435), .B(G2427), .Z(n820) );
  XNOR2_X1 U914 ( .A(KEYINPUT106), .B(G2438), .ZN(n819) );
  XNOR2_X1 U915 ( .A(n820), .B(n819), .ZN(n821) );
  XOR2_X1 U916 ( .A(n821), .B(G2443), .Z(n823) );
  XOR2_X1 U917 ( .A(G1348), .B(n966), .Z(n822) );
  XNOR2_X1 U918 ( .A(n823), .B(n822), .ZN(n824) );
  XNOR2_X1 U919 ( .A(n825), .B(n824), .ZN(n826) );
  XNOR2_X1 U920 ( .A(n827), .B(n826), .ZN(n828) );
  NAND2_X1 U921 ( .A1(n828), .A2(G14), .ZN(n907) );
  XNOR2_X1 U922 ( .A(KEYINPUT107), .B(n907), .ZN(G401) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n913), .ZN(G217) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U925 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n830) );
  XNOR2_X1 U927 ( .A(KEYINPUT108), .B(n830), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n832), .A2(n831), .ZN(G188) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G108), .ZN(G238) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  INV_X1 U933 ( .A(G69), .ZN(G235) );
  NOR2_X1 U934 ( .A1(n834), .A2(n833), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  XOR2_X1 U936 ( .A(KEYINPUT42), .B(G2090), .Z(n836) );
  XNOR2_X1 U937 ( .A(G2078), .B(G2084), .ZN(n835) );
  XNOR2_X1 U938 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U939 ( .A(n837), .B(G2096), .Z(n839) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2072), .ZN(n838) );
  XNOR2_X1 U941 ( .A(n839), .B(n838), .ZN(n844) );
  XOR2_X1 U942 ( .A(KEYINPUT43), .B(G2678), .Z(n842) );
  XOR2_X1 U943 ( .A(KEYINPUT109), .B(n840), .Z(n841) );
  XNOR2_X1 U944 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U945 ( .A(n844), .B(n843), .Z(G227) );
  XOR2_X1 U946 ( .A(KEYINPUT111), .B(G1986), .Z(n846) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1991), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U949 ( .A(n847), .B(KEYINPUT41), .Z(n849) );
  XNOR2_X1 U950 ( .A(G1961), .B(G1966), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U952 ( .A(G1956), .B(G1971), .Z(n851) );
  XNOR2_X1 U953 ( .A(G1981), .B(G1976), .ZN(n850) );
  XNOR2_X1 U954 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U955 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U956 ( .A(KEYINPUT110), .B(G2474), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(G229) );
  INV_X1 U958 ( .A(n856), .ZN(G319) );
  NAND2_X1 U959 ( .A1(n885), .A2(G124), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n857), .B(KEYINPUT44), .ZN(n859) );
  NAND2_X1 U961 ( .A1(G100), .A2(n881), .ZN(n858) );
  NAND2_X1 U962 ( .A1(n859), .A2(n858), .ZN(n863) );
  NAND2_X1 U963 ( .A1(G136), .A2(n882), .ZN(n861) );
  NAND2_X1 U964 ( .A1(G112), .A2(n886), .ZN(n860) );
  NAND2_X1 U965 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U966 ( .A1(n863), .A2(n862), .ZN(G162) );
  NAND2_X1 U967 ( .A1(G130), .A2(n885), .ZN(n865) );
  NAND2_X1 U968 ( .A1(G118), .A2(n886), .ZN(n864) );
  NAND2_X1 U969 ( .A1(n865), .A2(n864), .ZN(n871) );
  NAND2_X1 U970 ( .A1(G106), .A2(n881), .ZN(n867) );
  NAND2_X1 U971 ( .A1(G142), .A2(n882), .ZN(n866) );
  NAND2_X1 U972 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U973 ( .A(KEYINPUT45), .B(n868), .Z(n869) );
  XNOR2_X1 U974 ( .A(KEYINPUT112), .B(n869), .ZN(n870) );
  NOR2_X1 U975 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U976 ( .A(n872), .B(n928), .Z(n875) );
  XNOR2_X1 U977 ( .A(G164), .B(n873), .ZN(n874) );
  XNOR2_X1 U978 ( .A(n875), .B(n874), .ZN(n880) );
  XOR2_X1 U979 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n878) );
  XOR2_X1 U980 ( .A(n876), .B(G162), .Z(n877) );
  XNOR2_X1 U981 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U982 ( .A(n880), .B(n879), .Z(n895) );
  NAND2_X1 U983 ( .A1(G103), .A2(n881), .ZN(n884) );
  NAND2_X1 U984 ( .A1(G139), .A2(n882), .ZN(n883) );
  NAND2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n893) );
  XNOR2_X1 U986 ( .A(KEYINPUT114), .B(KEYINPUT47), .ZN(n891) );
  NAND2_X1 U987 ( .A1(n885), .A2(G127), .ZN(n889) );
  NAND2_X1 U988 ( .A1(n886), .A2(G115), .ZN(n887) );
  XOR2_X1 U989 ( .A(KEYINPUT113), .B(n887), .Z(n888) );
  NAND2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U991 ( .A(n891), .B(n890), .Z(n892) );
  NOR2_X1 U992 ( .A1(n893), .A2(n892), .ZN(n914) );
  XNOR2_X1 U993 ( .A(G160), .B(n914), .ZN(n894) );
  XNOR2_X1 U994 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U995 ( .A(n897), .B(n896), .Z(n898) );
  NOR2_X1 U996 ( .A1(G37), .A2(n898), .ZN(n899) );
  XOR2_X1 U997 ( .A(KEYINPUT115), .B(n899), .Z(G395) );
  XOR2_X1 U998 ( .A(n900), .B(n965), .Z(n902) );
  XOR2_X1 U999 ( .A(G301), .B(n978), .Z(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1001 ( .A(G286), .B(n903), .Z(n904) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n904), .ZN(G397) );
  XNOR2_X1 U1003 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n906) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n905) );
  XNOR2_X1 U1005 ( .A(n906), .B(n905), .ZN(n909) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n907), .ZN(n908) );
  NOR2_X1 U1007 ( .A1(n909), .A2(n908), .ZN(n910) );
  XOR2_X1 U1008 ( .A(KEYINPUT117), .B(n910), .Z(n912) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1010 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(n913), .ZN(G223) );
  INV_X1 U1013 ( .A(G301), .ZN(G171) );
  INV_X1 U1014 ( .A(KEYINPUT55), .ZN(n961) );
  XOR2_X1 U1015 ( .A(G2072), .B(n914), .Z(n916) );
  XOR2_X1 U1016 ( .A(G164), .B(G2078), .Z(n915) );
  NOR2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1018 ( .A(KEYINPUT50), .B(n917), .ZN(n922) );
  XOR2_X1 U1019 ( .A(G2090), .B(G162), .Z(n918) );
  NOR2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1021 ( .A(KEYINPUT51), .B(n920), .Z(n921) );
  NAND2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n936) );
  XNOR2_X1 U1023 ( .A(G160), .B(G2084), .ZN(n923) );
  XNOR2_X1 U1024 ( .A(n923), .B(KEYINPUT118), .ZN(n924) );
  NAND2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n931) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(KEYINPUT119), .B(n932), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(KEYINPUT52), .B(n937), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n961), .A2(n938), .ZN(n939) );
  NAND2_X1 U1034 ( .A1(n939), .A2(G29), .ZN(n1019) );
  XNOR2_X1 U1035 ( .A(G2067), .B(G26), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(G2072), .B(G33), .ZN(n940) );
  NOR2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n953) );
  XOR2_X1 U1038 ( .A(n942), .B(G27), .Z(n945) );
  XOR2_X1 U1039 ( .A(G32), .B(KEYINPUT122), .Z(n943) );
  XNOR2_X1 U1040 ( .A(G1996), .B(n943), .ZN(n944) );
  NAND2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n951) );
  XNOR2_X1 U1042 ( .A(KEYINPUT120), .B(G25), .ZN(n947) );
  XNOR2_X1 U1043 ( .A(n947), .B(n946), .ZN(n948) );
  NAND2_X1 U1044 ( .A1(n948), .A2(G28), .ZN(n949) );
  XOR2_X1 U1045 ( .A(KEYINPUT121), .B(n949), .Z(n950) );
  NOR2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(n954), .B(KEYINPUT53), .ZN(n957) );
  XOR2_X1 U1049 ( .A(G2084), .B(G34), .Z(n955) );
  XNOR2_X1 U1050 ( .A(KEYINPUT54), .B(n955), .ZN(n956) );
  NAND2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(G35), .B(G2090), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(n961), .B(n960), .ZN(n962) );
  NOR2_X1 U1055 ( .A1(G29), .A2(n962), .ZN(n1015) );
  INV_X1 U1056 ( .A(G16), .ZN(n1011) );
  XOR2_X1 U1057 ( .A(n1011), .B(KEYINPUT56), .Z(n987) );
  NAND2_X1 U1058 ( .A1(G1971), .A2(G303), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n970) );
  XOR2_X1 U1060 ( .A(G299), .B(G1956), .Z(n968) );
  XOR2_X1 U1061 ( .A(n966), .B(n965), .Z(n967) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n977) );
  XNOR2_X1 U1065 ( .A(G168), .B(G1966), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1067 ( .A(KEYINPUT57), .B(n975), .Z(n976) );
  NOR2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n985) );
  XOR2_X1 U1069 ( .A(G171), .B(G1961), .Z(n980) );
  XOR2_X1 U1070 ( .A(n978), .B(G1348), .Z(n979) );
  NOR2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(n981), .B(KEYINPUT123), .ZN(n982) );
  NOR2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1074 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1075 ( .A1(n987), .A2(n986), .ZN(n1013) );
  XOR2_X1 U1076 ( .A(G1986), .B(G24), .Z(n990) );
  XNOR2_X1 U1077 ( .A(G22), .B(KEYINPUT125), .ZN(n988) );
  XNOR2_X1 U1078 ( .A(n988), .B(G1971), .ZN(n989) );
  NAND2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n992) );
  XNOR2_X1 U1080 ( .A(G23), .B(G1976), .ZN(n991) );
  NOR2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1082 ( .A(KEYINPUT58), .B(n993), .Z(n1008) );
  XOR2_X1 U1083 ( .A(G1961), .B(G5), .Z(n1003) );
  XOR2_X1 U1084 ( .A(G19), .B(G1341), .Z(n997) );
  XNOR2_X1 U1085 ( .A(G1981), .B(G6), .ZN(n995) );
  XNOR2_X1 U1086 ( .A(G20), .B(G1956), .ZN(n994) );
  NOR2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n1000) );
  XOR2_X1 U1089 ( .A(KEYINPUT59), .B(G1348), .Z(n998) );
  XNOR2_X1 U1090 ( .A(G4), .B(n998), .ZN(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(KEYINPUT60), .B(n1001), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(G21), .B(G1966), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1096 ( .A(KEYINPUT124), .B(n1006), .Z(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(KEYINPUT61), .B(n1009), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1102 ( .A1(G11), .A2(n1016), .ZN(n1017) );
  XOR2_X1 U1103 ( .A(KEYINPUT126), .B(n1017), .Z(n1018) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1020), .ZN(G150) );
  INV_X1 U1106 ( .A(G150), .ZN(G311) );
endmodule

