//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  OR2_X1    g000(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G137), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G134), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n187), .A2(new_n189), .A3(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(KEYINPUT65), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G137), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT11), .A2(G134), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n188), .A2(G134), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n191), .A2(new_n196), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G131), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n191), .A2(new_n196), .A3(new_n201), .A4(new_n198), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT75), .ZN(new_n204));
  INV_X1    g018(.A(G107), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G104), .ZN(new_n206));
  INV_X1    g020(.A(G104), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT3), .B1(new_n207), .B2(G107), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n205), .A3(G104), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(KEYINPUT75), .A3(G107), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n206), .A2(new_n208), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT76), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(G101), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT4), .B1(new_n212), .B2(G101), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n213), .B1(new_n212), .B2(G101), .ZN(new_n217));
  NOR3_X1   g031(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G143), .ZN(new_n220));
  INV_X1    g034(.A(G143), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G146), .ZN(new_n222));
  OR2_X1    g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  NAND2_X1  g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n220), .A2(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n220), .A2(new_n222), .A3(new_n224), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT4), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n212), .A2(new_n229), .A3(G101), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G101), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n205), .A2(G104), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n207), .A2(G107), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AND4_X1   g049(.A1(new_n206), .A2(new_n208), .A3(new_n210), .A4(new_n211), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(new_n232), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n220), .A2(new_n222), .A3(new_n239), .A4(G128), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n221), .A2(KEYINPUT1), .A3(G146), .ZN(new_n241));
  XNOR2_X1  g055(.A(G143), .B(G146), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n240), .B(new_n241), .C1(G128), .C2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT10), .ZN(new_n244));
  OAI22_X1  g058(.A1(new_n218), .A2(new_n231), .B1(new_n238), .B2(new_n244), .ZN(new_n245));
  XOR2_X1   g059(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n246));
  INV_X1    g060(.A(KEYINPUT77), .ZN(new_n247));
  AOI21_X1  g061(.A(G128), .B1(new_n220), .B2(new_n222), .ZN(new_n248));
  INV_X1    g062(.A(new_n241), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OAI211_X1 g064(.A(KEYINPUT77), .B(new_n241), .C1(new_n242), .C2(G128), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n240), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT78), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n252), .A2(new_n253), .A3(new_n237), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n253), .B1(new_n252), .B2(new_n237), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n246), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT80), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  OAI211_X1 g072(.A(KEYINPUT80), .B(new_n246), .C1(new_n254), .C2(new_n255), .ZN(new_n259));
  AOI211_X1 g073(.A(new_n203), .B(new_n245), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(G110), .B(G140), .ZN(new_n261));
  INV_X1    g075(.A(G953), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n262), .A2(G227), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n261), .B(new_n263), .Z(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  OAI22_X1  g080(.A1(new_n254), .A2(new_n255), .B1(new_n243), .B2(new_n237), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT12), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n203), .A2(KEYINPUT81), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n268), .B1(new_n267), .B2(new_n269), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n266), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n245), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n252), .A2(new_n237), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT78), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n252), .A2(new_n237), .A3(new_n253), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT80), .B1(new_n279), .B2(new_n246), .ZN(new_n280));
  INV_X1    g094(.A(new_n259), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n275), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT83), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n283), .A3(new_n203), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n245), .B1(new_n258), .B2(new_n259), .ZN(new_n285));
  INV_X1    g099(.A(new_n203), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT83), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n260), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n274), .B1(new_n288), .B2(new_n264), .ZN(new_n289));
  INV_X1    g103(.A(G469), .ZN(new_n290));
  INV_X1    g104(.A(G902), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT82), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n267), .A2(new_n269), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT12), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n270), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n293), .B1(new_n260), .B2(new_n296), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n286), .B(new_n275), .C1(new_n280), .C2(new_n281), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n273), .A2(new_n298), .A3(KEYINPUT82), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(new_n265), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n283), .B1(new_n282), .B2(new_n203), .ZN(new_n301));
  NOR3_X1   g115(.A1(new_n285), .A2(KEYINPUT83), .A3(new_n286), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n266), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n291), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT84), .B1(new_n305), .B2(G469), .ZN(new_n306));
  AOI21_X1  g120(.A(G902), .B1(new_n300), .B2(new_n303), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT84), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n307), .A2(new_n308), .A3(new_n290), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n292), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT23), .ZN(new_n311));
  INV_X1    g125(.A(G119), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n311), .B1(new_n312), .B2(G128), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(G128), .ZN(new_n314));
  INV_X1    g128(.A(G128), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(KEYINPUT23), .A3(G119), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n313), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  XOR2_X1   g131(.A(KEYINPUT24), .B(G110), .Z(new_n318));
  XNOR2_X1  g132(.A(G119), .B(G128), .ZN(new_n319));
  AOI22_X1  g133(.A1(G110), .A2(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G125), .ZN(new_n322));
  INV_X1    g136(.A(G125), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G140), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n324), .A3(KEYINPUT16), .ZN(new_n325));
  OR3_X1    g139(.A1(new_n323), .A2(KEYINPUT16), .A3(G140), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n326), .A3(G146), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(G146), .B1(new_n325), .B2(new_n326), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n320), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI22_X1  g144(.A1(new_n317), .A2(G110), .B1(new_n318), .B2(new_n319), .ZN(new_n331));
  XNOR2_X1  g145(.A(G125), .B(G140), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n219), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n327), .A3(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT22), .B(G137), .ZN(new_n335));
  INV_X1    g149(.A(G221), .ZN(new_n336));
  INV_X1    g150(.A(G234), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n336), .A2(new_n337), .A3(G953), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n335), .B(new_n338), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n330), .A2(new_n334), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n339), .B1(new_n330), .B2(new_n334), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n291), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT74), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT25), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  OAI221_X1 g160(.A(new_n291), .B1(new_n343), .B2(new_n344), .C1(new_n340), .C2(new_n341), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n346), .A2(new_n347), .B1(new_n343), .B2(new_n344), .ZN(new_n348));
  INV_X1    g162(.A(G217), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n349), .B1(G234), .B2(new_n291), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n340), .A2(new_n341), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n350), .A2(G902), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n352), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT71), .ZN(new_n358));
  INV_X1    g172(.A(G113), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT2), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT2), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G113), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(G116), .B(G119), .ZN(new_n364));
  NOR3_X1   g178(.A1(new_n363), .A2(new_n364), .A3(KEYINPUT69), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT69), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n312), .A2(G116), .ZN(new_n367));
  INV_X1    g181(.A(G116), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G119), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT2), .B(G113), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n366), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n370), .A2(new_n371), .ZN(new_n373));
  OAI22_X1  g187(.A1(new_n365), .A2(new_n372), .B1(KEYINPUT68), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT69), .B1(new_n363), .B2(new_n364), .ZN(new_n375));
  AOI21_X1  g189(.A(KEYINPUT68), .B1(new_n363), .B2(new_n364), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n370), .A2(new_n371), .A3(new_n366), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n243), .A2(new_n202), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n189), .A2(KEYINPUT67), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT65), .B(G137), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n381), .B1(new_n382), .B2(G134), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n192), .A2(new_n194), .ZN(new_n384));
  INV_X1    g198(.A(G134), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(KEYINPUT67), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n201), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n380), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n227), .B1(new_n200), .B2(new_n202), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n379), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT26), .B(G101), .ZN(new_n391));
  NOR2_X1   g205(.A1(G237), .A2(G953), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G210), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n391), .B(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n394), .B(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n358), .B1(new_n390), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n379), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n197), .B1(new_n382), .B2(new_n195), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n201), .B1(new_n400), .B2(new_n191), .ZN(new_n401));
  AND4_X1   g215(.A1(new_n201), .A2(new_n191), .A3(new_n196), .A4(new_n198), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n228), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n384), .A2(new_n385), .B1(KEYINPUT67), .B2(new_n189), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT67), .ZN(new_n405));
  AOI211_X1 g219(.A(new_n405), .B(G134), .C1(new_n192), .C2(new_n194), .ZN(new_n406));
  OAI21_X1  g220(.A(G131), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(new_n202), .A3(new_n243), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n399), .A2(new_n403), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(KEYINPUT71), .A3(new_n396), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n398), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n403), .A2(KEYINPUT66), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT30), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT66), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n203), .A2(new_n414), .A3(new_n228), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n412), .A2(new_n413), .A3(new_n408), .A4(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT30), .B1(new_n388), .B2(new_n389), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n399), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT31), .B1(new_n411), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n416), .A2(new_n417), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n379), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT31), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n421), .A2(new_n422), .A3(new_n398), .A4(new_n410), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT72), .B(KEYINPUT28), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n408), .B1(new_n389), .B2(new_n414), .ZN(new_n425));
  AOI211_X1 g239(.A(KEYINPUT66), .B(new_n227), .C1(new_n200), .C2(new_n202), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n379), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n424), .B1(new_n427), .B2(new_n409), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n390), .A2(KEYINPUT28), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n397), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n419), .A2(new_n423), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G472), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n432), .A3(new_n291), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT32), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT32), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n431), .A2(new_n435), .A3(new_n432), .A4(new_n291), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT29), .ZN(new_n438));
  INV_X1    g252(.A(new_n428), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT28), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n409), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n397), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n418), .A2(new_n396), .A3(new_n390), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n438), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT73), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n429), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n441), .A2(KEYINPUT73), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n379), .B1(new_n388), .B2(new_n389), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n409), .A2(new_n448), .ZN(new_n449));
  AOI22_X1  g263(.A1(new_n446), .A2(new_n447), .B1(KEYINPUT28), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n397), .A2(new_n438), .ZN(new_n451));
  AOI21_X1  g265(.A(G902), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n444), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G472), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n357), .B1(new_n437), .B2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT9), .B(G234), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n336), .B1(new_n457), .B2(new_n291), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(G110), .B(G122), .ZN(new_n460));
  INV_X1    g274(.A(new_n216), .ZN(new_n461));
  INV_X1    g275(.A(new_n217), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n462), .A3(new_n214), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(new_n379), .A3(new_n230), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n364), .A2(KEYINPUT5), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n368), .A2(G119), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT5), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n359), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT86), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT86), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n465), .A2(new_n471), .A3(new_n468), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n373), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n474), .A3(new_n237), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n460), .B1(new_n464), .B2(new_n475), .ZN(new_n476));
  OR2_X1    g290(.A1(new_n476), .A2(KEYINPUT6), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n376), .B1(new_n375), .B2(new_n377), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n230), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n475), .B(new_n460), .C1(new_n480), .C2(new_n218), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT87), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n464), .A2(KEYINPUT87), .A3(new_n475), .A4(new_n460), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n476), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n477), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n227), .A2(new_n323), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n488), .B1(new_n323), .B2(new_n243), .ZN(new_n489));
  INV_X1    g303(.A(G224), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(G953), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n489), .B(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(G210), .B1(G237), .B2(G902), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n473), .A2(new_n238), .A3(new_n474), .ZN(new_n495));
  INV_X1    g309(.A(new_n469), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n237), .B1(new_n373), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n460), .B(KEYINPUT8), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  OR2_X1    g313(.A1(new_n499), .A2(KEYINPUT88), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(KEYINPUT88), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT89), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n489), .B1(new_n502), .B2(KEYINPUT7), .ZN(new_n503));
  INV_X1    g317(.A(new_n491), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT7), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g320(.A(KEYINPUT7), .B(new_n504), .C1(new_n489), .C2(new_n502), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n500), .A2(new_n501), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n483), .A2(new_n484), .ZN(new_n509));
  AOI21_X1  g323(.A(G902), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n493), .A2(new_n494), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n494), .B1(new_n493), .B2(new_n510), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(G214), .B1(G237), .B2(G902), .ZN(new_n514));
  XOR2_X1   g328(.A(new_n514), .B(KEYINPUT85), .Z(new_n515));
  INV_X1    g329(.A(G475), .ZN(new_n516));
  AOI21_X1  g330(.A(G143), .B1(new_n392), .B2(G214), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n392), .A2(G143), .A3(G214), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT18), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n518), .B(new_n519), .C1(new_n520), .C2(new_n201), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n322), .A2(new_n324), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(G146), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n333), .ZN(new_n524));
  INV_X1    g338(.A(new_n519), .ZN(new_n525));
  OAI21_X1  g339(.A(G131), .B1(new_n525), .B2(new_n517), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n521), .B(new_n524), .C1(new_n526), .C2(new_n520), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n518), .A2(new_n201), .A3(new_n519), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(KEYINPUT17), .ZN(new_n530));
  INV_X1    g344(.A(new_n329), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n531), .B(new_n327), .C1(new_n526), .C2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n527), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(G113), .B(G122), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT92), .B(G104), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n537), .B(new_n527), .C1(new_n530), .C2(new_n533), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n516), .B1(new_n541), .B2(new_n291), .ZN(new_n542));
  NOR2_X1   g356(.A1(G475), .A2(G902), .ZN(new_n543));
  XOR2_X1   g357(.A(new_n543), .B(KEYINPUT94), .Z(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT19), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n522), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n332), .A2(KEYINPUT19), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n219), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT91), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n550), .A3(new_n327), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n522), .A2(new_n546), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n332), .A2(KEYINPUT19), .ZN(new_n553));
  AOI21_X1  g367(.A(G146), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT91), .B1(new_n554), .B2(new_n328), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n551), .A2(new_n555), .A3(new_n529), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n527), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(KEYINPUT93), .A3(new_n538), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n540), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n537), .B1(new_n556), .B2(new_n527), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n560), .A2(KEYINPUT93), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n545), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  XOR2_X1   g376(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n540), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(KEYINPUT93), .B2(new_n560), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n557), .A2(new_n538), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT93), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT20), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n572), .A3(new_n545), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n542), .B1(new_n565), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(G478), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(KEYINPUT15), .ZN(new_n576));
  INV_X1    g390(.A(G122), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(G116), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n368), .A2(G122), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(KEYINPUT14), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n581), .A3(G107), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n578), .B(new_n579), .C1(KEYINPUT14), .C2(new_n205), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT95), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n221), .A2(G128), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n315), .A2(G143), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n586), .A2(new_n587), .A3(new_n585), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(G134), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n590), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n385), .B1(new_n592), .B2(new_n588), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n584), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(G116), .B(G122), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(new_n205), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT13), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n586), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n587), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n586), .A2(new_n597), .ZN(new_n600));
  OAI21_X1  g414(.A(G134), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n593), .A2(new_n596), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT96), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT96), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n593), .A2(new_n596), .A3(new_n601), .A4(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n594), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n457), .A2(G217), .A3(new_n262), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  AOI211_X1 g423(.A(new_n594), .B(new_n607), .C1(new_n603), .C2(new_n605), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n291), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT97), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n576), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OR2_X1    g427(.A1(new_n606), .A2(new_n608), .ZN(new_n614));
  INV_X1    g428(.A(new_n610), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n576), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n616), .A2(KEYINPUT97), .A3(new_n291), .A4(new_n617), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n262), .A2(G952), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(G234), .B2(G237), .ZN(new_n621));
  NAND2_X1  g435(.A1(G234), .A2(G237), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(G902), .A3(G953), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n623), .B(KEYINPUT98), .Z(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT21), .B(G898), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n574), .A2(new_n619), .A3(new_n627), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n513), .A2(new_n515), .A3(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n310), .A2(new_n455), .A3(new_n459), .A4(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G101), .ZN(G3));
  NAND3_X1  g445(.A1(new_n305), .A2(KEYINPUT84), .A3(G469), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n308), .B1(new_n307), .B2(new_n290), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n458), .B1(new_n634), .B2(new_n292), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n431), .A2(new_n291), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G472), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n637), .A2(new_n433), .A3(new_n356), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n515), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n641), .B(new_n627), .C1(new_n511), .C2(new_n512), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT33), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n614), .B(new_n615), .C1(KEYINPUT99), .C2(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(KEYINPUT99), .B1(new_n606), .B2(new_n608), .ZN(new_n645));
  OAI211_X1 g459(.A(new_n645), .B(KEYINPUT33), .C1(new_n609), .C2(new_n610), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n575), .A2(G902), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(KEYINPUT100), .A3(new_n648), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT100), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n611), .B2(new_n575), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n649), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n574), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n642), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n640), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT34), .B(G104), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G6));
  AOI21_X1  g473(.A(new_n542), .B1(new_n613), .B2(new_n618), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n571), .A2(new_n545), .A3(new_n563), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n565), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n642), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n640), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT35), .B(G107), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  NAND2_X1  g481(.A1(new_n330), .A2(new_n334), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n339), .A2(KEYINPUT36), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n355), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n671), .B1(new_n348), .B2(new_n351), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n637), .A2(new_n433), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT101), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n637), .A2(KEYINPUT101), .A3(new_n433), .A4(new_n672), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n310), .A2(new_n459), .A3(new_n629), .A4(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT102), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n680), .B(KEYINPUT103), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n678), .B(new_n681), .ZN(G12));
  AOI22_X1  g496(.A1(new_n434), .A2(new_n436), .B1(new_n453), .B2(G472), .ZN(new_n683));
  INV_X1    g497(.A(G900), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n624), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n621), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n660), .A2(new_n662), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n660), .A2(new_n662), .A3(KEYINPUT104), .A4(new_n687), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n641), .B(new_n672), .C1(new_n511), .C2(new_n512), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n683), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n310), .A2(new_n694), .A3(new_n459), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT105), .B(G128), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G30));
  XOR2_X1   g511(.A(new_n513), .B(KEYINPUT38), .Z(new_n698));
  NOR2_X1   g512(.A1(new_n411), .A2(new_n418), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n397), .B2(new_n449), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n700), .B2(G902), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n437), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n565), .A2(new_n573), .ZN(new_n703));
  INV_X1    g517(.A(new_n542), .ZN(new_n704));
  AOI22_X1  g518(.A1(new_n703), .A2(new_n704), .B1(new_n618), .B2(new_n613), .ZN(new_n705));
  INV_X1    g519(.A(new_n672), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n641), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT106), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n698), .A2(new_n702), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n687), .B(KEYINPUT39), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n635), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n709), .B1(new_n711), .B2(KEYINPUT40), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n712), .B1(KEYINPUT40), .B2(new_n711), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G143), .ZN(G45));
  NAND3_X1  g528(.A1(new_n653), .A2(new_n654), .A3(new_n687), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n683), .A2(new_n693), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n310), .A2(new_n459), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  AND3_X1   g532(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n290), .B1(new_n289), .B2(new_n291), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n719), .A2(new_n720), .A3(new_n458), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n455), .A3(new_n656), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NOR2_X1   g538(.A1(new_n719), .A2(new_n720), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(new_n664), .A3(new_n455), .A4(new_n459), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G116), .ZN(G18));
  NOR3_X1   g541(.A1(new_n683), .A2(new_n693), .A3(new_n628), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n721), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  OAI211_X1 g544(.A(new_n705), .B(new_n641), .C1(new_n511), .C2(new_n512), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n419), .B(new_n423), .C1(new_n450), .C2(new_n396), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n432), .A3(new_n291), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n637), .A2(new_n733), .A3(new_n356), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n731), .A2(new_n734), .A3(new_n626), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n721), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G122), .ZN(G24));
  NOR3_X1   g551(.A1(new_n260), .A2(new_n296), .A3(new_n265), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n298), .B1(new_n301), .B2(new_n302), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n738), .B1(new_n739), .B2(new_n265), .ZN(new_n740));
  OAI21_X1  g554(.A(G469), .B1(new_n740), .B2(G902), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n493), .A2(new_n510), .ZN(new_n742));
  INV_X1    g556(.A(new_n494), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n493), .A2(new_n494), .A3(new_n510), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n515), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n741), .A2(new_n746), .A3(new_n459), .A4(new_n292), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n637), .A2(new_n733), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n647), .A2(KEYINPUT100), .A3(new_n648), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n652), .B1(new_n647), .B2(new_n648), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n574), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n748), .A2(new_n752), .A3(new_n672), .A4(new_n687), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n747), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n323), .ZN(G27));
  OAI21_X1  g569(.A(new_n292), .B1(new_n290), .B2(new_n307), .ZN(new_n756));
  INV_X1    g570(.A(new_n715), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n744), .A2(new_n459), .A3(new_n641), .A4(new_n745), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n455), .A2(new_n756), .A3(new_n757), .A4(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT42), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT107), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n437), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n434), .A2(KEYINPUT107), .A3(new_n436), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n454), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n305), .A2(G469), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n758), .B1(new_n767), .B2(new_n292), .ZN(new_n768));
  INV_X1    g582(.A(new_n687), .ZN(new_n769));
  NOR4_X1   g583(.A1(new_n751), .A2(new_n761), .A3(new_n574), .A4(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n766), .A2(new_n768), .A3(new_n356), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n762), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G131), .ZN(G33));
  AND2_X1   g587(.A1(new_n690), .A2(new_n691), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n455), .A2(new_n756), .A3(new_n774), .A4(new_n759), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G134), .ZN(G36));
  INV_X1    g590(.A(KEYINPUT109), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT43), .B1(new_n574), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n778), .B1(new_n751), .B2(new_n654), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n653), .B(new_n574), .C1(new_n777), .C2(KEYINPUT43), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n706), .B1(new_n637), .B2(new_n433), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n781), .A2(KEYINPUT44), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT44), .B1(new_n781), .B2(new_n782), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n511), .A2(new_n512), .A3(new_n515), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n783), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT46), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n304), .A2(KEYINPUT45), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT45), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n300), .A2(new_n303), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n788), .B(G469), .C1(new_n792), .C2(G902), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT108), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT108), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n290), .B1(new_n789), .B2(new_n791), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n290), .A2(new_n291), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n795), .B(new_n788), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n791), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n790), .B1(new_n300), .B2(new_n303), .ZN(new_n800));
  OAI21_X1  g614(.A(G469), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n797), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(KEYINPUT46), .A3(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n794), .A2(new_n292), .A3(new_n798), .A4(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n787), .A2(new_n804), .A3(new_n459), .A4(new_n710), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G137), .ZN(G39));
  NAND2_X1  g620(.A1(new_n437), .A2(new_n454), .ZN(new_n807));
  NOR4_X1   g621(.A1(new_n786), .A2(new_n807), .A3(new_n356), .A4(new_n715), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n804), .A2(KEYINPUT47), .A3(new_n459), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT47), .B1(new_n804), .B2(new_n459), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G140), .ZN(G42));
  NOR2_X1   g627(.A1(new_n458), .A2(new_n515), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n653), .A2(new_n356), .A3(new_n574), .A4(new_n814), .ZN(new_n815));
  XOR2_X1   g629(.A(new_n815), .B(KEYINPUT110), .Z(new_n816));
  INV_X1    g630(.A(KEYINPUT49), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n816), .B1(new_n817), .B2(new_n725), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT111), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  AOI211_X1 g635(.A(new_n702), .B(new_n698), .C1(new_n817), .C2(new_n725), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n823), .B(KEYINPUT112), .Z(new_n824));
  NAND3_X1  g638(.A1(new_n637), .A2(new_n733), .A3(new_n672), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n715), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n721), .A2(new_n746), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n731), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n706), .A2(new_n459), .A3(new_n687), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n756), .A2(new_n828), .A3(new_n702), .A4(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n695), .A2(new_n717), .A3(new_n827), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n754), .B1(new_n635), .B2(new_n694), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n835), .A2(KEYINPUT52), .A3(new_n717), .A4(new_n831), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n542), .A2(new_n769), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n672), .A2(new_n618), .A3(new_n613), .A4(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n563), .B1(new_n571), .B2(new_n545), .ZN(new_n840));
  AOI211_X1 g654(.A(new_n544), .B(new_n564), .C1(new_n567), .C2(new_n570), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n843), .A2(new_n744), .A3(new_n641), .A4(new_n745), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n683), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n310), .A2(new_n459), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n826), .A2(new_n756), .A3(new_n759), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n775), .A3(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n765), .A2(new_n454), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n357), .B1(new_n849), .B2(new_n764), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n756), .A2(new_n759), .A3(new_n770), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n850), .A2(new_n851), .B1(new_n760), .B2(new_n761), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n654), .A2(new_n619), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n642), .B1(new_n655), .B2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n310), .A2(new_n459), .A3(new_n638), .A4(new_n855), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n630), .A2(new_n678), .A3(new_n856), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n722), .A2(new_n729), .A3(new_n736), .A4(new_n726), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n853), .A2(KEYINPUT53), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n837), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n719), .B1(new_n632), .B2(new_n633), .ZN(new_n861));
  INV_X1    g675(.A(new_n844), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n807), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n861), .A2(new_n863), .A3(new_n458), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n775), .A2(new_n847), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n858), .A2(new_n866), .A3(new_n772), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n630), .A2(new_n678), .A3(new_n856), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT113), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n834), .A2(new_n836), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT113), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n853), .A2(new_n871), .A3(new_n857), .A4(new_n858), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n860), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n873), .B(new_n874), .ZN(new_n876));
  MUX2_X1   g690(.A(new_n875), .B(new_n876), .S(KEYINPUT54), .Z(new_n877));
  AOI21_X1  g691(.A(new_n686), .B1(new_n779), .B2(new_n780), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n850), .A2(new_n725), .A3(new_n759), .A4(new_n878), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n879), .A2(KEYINPUT116), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(KEYINPUT116), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(KEYINPUT48), .A3(new_n881), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n620), .B(KEYINPUT115), .Z(new_n883));
  NAND3_X1  g697(.A1(new_n878), .A2(new_n356), .A3(new_n748), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n884), .A2(new_n747), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n725), .A2(new_n759), .ZN(new_n886));
  NOR4_X1   g700(.A1(new_n886), .A2(new_n357), .A3(new_n686), .A4(new_n702), .ZN(new_n887));
  AOI211_X1 g701(.A(new_n883), .B(new_n885), .C1(new_n887), .C2(new_n752), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT48), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n879), .A2(KEYINPUT116), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n882), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n884), .A2(new_n786), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n810), .A2(new_n811), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n725), .A2(new_n458), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n892), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n878), .A2(new_n725), .A3(new_n759), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n897), .A2(new_n825), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n653), .A2(new_n654), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n898), .B1(new_n887), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n721), .ZN(new_n901));
  NOR4_X1   g715(.A1(new_n698), .A2(new_n884), .A3(new_n901), .A4(new_n641), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n902), .A2(KEYINPUT50), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(KEYINPUT50), .ZN(new_n904));
  OAI211_X1 g718(.A(KEYINPUT51), .B(new_n900), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n891), .B1(new_n896), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n893), .A2(KEYINPUT114), .ZN(new_n909));
  OR3_X1    g723(.A1(new_n810), .A2(KEYINPUT114), .A3(new_n811), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n909), .A2(new_n910), .A3(new_n894), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n908), .B1(new_n911), .B2(new_n892), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n907), .B1(new_n912), .B2(KEYINPUT51), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n877), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(G952), .A2(G953), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n824), .B1(new_n914), .B2(new_n915), .ZN(G75));
  NOR2_X1   g730(.A1(new_n262), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n875), .A2(new_n291), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT56), .B1(new_n919), .B2(G210), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n487), .B(new_n492), .Z(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT55), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n918), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n923), .B1(new_n920), .B2(new_n922), .ZN(G51));
  XNOR2_X1  g738(.A(new_n875), .B(KEYINPUT54), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n797), .B(KEYINPUT117), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT57), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n289), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n919), .A2(new_n796), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n917), .B1(new_n928), .B2(new_n929), .ZN(G54));
  AND2_X1   g744(.A1(KEYINPUT58), .A2(G475), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n919), .A2(new_n571), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n571), .B1(new_n919), .B2(new_n931), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n932), .A2(new_n933), .A3(new_n917), .ZN(G60));
  NAND2_X1  g748(.A1(G478), .A2(G902), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT59), .Z(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n647), .B1(new_n877), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n647), .A2(new_n937), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n918), .B1(new_n925), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n938), .A2(new_n940), .ZN(G63));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT60), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n353), .B1(new_n875), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT119), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n875), .A2(new_n943), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n670), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n944), .A2(new_n945), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n918), .A2(KEYINPUT61), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n946), .A2(new_n948), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT118), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n944), .A2(new_n952), .A3(new_n918), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n944), .B2(new_n918), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n947), .A2(new_n670), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n951), .B1(new_n956), .B2(KEYINPUT61), .ZN(G66));
  NAND2_X1  g771(.A1(new_n857), .A2(new_n858), .ZN(new_n958));
  NAND2_X1  g772(.A1(G224), .A2(G953), .ZN(new_n959));
  OAI22_X1  g773(.A1(new_n958), .A2(G953), .B1(new_n625), .B2(new_n959), .ZN(new_n960));
  OAI221_X1 g774(.A(new_n477), .B1(G898), .B2(new_n262), .C1(new_n485), .C2(new_n486), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n960), .B(new_n961), .Z(G69));
  NAND2_X1  g776(.A1(new_n552), .A2(new_n553), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT120), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n420), .B(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n854), .A2(new_n655), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n455), .A2(new_n785), .A3(new_n966), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n711), .A2(new_n967), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n805), .A2(new_n968), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n835), .A2(new_n717), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n713), .A2(KEYINPUT62), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(KEYINPUT62), .B1(new_n713), .B2(new_n970), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n812), .B(new_n969), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n965), .B1(new_n974), .B2(G953), .ZN(new_n975));
  INV_X1    g789(.A(new_n965), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n262), .A2(G900), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT122), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n798), .A2(new_n292), .A3(new_n803), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n458), .B1(new_n979), .B2(new_n794), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT123), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n766), .A2(new_n356), .A3(new_n828), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n980), .A2(new_n981), .A3(new_n710), .A4(new_n983), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n804), .A2(new_n459), .A3(new_n710), .A4(new_n983), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(KEYINPUT123), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n775), .ZN(new_n988));
  OR3_X1    g802(.A1(new_n852), .A2(KEYINPUT124), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(KEYINPUT124), .B1(new_n852), .B2(new_n988), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n805), .A2(new_n970), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n987), .A2(new_n812), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n978), .B1(new_n993), .B2(new_n262), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n976), .B1(new_n994), .B2(KEYINPUT125), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT125), .ZN(new_n996));
  AOI211_X1 g810(.A(new_n996), .B(new_n978), .C1(new_n993), .C2(new_n262), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n975), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT121), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n999), .B1(new_n995), .B2(new_n997), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n262), .B1(G227), .B2(G900), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n998), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  OAI221_X1 g817(.A(new_n975), .B1(new_n999), .B2(new_n1001), .C1(new_n995), .C2(new_n997), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n1003), .A2(new_n1004), .ZN(G72));
  NAND2_X1  g819(.A1(G472), .A2(G902), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT63), .Z(new_n1007));
  NOR2_X1   g821(.A1(new_n418), .A2(new_n390), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1008), .A2(new_n396), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1007), .B1(new_n1009), .B2(new_n699), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1010), .B(KEYINPUT126), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n876), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT127), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1007), .B1(new_n973), .B2(new_n958), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n1014), .B(new_n396), .C1(new_n418), .C2(new_n390), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1007), .B1(new_n993), .B2(new_n958), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n443), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1015), .A2(new_n918), .A3(new_n1017), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1013), .A2(new_n1018), .ZN(G57));
endmodule


