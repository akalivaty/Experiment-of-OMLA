//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n449, new_n451, new_n453, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n631, new_n632,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1202,
    new_n1203;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G108), .Z(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT66), .Z(G173));
  XNOR2_X1  g022(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT68), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NOR4_X1   g031(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT69), .Z(new_n462));
  INV_X1    g037(.A(new_n456), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2106), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n471));
  AND3_X1   g046(.A1(new_n469), .A2(new_n471), .A3(KEYINPUT70), .ZN(new_n472));
  AOI21_X1  g047(.A(KEYINPUT70), .B1(new_n469), .B2(new_n471), .ZN(new_n473));
  OAI21_X1  g048(.A(G125), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n467), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n470), .A2(KEYINPUT71), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT71), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n480), .A2(G101), .A3(new_n467), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT72), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(G2105), .B1(new_n477), .B2(new_n479), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(KEYINPUT72), .A3(G101), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n477), .A2(new_n479), .A3(KEYINPUT3), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n486), .A2(G137), .A3(new_n467), .A4(new_n469), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n476), .A2(new_n488), .ZN(G160));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n469), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(new_n467), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n492), .B(KEYINPUT73), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n490), .A2(G2105), .ZN(new_n494));
  MUX2_X1   g069(.A(G100), .B(G112), .S(G2105), .Z(new_n495));
  AOI22_X1  g070(.A1(new_n494), .A2(G136), .B1(G2104), .B2(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n493), .A2(new_n496), .ZN(G162));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  AND2_X1   g073(.A1(KEYINPUT74), .A2(G114), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT74), .A2(G114), .ZN(new_n500));
  OAI21_X1  g075(.A(G2105), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT75), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT75), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n503), .B(G2105), .C1(new_n499), .C2(new_n500), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n498), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n486), .A2(G126), .A3(G2105), .A4(new_n469), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n486), .A2(G138), .A3(new_n467), .A4(new_n469), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT4), .ZN(new_n510));
  INV_X1    g085(.A(G138), .ZN(new_n511));
  NOR3_X1   g086(.A1(new_n511), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n512), .B1(new_n472), .B2(new_n473), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT76), .A2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(KEYINPUT76), .A2(KEYINPUT5), .A3(G543), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G62), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n517), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT77), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n524), .A2(new_n525), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n520), .A2(new_n521), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n527), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G651), .ZN(new_n529));
  OAI21_X1  g104(.A(KEYINPUT77), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(KEYINPUT6), .A2(G651), .ZN(new_n532));
  NOR2_X1   g107(.A1(KEYINPUT6), .A2(G651), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n522), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n519), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n535), .A2(G88), .B1(G50), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n531), .A2(new_n537), .ZN(G303));
  INV_X1    g113(.A(G303), .ZN(G166));
  AND2_X1   g114(.A1(new_n535), .A2(G89), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT7), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n527), .A2(G63), .A3(G651), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n532), .A2(new_n533), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G51), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n542), .B(new_n543), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n540), .A2(new_n547), .ZN(G168));
  INV_X1    g123(.A(G52), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n544), .A2(new_n527), .ZN(new_n550));
  INV_X1    g125(.A(G90), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n549), .A2(new_n545), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n529), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n552), .A2(new_n554), .ZN(G171));
  AOI22_X1  g130(.A1(new_n527), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(new_n529), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n536), .A2(G43), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT79), .ZN(new_n559));
  XOR2_X1   g134(.A(KEYINPUT78), .B(G81), .Z(new_n560));
  OAI211_X1 g135(.A(new_n558), .B(new_n559), .C1(new_n550), .C2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  OR3_X1    g137(.A1(new_n522), .A2(new_n560), .A3(new_n534), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n559), .B1(new_n563), .B2(new_n558), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n557), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(KEYINPUT80), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT80), .ZN(new_n567));
  OAI211_X1 g142(.A(new_n567), .B(new_n557), .C1(new_n562), .C2(new_n564), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  AND3_X1   g145(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G36), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(G188));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G65), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n522), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(G651), .B1(new_n535), .B2(G91), .ZN(new_n579));
  INV_X1    g154(.A(G53), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT9), .B1(new_n545), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT9), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n536), .A2(new_n582), .A3(G53), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n579), .A2(new_n584), .ZN(G299));
  INV_X1    g160(.A(G171), .ZN(G301));
  INV_X1    g161(.A(G168), .ZN(G286));
  NAND2_X1  g162(.A1(new_n535), .A2(G87), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n536), .A2(G49), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G288));
  AOI22_X1  g166(.A1(new_n535), .A2(G86), .B1(G48), .B2(new_n536), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT81), .ZN(new_n594));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n520), .B2(new_n521), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(KEYINPUT82), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT82), .ZN(new_n599));
  OAI211_X1 g174(.A(new_n599), .B(G651), .C1(new_n594), .C2(new_n596), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n592), .A2(new_n598), .A3(new_n600), .ZN(G305));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  XNOR2_X1  g177(.A(KEYINPUT85), .B(G47), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n602), .A2(new_n550), .B1(new_n545), .B2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G60), .ZN(new_n606));
  INV_X1    g181(.A(G72), .ZN(new_n607));
  OAI22_X1  g182(.A1(new_n522), .A2(new_n606), .B1(new_n607), .B2(new_n519), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(KEYINPUT83), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT83), .ZN(new_n610));
  OAI221_X1 g185(.A(new_n610), .B1(new_n607), .B2(new_n519), .C1(new_n522), .C2(new_n606), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n609), .A2(G651), .A3(new_n611), .ZN(new_n612));
  AND2_X1   g187(.A1(new_n612), .A2(KEYINPUT84), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n612), .A2(KEYINPUT84), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n605), .B1(new_n613), .B2(new_n614), .ZN(G290));
  XOR2_X1   g190(.A(KEYINPUT86), .B(KEYINPUT10), .Z(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n535), .A2(G92), .A3(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G92), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n616), .B1(new_n550), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(G79), .A2(G543), .ZN(new_n622));
  INV_X1    g197(.A(G66), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n522), .B2(new_n623), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n624), .A2(G651), .B1(new_n536), .B2(G54), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  MUX2_X1   g201(.A(new_n626), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g202(.A(new_n626), .B(G301), .S(G868), .Z(G321));
  MUX2_X1   g203(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g204(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g205(.A(new_n626), .ZN(new_n631));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(G860), .ZN(G148));
  INV_X1    g208(.A(G868), .ZN(new_n634));
  NOR3_X1   g209(.A1(new_n626), .A2(G559), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n569), .B2(new_n634), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n469), .A2(new_n471), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT70), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n469), .A2(new_n471), .A3(KEYINPUT70), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(new_n484), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT12), .ZN(new_n644));
  INV_X1    g219(.A(G2100), .ZN(new_n645));
  AOI22_X1  g220(.A1(new_n644), .A2(KEYINPUT13), .B1(KEYINPUT87), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(KEYINPUT13), .B2(new_n644), .ZN(new_n647));
  OR3_X1    g222(.A1(new_n647), .A2(KEYINPUT87), .A3(new_n645), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n647), .B1(KEYINPUT87), .B2(new_n645), .ZN(new_n649));
  MUX2_X1   g224(.A(G99), .B(G111), .S(G2105), .Z(new_n650));
  AOI22_X1  g225(.A1(new_n491), .A2(G123), .B1(G2104), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n494), .A2(G135), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(G2096), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n648), .A2(new_n649), .A3(new_n655), .ZN(G156));
  INV_X1    g231(.A(KEYINPUT14), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT15), .B(G2435), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2427), .ZN(new_n660));
  INV_X1    g235(.A(G2430), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n657), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n661), .B2(new_n660), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2451), .B(G2454), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT16), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1341), .B(G1348), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n663), .A2(new_n669), .ZN(new_n671));
  AND3_X1   g246(.A1(new_n670), .A2(G14), .A3(new_n671), .ZN(G401));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT88), .ZN(new_n674));
  NOR2_X1   g249(.A1(G2072), .A2(G2078), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n442), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2084), .B(G2090), .Z(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n676), .B(KEYINPUT17), .Z(new_n681));
  OAI211_X1 g256(.A(new_n678), .B(new_n680), .C1(new_n681), .C2(new_n674), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n681), .A2(new_n674), .A3(new_n679), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n676), .A2(new_n679), .A3(new_n673), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT18), .Z(new_n685));
  NAND3_X1  g260(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(new_n654), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G2100), .ZN(G227));
  XNOR2_X1  g263(.A(G1956), .B(G2474), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT89), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1961), .B(G1966), .Z(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1971), .B(G1976), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT19), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n691), .A2(new_n692), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n693), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n697), .A2(KEYINPUT90), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(KEYINPUT90), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n695), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT91), .B(KEYINPUT20), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n696), .B(new_n698), .C1(new_n701), .C2(new_n703), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n701), .A2(new_n703), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1991), .B(G1996), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n708), .B(new_n709), .Z(new_n710));
  XNOR2_X1  g285(.A(G1981), .B(G1986), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT92), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n708), .B(new_n709), .ZN(new_n714));
  INV_X1    g289(.A(new_n712), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n713), .A2(new_n716), .ZN(G229));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n569), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n718), .B2(G19), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G1341), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G33), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT25), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n642), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n726), .A2(new_n467), .ZN(new_n727));
  AOI211_X1 g302(.A(new_n725), .B(new_n727), .C1(G139), .C2(new_n494), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n723), .B1(new_n728), .B2(new_n722), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G2072), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n718), .A2(G5), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G171), .B2(new_n718), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n732), .A2(G1961), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(G1961), .ZN(new_n734));
  NOR2_X1   g309(.A1(G168), .A2(new_n718), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n718), .B2(G21), .ZN(new_n736));
  INV_X1    g311(.A(G1966), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n733), .B(new_n734), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n722), .A2(G32), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n494), .A2(G141), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n491), .A2(G129), .ZN(new_n741));
  NAND3_X1  g316(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT26), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  AOI22_X1  g320(.A1(G105), .A2(new_n484), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n740), .A2(new_n741), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n739), .B1(new_n748), .B2(new_n722), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT27), .B(G1996), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT24), .B(G34), .Z(new_n752));
  NOR2_X1   g327(.A1(new_n752), .A2(G29), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G160), .B2(G29), .ZN(new_n754));
  NOR2_X1   g329(.A1(G4), .A2(G16), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n631), .B2(G16), .ZN(new_n756));
  OAI221_X1 g331(.A(new_n751), .B1(G2084), .B2(new_n754), .C1(G1348), .C2(new_n756), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT31), .B(G11), .Z(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT30), .B(G28), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n758), .B1(new_n722), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n653), .B2(new_n722), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n736), .B2(new_n737), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n756), .A2(G1348), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n749), .A2(new_n750), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n754), .A2(G2084), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n762), .A2(new_n763), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  NOR4_X1   g341(.A1(new_n730), .A2(new_n738), .A3(new_n757), .A4(new_n766), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n721), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(G162), .A2(G29), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G29), .B2(G35), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT29), .ZN(new_n771));
  INV_X1    g346(.A(G2090), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n718), .A2(G20), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT23), .Z(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G299), .B2(G16), .ZN(new_n776));
  INV_X1    g351(.A(G1956), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G27), .A2(G29), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G164), .B2(G29), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G2078), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n773), .A2(new_n778), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n771), .A2(new_n772), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT100), .B(KEYINPUT28), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n722), .A2(G26), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n494), .A2(G140), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n491), .A2(G128), .ZN(new_n788));
  OAI21_X1  g363(.A(KEYINPUT98), .B1(G104), .B2(G2105), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NOR3_X1   g365(.A1(KEYINPUT98), .A2(G104), .A3(G2105), .ZN(new_n791));
  OAI221_X1 g366(.A(G2104), .B1(G116), .B2(new_n467), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n787), .A2(new_n788), .A3(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT99), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n787), .A2(new_n788), .A3(KEYINPUT99), .A4(new_n792), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n786), .B1(new_n797), .B2(G29), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2067), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n768), .A2(new_n782), .A3(new_n783), .A4(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT36), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n491), .A2(G119), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT93), .ZN(new_n803));
  MUX2_X1   g378(.A(G95), .B(G107), .S(G2105), .Z(new_n804));
  AOI22_X1  g379(.A1(new_n494), .A2(G131), .B1(G2104), .B2(new_n804), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(G29), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G25), .B2(G29), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT94), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT35), .B(G1991), .Z(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT94), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n808), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(new_n810), .ZN(new_n815));
  NOR2_X1   g390(.A1(G16), .A2(G24), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n612), .A2(KEYINPUT84), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n612), .A2(KEYINPUT84), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n604), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n816), .B1(new_n819), .B2(G16), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(G1986), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(G1986), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n812), .A2(new_n815), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n718), .A2(G22), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT96), .Z(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G166), .B2(new_n718), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT97), .B(G1971), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n826), .B(new_n827), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n718), .A2(G23), .ZN(new_n829));
  INV_X1    g404(.A(G288), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(new_n718), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT33), .B(G1976), .Z(new_n832));
  XOR2_X1   g407(.A(new_n831), .B(new_n832), .Z(new_n833));
  MUX2_X1   g408(.A(G6), .B(G305), .S(G16), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT95), .ZN(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT32), .B(G1981), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n828), .B(new_n833), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n839), .A2(KEYINPUT34), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n823), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(KEYINPUT34), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n801), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n841), .A2(new_n801), .A3(new_n842), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n800), .B1(new_n844), .B2(new_n845), .ZN(G311));
  INV_X1    g421(.A(new_n800), .ZN(new_n847));
  INV_X1    g422(.A(new_n845), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(new_n848), .B2(new_n843), .ZN(G150));
  AOI22_X1  g424(.A1(new_n535), .A2(G93), .B1(G55), .B2(new_n536), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n527), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n850), .B1(new_n529), .B2(new_n851), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(KEYINPUT101), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(KEYINPUT101), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(G860), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  NAND3_X1  g432(.A1(new_n566), .A2(new_n568), .A3(new_n852), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n853), .A2(new_n565), .A3(new_n854), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT38), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n631), .A2(G559), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n864));
  INV_X1    g439(.A(G860), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(new_n863), .B2(KEYINPUT39), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n857), .B1(new_n864), .B2(new_n866), .ZN(G145));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n728), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n728), .A2(new_n868), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n795), .A2(G164), .A3(new_n796), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(G164), .B1(new_n795), .B2(new_n796), .ZN(new_n873));
  NOR3_X1   g448(.A1(new_n872), .A2(new_n873), .A3(new_n748), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n797), .A2(new_n515), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n747), .B1(new_n875), .B2(new_n871), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n869), .B(new_n870), .C1(new_n874), .C2(new_n876), .ZN(new_n877));
  MUX2_X1   g452(.A(G106), .B(G118), .S(G2105), .Z(new_n878));
  AOI22_X1  g453(.A1(new_n491), .A2(G130), .B1(G2104), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n494), .A2(G142), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n644), .B(new_n881), .Z(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n806), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n748), .B1(new_n872), .B2(new_n873), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n875), .A2(new_n747), .A3(new_n871), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n884), .A2(new_n885), .A3(new_n868), .A4(new_n728), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n877), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n877), .A2(new_n883), .A3(KEYINPUT103), .A4(new_n886), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n877), .A2(new_n886), .ZN(new_n891));
  INV_X1    g466(.A(new_n883), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n889), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n653), .B(G160), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(G162), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(G37), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n883), .B1(new_n877), .B2(new_n886), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n900), .A2(new_n896), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n899), .B1(new_n901), .B2(new_n887), .ZN(new_n902));
  INV_X1    g477(.A(new_n887), .ZN(new_n903));
  NOR4_X1   g478(.A1(new_n903), .A2(new_n900), .A3(KEYINPUT104), .A4(new_n896), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n897), .B(new_n898), .C1(new_n902), .C2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g481(.A1(new_n855), .A2(G868), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n626), .A2(G559), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n860), .B(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n626), .A2(G299), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n621), .A2(new_n579), .A3(new_n584), .A4(new_n625), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n912), .ZN(new_n914));
  XNOR2_X1  g489(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  AOI22_X1  g491(.A1(new_n913), .A2(KEYINPUT106), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n914), .A2(KEYINPUT106), .A3(new_n916), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n909), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n910), .A2(new_n912), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n909), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n819), .A2(new_n830), .ZN(new_n925));
  NAND2_X1  g500(.A1(G290), .A2(G288), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XOR2_X1   g502(.A(G303), .B(G305), .Z(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n932), .B1(new_n933), .B2(KEYINPUT42), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n924), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n934), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(new_n921), .A3(new_n923), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n933), .A2(KEYINPUT42), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n935), .A2(new_n933), .A3(new_n937), .A4(KEYINPUT42), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n907), .B1(new_n942), .B2(G868), .ZN(G295));
  AOI21_X1  g518(.A(new_n907), .B1(new_n942), .B2(G868), .ZN(G331));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n945));
  XNOR2_X1  g520(.A(G168), .B(G171), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n858), .A2(new_n859), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n946), .B1(new_n858), .B2(new_n859), .ZN(new_n948));
  OAI22_X1  g523(.A1(new_n947), .A2(new_n948), .B1(new_n919), .B2(new_n917), .ZN(new_n949));
  INV_X1    g524(.A(new_n946), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n860), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n858), .A2(new_n859), .A3(new_n946), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n922), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n949), .A2(new_n932), .A3(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n954), .A2(new_n898), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT108), .B1(new_n922), .B2(new_n911), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n914), .A2(new_n957), .A3(KEYINPUT41), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n922), .A2(new_n915), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(new_n947), .B2(new_n948), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n947), .A2(new_n948), .ZN(new_n962));
  AOI22_X1  g537(.A1(new_n961), .A2(KEYINPUT109), .B1(new_n962), .B2(new_n922), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n960), .B(new_n964), .C1(new_n947), .C2(new_n948), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n932), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n955), .B1(new_n966), .B2(KEYINPUT110), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT110), .ZN(new_n968));
  AOI211_X1 g543(.A(new_n968), .B(new_n932), .C1(new_n963), .C2(new_n965), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n945), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n930), .A2(new_n931), .ZN(new_n972));
  INV_X1    g547(.A(new_n917), .ZN(new_n973));
  AOI22_X1  g548(.A1(new_n951), .A2(new_n952), .B1(new_n973), .B2(new_n918), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n947), .A2(new_n948), .A3(new_n914), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n955), .A2(KEYINPUT43), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n970), .A2(new_n971), .A3(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n976), .A2(new_n945), .A3(new_n898), .A4(new_n954), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n979), .A2(KEYINPUT111), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT44), .B1(new_n979), .B2(KEYINPUT111), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT43), .B1(new_n967), .B2(new_n969), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n978), .A2(new_n984), .ZN(G397));
  INV_X1    g560(.A(KEYINPUT62), .ZN(new_n986));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  INV_X1    g562(.A(new_n498), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT74), .B(G114), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n503), .B1(new_n989), .B2(G2105), .ZN(new_n990));
  INV_X1    g565(.A(new_n504), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n506), .ZN(new_n993));
  AOI22_X1  g568(.A1(new_n642), .A2(new_n512), .B1(new_n509), .B2(KEYINPUT4), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n987), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G40), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n476), .A2(new_n488), .A3(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(KEYINPUT45), .B(new_n987), .C1(new_n993), .C2(new_n994), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n737), .ZN(new_n1002));
  INV_X1    g577(.A(G2084), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT50), .B1(new_n515), .B2(new_n987), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n1005));
  AOI211_X1 g580(.A(new_n1005), .B(G1384), .C1(new_n508), .C2(new_n514), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1003), .B(new_n999), .C1(new_n1004), .C2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1002), .A2(G168), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(G8), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT51), .ZN(new_n1010));
  AOI21_X1  g585(.A(G168), .B1(new_n1002), .B2(new_n1007), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n1012));
  OAI211_X1 g587(.A(G8), .B(new_n1008), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT121), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1010), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1014), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n986), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT121), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1010), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(KEYINPUT62), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(G303), .A2(G8), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1022), .B(KEYINPUT55), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n483), .A2(new_n487), .A3(new_n485), .ZN(new_n1024));
  INV_X1    g599(.A(G125), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n640), .B2(new_n641), .ZN(new_n1026));
  INV_X1    g601(.A(new_n475), .ZN(new_n1027));
  OAI21_X1  g602(.A(G2105), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1024), .A2(new_n1028), .A3(G40), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n995), .A2(new_n1005), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n515), .A2(KEYINPUT50), .A3(new_n987), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT114), .B(G1971), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n772), .A2(new_n1032), .B1(new_n1001), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G8), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1023), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1034), .A2(new_n1035), .A3(new_n1023), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1036), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n995), .A2(new_n1029), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(new_n1035), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n999), .A2(new_n987), .A3(new_n515), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(KEYINPUT115), .A3(G8), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n598), .A2(new_n600), .A3(KEYINPUT116), .ZN(new_n1046));
  AOI21_X1  g621(.A(G305), .B1(G1981), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(G305), .A2(new_n1046), .A3(G1981), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(KEYINPUT49), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT49), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1049), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1051), .B1(new_n1052), .B2(new_n1047), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1045), .A2(new_n1050), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n830), .A2(G1976), .ZN(new_n1055));
  INV_X1    g630(.A(G1976), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT52), .B1(G288), .B2(new_n1056), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1041), .A2(new_n1040), .A3(new_n1035), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT115), .B1(new_n1043), .B2(G8), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1055), .B(new_n1057), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1054), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(new_n1045), .B2(new_n1055), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g639(.A(KEYINPUT117), .B(new_n1023), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT45), .B1(new_n515), .B2(new_n987), .ZN(new_n1066));
  AOI211_X1 g641(.A(new_n996), .B(G1384), .C1(new_n508), .C2(new_n514), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G2078), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1068), .A2(KEYINPUT53), .A3(new_n1069), .A4(new_n999), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n999), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1071));
  INV_X1    g646(.A(G1961), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n997), .A2(new_n1069), .A3(new_n999), .A4(new_n1000), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1070), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G171), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  AND4_X1   g654(.A1(new_n1039), .A2(new_n1064), .A3(new_n1065), .A4(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1017), .A2(new_n1021), .A3(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n626), .A2(KEYINPUT60), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n995), .A2(new_n1029), .A3(G2067), .ZN(new_n1084));
  INV_X1    g659(.A(G1348), .ZN(new_n1085));
  AOI211_X1 g660(.A(new_n1083), .B(new_n1084), .C1(new_n1071), .C2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1996), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n997), .A2(new_n1087), .A3(new_n999), .A4(new_n1000), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT58), .B(G1341), .Z(new_n1089));
  NAND2_X1  g664(.A1(new_n1043), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n569), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(new_n569), .A3(new_n1093), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1086), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT61), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT57), .B1(new_n584), .B2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n1100), .B(G299), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1071), .A2(new_n777), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT56), .B(G2072), .Z(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .A4(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1101), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1101), .B(new_n1105), .C1(new_n1032), .C2(G1956), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1098), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1071), .A2(new_n1085), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1084), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n626), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  AOI211_X1 g687(.A(new_n631), .B(new_n1084), .C1(new_n1071), .C2(new_n1085), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT60), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1105), .B1(new_n1032), .B2(G1956), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1101), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1117), .A2(KEYINPUT61), .A3(new_n1107), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1097), .A2(new_n1109), .A3(new_n1114), .A4(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1106), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1122));
  OR2_X1    g697(.A1(KEYINPUT124), .A2(G2078), .ZN(new_n1123));
  NAND2_X1  g698(.A1(KEYINPUT124), .A2(G2078), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1075), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT123), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1126), .B1(G160), .B2(G40), .ZN(new_n1127));
  NOR4_X1   g702(.A1(new_n476), .A2(new_n488), .A3(KEYINPUT123), .A4(new_n998), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1125), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n997), .A2(new_n1000), .ZN(new_n1130));
  OR2_X1    g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1131), .A2(G301), .A3(new_n1076), .A4(new_n1073), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1122), .B1(new_n1078), .B2(new_n1132), .ZN(new_n1133));
  OAI22_X1  g708(.A1(G1961), .A2(new_n1032), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1135));
  OAI21_X1  g710(.A(G171), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g713(.A(KEYINPUT125), .B(G171), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1077), .A2(G171), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1133), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1039), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1082), .A2(new_n1121), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1054), .A2(new_n1056), .A3(new_n830), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(G1981), .B2(G305), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1148), .A2(new_n1045), .B1(new_n1064), .B2(new_n1037), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1003), .A2(new_n1032), .B1(new_n1001), .B2(new_n737), .ZN(new_n1150));
  NAND2_X1  g725(.A1(G168), .A2(G8), .ZN(new_n1151));
  OAI21_X1  g726(.A(KEYINPUT118), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1002), .A2(new_n1007), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT118), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1153), .A2(new_n1154), .A3(G8), .A4(G168), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1039), .A2(new_n1064), .A3(new_n1065), .A4(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT63), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1037), .A2(new_n1158), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1064), .A2(new_n1160), .A3(new_n1036), .A4(new_n1156), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1081), .A2(new_n1146), .A3(new_n1149), .A4(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n997), .A2(new_n1029), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1087), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1165), .A2(new_n747), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1166), .B(KEYINPUT112), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n797), .B(G2067), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n748), .A2(new_n1087), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1164), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(KEYINPUT113), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT113), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1167), .A2(new_n1173), .A3(new_n1170), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n806), .B(new_n811), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1164), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1172), .A2(new_n1174), .A3(new_n1178), .ZN(new_n1179));
  OR2_X1    g754(.A1(G290), .A2(G1986), .ZN(new_n1180));
  NAND2_X1  g755(.A1(G290), .A2(G1986), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1176), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1163), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1164), .B1(new_n1168), .B2(new_n747), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1164), .A2(KEYINPUT46), .A3(new_n1087), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT46), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1165), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1185), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT47), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1180), .A2(new_n1176), .ZN(new_n1191));
  XOR2_X1   g766(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1192));
  XNOR2_X1  g767(.A(new_n1191), .B(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1190), .B1(new_n1179), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n806), .A2(new_n810), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1196), .B(KEYINPUT126), .ZN(new_n1197));
  OAI22_X1  g772(.A1(new_n1195), .A2(new_n1197), .B1(G2067), .B2(new_n797), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1194), .B1(new_n1198), .B2(new_n1164), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1184), .A2(new_n1199), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g775(.A1(G401), .A2(G227), .A3(new_n465), .ZN(new_n1202));
  AOI21_X1  g776(.A(new_n1202), .B1(new_n713), .B2(new_n716), .ZN(new_n1203));
  AND4_X1   g777(.A1(new_n905), .A2(new_n970), .A3(new_n1203), .A4(new_n977), .ZN(G308));
  NAND4_X1  g778(.A1(new_n970), .A2(new_n1203), .A3(new_n905), .A4(new_n977), .ZN(G225));
endmodule


