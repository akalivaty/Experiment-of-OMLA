//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT81), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G122), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT8), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G104), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n192), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G101), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(G104), .A3(new_n191), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G107), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n195), .A2(new_n196), .A3(new_n198), .A4(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n192), .A2(new_n200), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G101), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(KEYINPUT83), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT84), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G113), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT2), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT2), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G113), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(G116), .B(G119), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT67), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n211), .A2(new_n212), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n212), .A2(KEYINPUT5), .ZN(new_n217));
  INV_X1    g031(.A(G116), .ZN(new_n218));
  NOR3_X1   g032(.A1(new_n218), .A2(KEYINPUT5), .A3(G119), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(new_n207), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n214), .A2(new_n216), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n201), .A2(new_n203), .ZN(new_n222));
  OAI22_X1  g036(.A1(new_n206), .A2(new_n221), .B1(new_n205), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n217), .A2(new_n220), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n211), .A2(new_n212), .A3(new_n215), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n215), .B1(new_n211), .B2(new_n212), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n227), .B1(new_n205), .B2(new_n204), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n190), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G224), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(G953), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT7), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n234));
  INV_X1    g048(.A(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G143), .ZN(new_n236));
  INV_X1    g050(.A(G143), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G146), .ZN(new_n238));
  AOI21_X1  g052(.A(G128), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(KEYINPUT1), .A3(G146), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n234), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(G143), .B(G146), .ZN(new_n243));
  OAI211_X1 g057(.A(KEYINPUT66), .B(new_n240), .C1(new_n243), .C2(G128), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G125), .ZN(new_n246));
  INV_X1    g060(.A(G128), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(KEYINPUT1), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(new_n236), .A3(new_n238), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n245), .A2(KEYINPUT85), .A3(new_n246), .A4(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT0), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n243), .B1(new_n251), .B2(new_n247), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n247), .A3(KEYINPUT64), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT64), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n254), .B1(KEYINPUT0), .B2(G128), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n253), .A2(new_n255), .B1(KEYINPUT0), .B2(G128), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n252), .B1(new_n256), .B2(new_n243), .ZN(new_n257));
  OR2_X1    g071(.A1(new_n257), .A2(new_n246), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n250), .A2(new_n258), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n242), .A2(new_n244), .B1(new_n243), .B2(new_n248), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT85), .B1(new_n260), .B2(new_n246), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n233), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  OR2_X1    g076(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n263), .A2(new_n197), .B1(G104), .B2(new_n191), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n198), .A2(new_n200), .ZN(new_n265));
  OAI21_X1  g079(.A(G101), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT4), .A3(new_n201), .ZN(new_n267));
  INV_X1    g081(.A(new_n211), .ZN(new_n268));
  INV_X1    g082(.A(new_n212), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n225), .B2(new_n226), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT4), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n272), .B(G101), .C1(new_n264), .C2(new_n265), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n267), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n222), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n221), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n274), .A2(new_n276), .A3(new_n189), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n260), .A2(new_n246), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n278), .A2(new_n258), .A3(KEYINPUT7), .A4(new_n232), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n229), .A2(new_n262), .A3(new_n277), .A4(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G902), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n274), .A2(new_n276), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT82), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT6), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n274), .A2(new_n276), .A3(KEYINPUT82), .ZN(new_n287));
  INV_X1    g101(.A(new_n189), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n285), .A2(new_n286), .A3(new_n287), .A4(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n278), .A2(new_n258), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n290), .B(new_n231), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n274), .A2(new_n276), .A3(KEYINPUT82), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT82), .B1(new_n274), .B2(new_n276), .ZN(new_n293));
  NOR3_X1   g107(.A1(new_n292), .A2(new_n293), .A3(new_n189), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n277), .A2(KEYINPUT6), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n289), .B(new_n291), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(G210), .B1(G237), .B2(G902), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n282), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n297), .B1(new_n282), .B2(new_n296), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n188), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT86), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n282), .A2(new_n296), .ZN(new_n302));
  INV_X1    g116(.A(new_n297), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n282), .A2(new_n296), .A3(new_n297), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT86), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n307), .A3(new_n188), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n301), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G953), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G227), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n311), .B(KEYINPUT75), .ZN(new_n312));
  XNOR2_X1  g126(.A(G110), .B(G140), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n312), .B(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n249), .B(new_n240), .C1(G128), .C2(new_n243), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n201), .A3(new_n203), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n315), .A2(new_n201), .A3(KEYINPUT77), .A4(new_n203), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n257), .A2(new_n273), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n245), .A2(new_n249), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n201), .A2(KEYINPUT10), .A3(new_n203), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n267), .A2(new_n323), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT11), .ZN(new_n328));
  INV_X1    g142(.A(G134), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n328), .B1(new_n329), .B2(G137), .ZN(new_n330));
  INV_X1    g144(.A(G137), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT11), .A3(G134), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n329), .A2(G137), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G131), .ZN(new_n335));
  INV_X1    g149(.A(G131), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n330), .A2(new_n332), .A3(new_n336), .A4(new_n333), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(KEYINPUT79), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n322), .A2(new_n327), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT80), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT12), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n260), .A2(new_n222), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n320), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n344), .B1(new_n346), .B2(new_n338), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n318), .A2(new_n319), .B1(new_n260), .B2(new_n222), .ZN(new_n348));
  INV_X1    g162(.A(new_n338), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n348), .A2(new_n349), .A3(new_n343), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n314), .B(new_n341), .C1(new_n347), .C2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n321), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(new_n318), .B2(new_n319), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n266), .A2(KEYINPUT4), .A3(new_n201), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n257), .A2(new_n273), .ZN(new_n355));
  OAI22_X1  g169(.A1(new_n354), .A2(new_n355), .B1(new_n260), .B2(new_n325), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n338), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n341), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n314), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n351), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G469), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(new_n281), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n353), .A2(new_n356), .A3(new_n339), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(new_n359), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n357), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n346), .A2(new_n338), .A3(new_n344), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n343), .B1(new_n348), .B2(new_n349), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n364), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n366), .B(G469), .C1(new_n314), .C2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n362), .A2(new_n281), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n363), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G221), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT9), .B(G234), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n374), .B1(new_n376), .B2(new_n281), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G113), .B(G122), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(new_n199), .ZN(new_n381));
  XNOR2_X1  g195(.A(G125), .B(G140), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n382), .A2(new_n235), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n235), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n383), .A2(KEYINPUT87), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n383), .B1(KEYINPUT87), .B2(new_n384), .ZN(new_n386));
  INV_X1    g200(.A(G237), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n310), .A3(G214), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n237), .ZN(new_n389));
  NOR2_X1   g203(.A1(G237), .A2(G953), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(G143), .A3(G214), .ZN(new_n391));
  AOI22_X1  g205(.A1(new_n389), .A2(new_n391), .B1(KEYINPUT18), .B2(G131), .ZN(new_n392));
  AND4_X1   g206(.A1(KEYINPUT18), .A2(new_n389), .A3(G131), .A4(new_n391), .ZN(new_n393));
  OAI22_X1  g207(.A1(new_n385), .A2(new_n386), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n390), .A2(G143), .A3(G214), .ZN(new_n395));
  AOI21_X1  g209(.A(G143), .B1(new_n390), .B2(G214), .ZN(new_n396));
  OAI21_X1  g210(.A(G131), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT17), .ZN(new_n398));
  OR2_X1    g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G140), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G125), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n246), .A2(G140), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n402), .A3(KEYINPUT16), .ZN(new_n403));
  OR3_X1    g217(.A1(new_n246), .A2(KEYINPUT16), .A3(G140), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(new_n404), .A3(G146), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(G146), .B1(new_n403), .B2(new_n404), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT89), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n403), .A2(new_n404), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n235), .ZN(new_n411));
  AOI21_X1  g225(.A(KEYINPUT89), .B1(new_n411), .B2(new_n405), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n399), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n389), .A2(new_n336), .A3(new_n391), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n397), .A2(new_n398), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT90), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT90), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n397), .A2(new_n414), .A3(new_n417), .A4(new_n398), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n381), .B(new_n394), .C1(new_n413), .C2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n421));
  OR2_X1    g235(.A1(new_n382), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT19), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n382), .B1(KEYINPUT88), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n422), .A2(new_n235), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n397), .A2(new_n414), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n405), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n394), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n381), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n420), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n432));
  NOR2_X1   g246(.A1(G475), .A2(G902), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT91), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n420), .A2(new_n435), .A3(new_n430), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n435), .B1(new_n420), .B2(new_n430), .ZN(new_n437));
  INV_X1    g251(.A(new_n433), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n434), .B1(new_n439), .B2(new_n432), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n394), .B1(new_n413), .B2(new_n419), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n429), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n420), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n281), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G475), .ZN(new_n445));
  INV_X1    g259(.A(G122), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G116), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n218), .A2(G122), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT92), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n449), .B1(new_n447), .B2(new_n448), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n191), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n237), .A2(G128), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n247), .A2(G143), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G134), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n453), .A2(new_n454), .A3(new_n329), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n446), .A2(G116), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n191), .B1(new_n459), .B2(KEYINPUT14), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n447), .A2(new_n448), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n460), .B1(KEYINPUT14), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n452), .A2(new_n458), .A3(new_n462), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n450), .A2(new_n451), .A3(new_n191), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n218), .A2(G122), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT92), .B1(new_n465), .B2(new_n459), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n467));
  AOI21_X1  g281(.A(G107), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n457), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT13), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n470), .B1(new_n247), .B2(G143), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n237), .A2(KEYINPUT13), .A3(G128), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n454), .A3(new_n472), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n473), .A2(KEYINPUT93), .A3(G134), .ZN(new_n474));
  AOI21_X1  g288(.A(KEYINPUT93), .B1(new_n473), .B2(G134), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n463), .B1(new_n469), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT70), .B(G217), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n478), .A2(new_n375), .A3(G953), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n466), .A2(G107), .A3(new_n467), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n452), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n483), .B(new_n457), .C1(new_n475), .C2(new_n474), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n479), .B1(new_n484), .B2(new_n463), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n281), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G478), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(KEYINPUT15), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n477), .A2(new_n480), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n484), .A2(new_n463), .A3(new_n479), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n488), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n281), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n310), .A2(G952), .ZN(new_n496));
  INV_X1    g310(.A(G234), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n496), .B1(new_n497), .B2(new_n387), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT21), .B(G898), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(KEYINPUT95), .ZN(new_n501));
  OAI211_X1 g315(.A(G902), .B(G953), .C1(new_n497), .C2(new_n387), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(KEYINPUT94), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n495), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n440), .A2(new_n445), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n379), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n309), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT32), .ZN(new_n509));
  XOR2_X1   g323(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n510));
  NAND2_X1  g324(.A1(new_n390), .A2(G210), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT26), .B(G101), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n271), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n338), .A2(new_n257), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n329), .A2(G137), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n331), .A2(G134), .ZN(new_n518));
  OAI21_X1  g332(.A(G131), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n337), .A2(new_n519), .A3(KEYINPUT68), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT68), .B1(new_n337), .B2(new_n519), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n515), .B(new_n516), .C1(new_n522), .C2(new_n260), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT28), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n337), .A2(new_n519), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT68), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n337), .A2(new_n519), .A3(KEYINPUT68), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n324), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT28), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n515), .A4(new_n516), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n524), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT65), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n337), .A2(new_n519), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n534), .B1(new_n337), .B2(new_n519), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n260), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n516), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n271), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n514), .B1(new_n533), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT31), .ZN(new_n542));
  INV_X1    g356(.A(new_n537), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n324), .A2(new_n535), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT30), .B1(new_n544), .B2(new_n516), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n249), .A2(new_n245), .B1(new_n527), .B2(new_n528), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n516), .A2(KEYINPUT30), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n271), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n523), .A2(new_n514), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n542), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT30), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(new_n538), .B2(new_n539), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n552), .B1(new_n338), .B2(new_n257), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n515), .B1(new_n530), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n550), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT31), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n541), .B1(new_n551), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(G472), .A2(G902), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n509), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n533), .A2(new_n540), .ZN(new_n563));
  INV_X1    g377(.A(new_n514), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n549), .A2(new_n542), .A3(new_n550), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT31), .B1(new_n556), .B2(new_n557), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n568), .A2(KEYINPUT32), .A3(new_n560), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n515), .B1(new_n530), .B2(new_n516), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n570), .B1(new_n524), .B2(new_n532), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT29), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n564), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(G902), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n523), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(new_n553), .B2(new_n555), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n572), .B1(new_n576), .B2(new_n514), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n533), .A2(new_n540), .A3(new_n514), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n574), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G472), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n562), .A2(new_n569), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT25), .ZN(new_n582));
  INV_X1    g396(.A(G119), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G128), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n247), .A2(G119), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT24), .B(G110), .ZN(new_n587));
  OR2_X1    g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n247), .A2(KEYINPUT23), .A3(G119), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n583), .A2(G128), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n589), .B(new_n584), .C1(new_n590), .C2(KEYINPUT23), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n591), .A2(KEYINPUT71), .A3(G110), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT71), .B1(new_n591), .B2(G110), .ZN(new_n593));
  OAI221_X1 g407(.A(new_n588), .B1(new_n406), .B2(new_n407), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n586), .A2(new_n587), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT73), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT72), .B(G110), .Z(new_n598));
  INV_X1    g412(.A(KEYINPUT23), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n585), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n598), .A2(new_n589), .A3(new_n584), .A4(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT73), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n597), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n405), .A2(new_n384), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n594), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT22), .B(G137), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n374), .A2(new_n497), .A3(G953), .ZN(new_n608));
  XOR2_X1   g422(.A(new_n607), .B(new_n608), .Z(new_n609));
  NAND2_X1  g423(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n606), .A2(KEYINPUT74), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT74), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n592), .A2(new_n593), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n588), .B1(new_n406), .B2(new_n407), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n605), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n609), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n611), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n582), .B1(new_n619), .B2(G902), .ZN(new_n620));
  INV_X1    g434(.A(new_n616), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n613), .B1(new_n594), .B2(new_n605), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n618), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n610), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n624), .A2(KEYINPUT25), .A3(new_n281), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n478), .B1(G234), .B2(new_n281), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(G902), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n626), .A2(new_n627), .B1(new_n624), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n581), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n508), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G101), .ZN(G3));
  OAI21_X1  g446(.A(G472), .B1(new_n559), .B2(G902), .ZN(new_n633));
  AOI21_X1  g447(.A(KEYINPUT25), .B1(new_n624), .B2(new_n281), .ZN(new_n634));
  AOI211_X1 g448(.A(new_n582), .B(G902), .C1(new_n623), .C2(new_n610), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n627), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n568), .A2(new_n560), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n624), .A2(new_n628), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n633), .A2(new_n636), .A3(new_n637), .A4(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(KEYINPUT96), .B1(new_n379), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(G902), .B1(new_n351), .B2(new_n360), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n371), .B1(new_n641), .B2(new_n362), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n377), .B1(new_n642), .B2(new_n370), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n633), .A2(new_n637), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT96), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n643), .A2(new_n644), .A3(new_n645), .A4(new_n629), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n504), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n187), .B(new_n649), .C1(new_n298), .C2(new_n299), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT97), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT33), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n492), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n490), .B(new_n491), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n653), .A2(G478), .A3(new_n281), .A4(new_n656), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n487), .A2(KEYINPUT98), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n487), .A2(KEYINPUT98), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n486), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n434), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n431), .A2(KEYINPUT91), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n420), .A2(new_n435), .A3(new_n430), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n663), .A2(new_n433), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n662), .B1(new_n665), .B2(KEYINPUT20), .ZN(new_n666));
  INV_X1    g480(.A(new_n445), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n661), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n650), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n648), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT34), .B(G104), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G6));
  NOR2_X1   g486(.A1(new_n436), .A2(new_n437), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n432), .B1(new_n673), .B2(new_n433), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n663), .A2(new_n432), .A3(new_n433), .A4(new_n664), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n445), .B(new_n495), .C1(new_n674), .C2(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n650), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n648), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT35), .B(G107), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G9));
  NOR2_X1   g495(.A1(new_n618), .A2(KEYINPUT36), .ZN(new_n682));
  XOR2_X1   g496(.A(new_n617), .B(new_n682), .Z(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n628), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n636), .A2(new_n684), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n685), .A2(new_n637), .A3(new_n633), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n508), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT37), .B(G110), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT99), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n687), .B(new_n689), .ZN(G12));
  INV_X1    g504(.A(new_n187), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(new_n304), .B2(new_n305), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n581), .A2(new_n692), .A3(new_n685), .ZN(new_n693));
  INV_X1    g507(.A(G900), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n499), .B1(new_n503), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n373), .A2(new_n378), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n677), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n693), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G128), .ZN(G30));
  XNOR2_X1  g514(.A(new_n695), .B(KEYINPUT39), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n379), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT101), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT40), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n702), .B(KEYINPUT101), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT40), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n306), .B(KEYINPUT38), .Z(new_n709));
  INV_X1    g523(.A(new_n570), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n514), .B1(new_n710), .B2(new_n523), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n711), .A2(KEYINPUT100), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n556), .A2(new_n557), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n713), .B1(new_n711), .B2(KEYINPUT100), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n281), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(G472), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n562), .A3(new_n569), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n626), .A2(new_n627), .B1(new_n628), .B2(new_n683), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(new_n187), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n495), .B1(new_n666), .B2(new_n667), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n709), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n706), .A2(new_n708), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G143), .ZN(G45));
  OAI211_X1 g537(.A(new_n661), .B(new_n696), .C1(new_n666), .C2(new_n667), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n379), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n693), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G146), .ZN(G48));
  NAND2_X1  g541(.A1(new_n367), .A2(new_n368), .ZN(new_n728));
  AOI22_X1  g542(.A1(new_n365), .A2(new_n728), .B1(new_n358), .B2(new_n359), .ZN(new_n729));
  OAI21_X1  g543(.A(G469), .B1(new_n729), .B2(G902), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n363), .A3(new_n378), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n630), .A2(new_n669), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT41), .B(G113), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G15));
  NAND4_X1  g549(.A1(new_n678), .A2(new_n581), .A3(new_n629), .A4(new_n732), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G116), .ZN(G18));
  OAI21_X1  g551(.A(new_n187), .B1(new_n298), .B2(new_n299), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n731), .ZN(new_n739));
  INV_X1    g553(.A(new_n506), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n739), .A2(new_n581), .A3(new_n740), .A4(new_n685), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G119), .ZN(G21));
  NOR2_X1   g556(.A1(new_n738), .A2(new_n720), .ZN(new_n743));
  OAI22_X1  g557(.A1(new_n566), .A2(new_n567), .B1(new_n514), .B2(new_n571), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n560), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n633), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n636), .A2(new_n638), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n730), .A2(new_n363), .A3(new_n378), .A4(new_n649), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n743), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G122), .ZN(G24));
  NOR2_X1   g566(.A1(new_n718), .A2(new_n746), .ZN(new_n753));
  INV_X1    g567(.A(new_n724), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(new_n739), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G125), .ZN(G27));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n754), .A2(new_n643), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n298), .A2(new_n299), .A3(new_n691), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n581), .A2(new_n629), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n757), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n304), .A2(new_n305), .A3(new_n187), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n379), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n562), .A2(KEYINPUT102), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT102), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n637), .A2(new_n765), .A3(new_n509), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n764), .A2(new_n766), .A3(new_n569), .A4(new_n580), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n724), .A2(new_n757), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n763), .A2(new_n767), .A3(new_n629), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n761), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G131), .ZN(G33));
  AND3_X1   g585(.A1(new_n581), .A2(new_n629), .A3(new_n759), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n698), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G134), .ZN(G36));
  NOR2_X1   g588(.A1(new_n666), .A2(new_n667), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n661), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT43), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n644), .A2(new_n718), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(KEYINPUT44), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT104), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT44), .B1(new_n778), .B2(new_n779), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n762), .B1(new_n782), .B2(KEYINPUT105), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n366), .B1(new_n314), .B2(new_n369), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT45), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n362), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n786), .B1(new_n785), .B2(new_n784), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(KEYINPUT46), .A3(new_n372), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT46), .B1(new_n787), .B2(new_n372), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT103), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n363), .B(new_n788), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n378), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n701), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n782), .A2(KEYINPUT105), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n781), .A2(new_n783), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G137), .ZN(G39));
  INV_X1    g611(.A(KEYINPUT47), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(KEYINPUT47), .B(new_n378), .C1(new_n791), .C2(new_n792), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n759), .A2(new_n747), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n802), .A2(new_n581), .A3(new_n724), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT106), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT106), .ZN(new_n805));
  INV_X1    g619(.A(new_n803), .ZN(new_n806));
  AOI211_X1 g620(.A(new_n805), .B(new_n806), .C1(new_n799), .C2(new_n800), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  XOR2_X1   g622(.A(KEYINPUT107), .B(G140), .Z(new_n809));
  XNOR2_X1  g623(.A(new_n808), .B(new_n809), .ZN(G42));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n811));
  INV_X1    g625(.A(new_n717), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n762), .A2(new_n731), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n812), .A2(new_n629), .A3(new_n813), .A4(new_n499), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n440), .A2(new_n445), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n814), .A2(new_n815), .A3(new_n661), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n778), .A2(new_n499), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n748), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n732), .A2(KEYINPUT111), .A3(new_n691), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT111), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n821), .B1(new_n731), .B2(new_n187), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n709), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  OR3_X1    g637(.A1(new_n818), .A2(new_n819), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n819), .B1(new_n818), .B2(new_n823), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n816), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT112), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n817), .A2(new_n827), .A3(new_n813), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n827), .B1(new_n817), .B2(new_n813), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n753), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n801), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n730), .A2(new_n363), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n377), .ZN(new_n834));
  AOI211_X1 g648(.A(new_n762), .B(new_n818), .C1(new_n832), .C2(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n811), .B1(new_n831), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n739), .ZN(new_n837));
  OAI221_X1 g651(.A(new_n496), .B1(new_n668), .B2(new_n814), .C1(new_n818), .C2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n765), .B1(new_n637), .B2(new_n509), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n569), .A2(new_n580), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n747), .B1(new_n841), .B2(new_n766), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n828), .B2(new_n829), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n843), .A2(KEYINPUT48), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(KEYINPUT48), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n838), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n832), .A2(KEYINPUT113), .A3(new_n834), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n847), .A2(new_n748), .A3(new_n759), .A4(new_n817), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT113), .B1(new_n832), .B2(new_n834), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n826), .A2(KEYINPUT51), .A3(new_n830), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n836), .B(new_n846), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n665), .A2(KEYINPUT20), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n675), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT108), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n493), .B1(new_n492), .B2(new_n281), .ZN(new_n856));
  AOI211_X1 g670(.A(G902), .B(new_n488), .C1(new_n490), .C2(new_n491), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n489), .A2(KEYINPUT108), .A3(new_n494), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n695), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n854), .A2(new_n445), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT109), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n854), .A2(new_n860), .A3(KEYINPUT109), .A4(new_n445), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n863), .A2(new_n581), .A3(new_n685), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n753), .A2(new_n754), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n763), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n504), .B1(new_n301), .B2(new_n308), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n858), .A2(new_n859), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n668), .B1(new_n815), .B2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n869), .A2(new_n640), .A3(new_n646), .A4(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n309), .B(new_n507), .C1(new_n630), .C2(new_n686), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n868), .A2(new_n773), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n749), .A2(new_n746), .A3(new_n747), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n738), .A2(new_n506), .A3(new_n731), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n581), .A2(new_n685), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n743), .A2(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n770), .A2(new_n733), .A3(new_n736), .A4(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n685), .A2(new_n695), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n743), .A2(new_n881), .A3(new_n643), .A4(new_n717), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n699), .A2(new_n726), .A3(new_n755), .A4(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT52), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n693), .B1(new_n698), .B2(new_n725), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n886), .A2(KEYINPUT52), .A3(new_n755), .A4(new_n882), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT53), .B1(new_n880), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n772), .A2(new_n725), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n759), .A2(new_n378), .A3(new_n373), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n815), .A2(KEYINPUT42), .A3(new_n661), .A4(new_n696), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI22_X1  g707(.A1(new_n890), .A2(new_n757), .B1(new_n842), .B2(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n733), .A2(new_n736), .A3(new_n741), .A4(new_n751), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT53), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n872), .A2(new_n873), .A3(new_n773), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n891), .B1(new_n865), .B2(new_n866), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n888), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT110), .ZN(new_n902));
  AND4_X1   g716(.A1(new_n733), .A2(new_n736), .A3(new_n741), .A4(new_n751), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(KEYINPUT53), .A3(new_n770), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n904), .A2(new_n874), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT110), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n905), .A2(new_n906), .A3(new_n888), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n889), .B1(new_n902), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT54), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n900), .A2(new_n770), .A3(new_n903), .ZN(new_n911));
  INV_X1    g725(.A(new_n888), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n896), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n901), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT54), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  OAI22_X1  g730(.A1(new_n852), .A2(new_n916), .B1(G952), .B2(G953), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT49), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n833), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n629), .A2(new_n188), .A3(new_n378), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n833), .A2(new_n918), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n776), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n922), .A2(new_n812), .A3(new_n709), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n917), .A2(new_n924), .ZN(G75));
  NOR2_X1   g739(.A1(new_n310), .A2(G952), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(G210), .A2(G902), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n908), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n289), .B1(new_n294), .B2(new_n295), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(new_n291), .ZN(new_n931));
  XNOR2_X1  g745(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n933), .A2(KEYINPUT56), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n927), .B1(new_n929), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT115), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n908), .B2(new_n928), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n906), .B1(new_n905), .B2(new_n888), .ZN(new_n938));
  AND4_X1   g752(.A1(new_n906), .A2(new_n888), .A3(new_n897), .A4(new_n900), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n913), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n928), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n940), .A2(KEYINPUT115), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT56), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n937), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n933), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(KEYINPUT116), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT116), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n944), .A2(new_n947), .A3(new_n933), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n935), .B1(new_n946), .B2(new_n948), .ZN(G51));
  NAND2_X1  g763(.A1(new_n940), .A2(KEYINPUT54), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT117), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n950), .A2(new_n910), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n940), .A2(KEYINPUT117), .A3(KEYINPUT54), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n371), .B(KEYINPUT57), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n361), .ZN(new_n956));
  OR3_X1    g770(.A1(new_n908), .A2(new_n281), .A3(new_n787), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n926), .B1(new_n956), .B2(new_n957), .ZN(G54));
  INV_X1    g772(.A(KEYINPUT118), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n908), .A2(new_n281), .ZN(new_n960));
  AND2_X1   g774(.A1(KEYINPUT58), .A2(G475), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n673), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n926), .B1(new_n962), .B2(new_n963), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n960), .A2(KEYINPUT118), .A3(new_n673), .A4(new_n961), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(G60));
  XNOR2_X1  g781(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n487), .A2(new_n281), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n968), .B(new_n969), .Z(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n910), .B2(new_n915), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n653), .A2(new_n656), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n927), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n952), .A2(new_n953), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n973), .A2(new_n970), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(G63));
  NAND2_X1  g791(.A1(G217), .A2(G902), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT60), .Z(new_n979));
  XNOR2_X1  g793(.A(new_n683), .B(KEYINPUT120), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n940), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n940), .A2(new_n979), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n927), .B(new_n981), .C1(new_n982), .C2(new_n624), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT61), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n983), .B(new_n984), .ZN(G66));
  OAI21_X1  g799(.A(G953), .B1(new_n501), .B2(new_n230), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n903), .A2(new_n872), .A3(new_n873), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n986), .B1(new_n988), .B2(G953), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n930), .B1(G898), .B2(new_n310), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(G69));
  AOI21_X1  g805(.A(new_n545), .B1(new_n530), .B2(new_n554), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT121), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n422), .A2(new_n424), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n993), .B(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n995), .B1(G900), .B2(G953), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n794), .A2(new_n743), .A3(new_n842), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n886), .A2(new_n755), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT123), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n796), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n770), .A2(new_n773), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT124), .Z(new_n1004));
  NOR3_X1   g818(.A1(new_n808), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n997), .B1(new_n1005), .B2(new_n310), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n310), .B1(G227), .B2(G900), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n722), .A2(new_n1001), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(KEYINPUT62), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n704), .A2(new_n772), .A3(new_n871), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n1011), .A2(new_n796), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n808), .ZN(new_n1014));
  OR2_X1    g828(.A1(new_n1010), .A2(KEYINPUT62), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  AND2_X1   g830(.A1(new_n1016), .A2(new_n310), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n995), .B(KEYINPUT122), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n1007), .B(new_n1009), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1018), .B1(new_n1016), .B2(new_n310), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1008), .B1(new_n1020), .B2(new_n1006), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1019), .A2(new_n1021), .ZN(G72));
  XNOR2_X1  g836(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1023));
  NAND2_X1  g837(.A1(G472), .A2(G902), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n576), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(new_n564), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1025), .B1(new_n1027), .B2(new_n713), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n926), .B1(new_n914), .B2(new_n1028), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1025), .B(KEYINPUT126), .Z(new_n1030));
  AOI21_X1  g844(.A(new_n1030), .B1(new_n1005), .B2(new_n988), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n576), .A2(new_n564), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g847(.A1(new_n1013), .A2(new_n1014), .A3(new_n988), .A4(new_n1015), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1030), .ZN(new_n1035));
  AOI21_X1  g849(.A(KEYINPUT127), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1026), .A2(new_n514), .ZN(new_n1037));
  NOR2_X1   g851(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1034), .A2(KEYINPUT127), .A3(new_n1035), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1033), .B1(new_n1038), .B2(new_n1039), .ZN(G57));
endmodule


