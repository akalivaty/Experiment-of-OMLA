

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U555 ( .A(n538), .B(KEYINPUT67), .ZN(n982) );
  XNOR2_X2 U556 ( .A(n558), .B(n557), .ZN(G160) );
  OR2_X1 U557 ( .A1(n715), .A2(n714), .ZN(n719) );
  OR2_X1 U558 ( .A1(n811), .A2(n810), .ZN(n826) );
  AND2_X1 U559 ( .A1(n912), .A2(n823), .ZN(n522) );
  NOR2_X1 U560 ( .A1(n708), .A2(n707), .ZN(n712) );
  NAND2_X1 U561 ( .A1(n697), .A2(n779), .ZN(n702) );
  XNOR2_X1 U562 ( .A(n588), .B(n587), .ZN(n589) );
  OR2_X1 U563 ( .A1(n809), .A2(n522), .ZN(n810) );
  NOR2_X1 U564 ( .A1(G543), .A2(n528), .ZN(n529) );
  NOR2_X2 U565 ( .A1(G2105), .A2(n541), .ZN(n987) );
  NAND2_X1 U566 ( .A1(n597), .A2(n596), .ZN(n1015) );
  NAND2_X1 U567 ( .A1(n556), .A2(n555), .ZN(n558) );
  NOR2_X1 U568 ( .A1(G651), .A2(G543), .ZN(n660) );
  NAND2_X1 U569 ( .A1(G89), .A2(n660), .ZN(n523) );
  XNOR2_X1 U570 ( .A(n523), .B(KEYINPUT78), .ZN(n524) );
  XNOR2_X1 U571 ( .A(n524), .B(KEYINPUT4), .ZN(n526) );
  XOR2_X1 U572 ( .A(G543), .B(KEYINPUT0), .Z(n649) );
  INV_X1 U573 ( .A(G651), .ZN(n528) );
  NOR2_X1 U574 ( .A1(n649), .A2(n528), .ZN(n664) );
  NAND2_X1 U575 ( .A1(G76), .A2(n664), .ZN(n525) );
  NAND2_X1 U576 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U577 ( .A(n527), .B(KEYINPUT5), .ZN(n534) );
  XOR2_X1 U578 ( .A(KEYINPUT1), .B(n529), .Z(n659) );
  NAND2_X1 U579 ( .A1(G63), .A2(n659), .ZN(n531) );
  NOR2_X2 U580 ( .A1(G651), .A2(n649), .ZN(n663) );
  NAND2_X1 U581 ( .A1(G51), .A2(n663), .ZN(n530) );
  NAND2_X1 U582 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U583 ( .A(KEYINPUT6), .B(n532), .Z(n533) );
  NAND2_X1 U584 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U585 ( .A(n535), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U586 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U587 ( .A1(G2104), .A2(G2105), .ZN(n536) );
  XOR2_X2 U588 ( .A(KEYINPUT17), .B(n536), .Z(n986) );
  NAND2_X1 U589 ( .A1(n986), .A2(G138), .ZN(n537) );
  XNOR2_X1 U590 ( .A(n537), .B(KEYINPUT92), .ZN(n540) );
  INV_X1 U591 ( .A(G2104), .ZN(n542) );
  NAND2_X1 U592 ( .A1(G2105), .A2(G2104), .ZN(n538) );
  NAND2_X1 U593 ( .A1(G114), .A2(n982), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n540), .A2(n539), .ZN(n547) );
  INV_X1 U595 ( .A(G2104), .ZN(n541) );
  NAND2_X1 U596 ( .A1(G102), .A2(n987), .ZN(n545) );
  NAND2_X1 U597 ( .A1(n542), .A2(G2105), .ZN(n543) );
  XNOR2_X1 U598 ( .A(n543), .B(KEYINPUT65), .ZN(n983) );
  NAND2_X1 U599 ( .A1(G126), .A2(n983), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X2 U601 ( .A1(n547), .A2(n546), .ZN(G164) );
  INV_X1 U602 ( .A(KEYINPUT23), .ZN(n549) );
  NAND2_X1 U603 ( .A1(G101), .A2(n987), .ZN(n548) );
  XNOR2_X1 U604 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U605 ( .A(n550), .B(KEYINPUT66), .ZN(n556) );
  AND2_X1 U606 ( .A1(G125), .A2(n983), .ZN(n554) );
  NAND2_X1 U607 ( .A1(G137), .A2(n986), .ZN(n552) );
  NAND2_X1 U608 ( .A1(G113), .A2(n982), .ZN(n551) );
  NAND2_X1 U609 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U610 ( .A1(n554), .A2(n553), .ZN(n555) );
  INV_X1 U611 ( .A(KEYINPUT64), .ZN(n557) );
  XOR2_X1 U612 ( .A(G2443), .B(G2446), .Z(n560) );
  XNOR2_X1 U613 ( .A(G2427), .B(G2451), .ZN(n559) );
  XNOR2_X1 U614 ( .A(n560), .B(n559), .ZN(n566) );
  XOR2_X1 U615 ( .A(G2430), .B(G2454), .Z(n562) );
  XNOR2_X1 U616 ( .A(G1341), .B(G1348), .ZN(n561) );
  XNOR2_X1 U617 ( .A(n562), .B(n561), .ZN(n564) );
  XOR2_X1 U618 ( .A(G2435), .B(G2438), .Z(n563) );
  XNOR2_X1 U619 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U620 ( .A(n566), .B(n565), .Z(n567) );
  AND2_X1 U621 ( .A1(G14), .A2(n567), .ZN(G401) );
  NAND2_X1 U622 ( .A1(n663), .A2(G52), .ZN(n568) );
  XNOR2_X1 U623 ( .A(KEYINPUT69), .B(n568), .ZN(n576) );
  NAND2_X1 U624 ( .A1(G90), .A2(n660), .ZN(n570) );
  NAND2_X1 U625 ( .A1(G77), .A2(n664), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U627 ( .A(n571), .B(KEYINPUT70), .ZN(n572) );
  XNOR2_X1 U628 ( .A(n572), .B(KEYINPUT9), .ZN(n574) );
  NAND2_X1 U629 ( .A1(n659), .A2(G64), .ZN(n573) );
  NAND2_X1 U630 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U631 ( .A1(n576), .A2(n575), .ZN(G171) );
  AND2_X1 U632 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U633 ( .A(G57), .ZN(G237) );
  INV_X1 U634 ( .A(G69), .ZN(G235) );
  INV_X1 U635 ( .A(G108), .ZN(G238) );
  INV_X1 U636 ( .A(G120), .ZN(G236) );
  INV_X1 U637 ( .A(G132), .ZN(G219) );
  INV_X1 U638 ( .A(G82), .ZN(G220) );
  NAND2_X1 U639 ( .A1(G88), .A2(n660), .ZN(n578) );
  NAND2_X1 U640 ( .A1(G75), .A2(n664), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n578), .A2(n577), .ZN(n583) );
  NAND2_X1 U642 ( .A1(G62), .A2(n659), .ZN(n579) );
  XOR2_X1 U643 ( .A(KEYINPUT87), .B(n579), .Z(n581) );
  NAND2_X1 U644 ( .A1(n663), .A2(G50), .ZN(n580) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U646 ( .A1(n583), .A2(n582), .ZN(G166) );
  XOR2_X1 U647 ( .A(KEYINPUT10), .B(KEYINPUT73), .Z(n585) );
  NAND2_X1 U648 ( .A1(G7), .A2(G661), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(G223) );
  INV_X1 U650 ( .A(G223), .ZN(n828) );
  NAND2_X1 U651 ( .A1(n828), .A2(G567), .ZN(n586) );
  XOR2_X1 U652 ( .A(KEYINPUT11), .B(n586), .Z(G234) );
  NAND2_X1 U653 ( .A1(G56), .A2(n659), .ZN(n588) );
  XOR2_X1 U654 ( .A(KEYINPUT14), .B(KEYINPUT75), .Z(n587) );
  XOR2_X1 U655 ( .A(KEYINPUT74), .B(n589), .Z(n595) );
  NAND2_X1 U656 ( .A1(n660), .A2(G81), .ZN(n590) );
  XNOR2_X1 U657 ( .A(n590), .B(KEYINPUT12), .ZN(n592) );
  NAND2_X1 U658 ( .A1(G68), .A2(n664), .ZN(n591) );
  NAND2_X1 U659 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U660 ( .A(KEYINPUT13), .B(n593), .Z(n594) );
  NOR2_X1 U661 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U662 ( .A1(n663), .A2(G43), .ZN(n596) );
  INV_X1 U663 ( .A(G860), .ZN(n955) );
  OR2_X1 U664 ( .A1(n1015), .A2(n955), .ZN(G153) );
  INV_X1 U665 ( .A(G171), .ZN(G301) );
  NAND2_X1 U666 ( .A1(G868), .A2(G301), .ZN(n608) );
  NAND2_X1 U667 ( .A1(G66), .A2(n659), .ZN(n599) );
  NAND2_X1 U668 ( .A1(G92), .A2(n660), .ZN(n598) );
  NAND2_X1 U669 ( .A1(n599), .A2(n598), .ZN(n605) );
  NAND2_X1 U670 ( .A1(n663), .A2(G54), .ZN(n600) );
  XNOR2_X1 U671 ( .A(n600), .B(KEYINPUT76), .ZN(n602) );
  NAND2_X1 U672 ( .A1(G79), .A2(n664), .ZN(n601) );
  NAND2_X1 U673 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U674 ( .A(KEYINPUT77), .B(n603), .Z(n604) );
  NOR2_X1 U675 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U676 ( .A(KEYINPUT15), .B(n606), .ZN(n710) );
  INV_X1 U677 ( .A(G868), .ZN(n677) );
  NAND2_X1 U678 ( .A1(n710), .A2(n677), .ZN(n607) );
  NAND2_X1 U679 ( .A1(n608), .A2(n607), .ZN(G284) );
  NAND2_X1 U680 ( .A1(n663), .A2(G53), .ZN(n609) );
  XOR2_X1 U681 ( .A(KEYINPUT71), .B(n609), .Z(n611) );
  NAND2_X1 U682 ( .A1(n659), .A2(G65), .ZN(n610) );
  NAND2_X1 U683 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U684 ( .A(KEYINPUT72), .B(n612), .Z(n616) );
  NAND2_X1 U685 ( .A1(G91), .A2(n660), .ZN(n614) );
  NAND2_X1 U686 ( .A1(G78), .A2(n664), .ZN(n613) );
  AND2_X1 U687 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n616), .A2(n615), .ZN(G299) );
  NOR2_X1 U689 ( .A1(G286), .A2(n677), .ZN(n617) );
  XOR2_X1 U690 ( .A(KEYINPUT79), .B(n617), .Z(n619) );
  NOR2_X1 U691 ( .A1(G868), .A2(G299), .ZN(n618) );
  NOR2_X1 U692 ( .A1(n619), .A2(n618), .ZN(G297) );
  NAND2_X1 U693 ( .A1(n955), .A2(G559), .ZN(n620) );
  INV_X1 U694 ( .A(n710), .ZN(n1012) );
  NAND2_X1 U695 ( .A1(n620), .A2(n1012), .ZN(n621) );
  XNOR2_X1 U696 ( .A(n621), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U697 ( .A1(n1012), .A2(G868), .ZN(n622) );
  NOR2_X1 U698 ( .A1(G559), .A2(n622), .ZN(n623) );
  XOR2_X1 U699 ( .A(KEYINPUT81), .B(n623), .Z(n626) );
  NOR2_X1 U700 ( .A1(G868), .A2(n1015), .ZN(n624) );
  XNOR2_X1 U701 ( .A(KEYINPUT80), .B(n624), .ZN(n625) );
  NOR2_X1 U702 ( .A1(n626), .A2(n625), .ZN(G282) );
  NAND2_X1 U703 ( .A1(G123), .A2(n983), .ZN(n627) );
  XNOR2_X1 U704 ( .A(n627), .B(KEYINPUT18), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G135), .A2(n986), .ZN(n628) );
  XNOR2_X1 U706 ( .A(n628), .B(KEYINPUT82), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U708 ( .A1(G111), .A2(n982), .ZN(n632) );
  NAND2_X1 U709 ( .A1(G99), .A2(n987), .ZN(n631) );
  NAND2_X1 U710 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U711 ( .A1(n634), .A2(n633), .ZN(n995) );
  XNOR2_X1 U712 ( .A(n995), .B(G2096), .ZN(n636) );
  INV_X1 U713 ( .A(G2100), .ZN(n635) );
  NAND2_X1 U714 ( .A1(n636), .A2(n635), .ZN(G156) );
  NAND2_X1 U715 ( .A1(n664), .A2(G73), .ZN(n638) );
  XNOR2_X1 U716 ( .A(KEYINPUT2), .B(KEYINPUT86), .ZN(n637) );
  XNOR2_X1 U717 ( .A(n638), .B(n637), .ZN(n645) );
  NAND2_X1 U718 ( .A1(G48), .A2(n663), .ZN(n640) );
  NAND2_X1 U719 ( .A1(G86), .A2(n660), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U721 ( .A1(G61), .A2(n659), .ZN(n641) );
  XNOR2_X1 U722 ( .A(KEYINPUT85), .B(n641), .ZN(n642) );
  NOR2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U724 ( .A1(n645), .A2(n644), .ZN(G305) );
  NAND2_X1 U725 ( .A1(G49), .A2(n663), .ZN(n647) );
  NAND2_X1 U726 ( .A1(G74), .A2(G651), .ZN(n646) );
  NAND2_X1 U727 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U728 ( .A1(n659), .A2(n648), .ZN(n651) );
  NAND2_X1 U729 ( .A1(n649), .A2(G87), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(G288) );
  NAND2_X1 U731 ( .A1(G60), .A2(n659), .ZN(n653) );
  NAND2_X1 U732 ( .A1(G47), .A2(n663), .ZN(n652) );
  NAND2_X1 U733 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U734 ( .A(KEYINPUT68), .B(n654), .Z(n658) );
  NAND2_X1 U735 ( .A1(G85), .A2(n660), .ZN(n656) );
  NAND2_X1 U736 ( .A1(G72), .A2(n664), .ZN(n655) );
  AND2_X1 U737 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U738 ( .A1(n658), .A2(n657), .ZN(G290) );
  NAND2_X1 U739 ( .A1(G67), .A2(n659), .ZN(n662) );
  NAND2_X1 U740 ( .A1(G93), .A2(n660), .ZN(n661) );
  NAND2_X1 U741 ( .A1(n662), .A2(n661), .ZN(n668) );
  NAND2_X1 U742 ( .A1(G55), .A2(n663), .ZN(n666) );
  NAND2_X1 U743 ( .A1(G80), .A2(n664), .ZN(n665) );
  NAND2_X1 U744 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U745 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U746 ( .A(KEYINPUT84), .B(n669), .Z(n954) );
  XNOR2_X1 U747 ( .A(KEYINPUT19), .B(G305), .ZN(n670) );
  XNOR2_X1 U748 ( .A(n670), .B(G288), .ZN(n671) );
  XNOR2_X1 U749 ( .A(n954), .B(n671), .ZN(n673) );
  XNOR2_X1 U750 ( .A(G290), .B(G166), .ZN(n672) );
  XNOR2_X1 U751 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U752 ( .A(n674), .B(G299), .ZN(n1013) );
  NAND2_X1 U753 ( .A1(G559), .A2(n1012), .ZN(n675) );
  XOR2_X1 U754 ( .A(n1015), .B(n675), .Z(n956) );
  XOR2_X1 U755 ( .A(n1013), .B(n956), .Z(n676) );
  NOR2_X1 U756 ( .A1(n677), .A2(n676), .ZN(n679) );
  NOR2_X1 U757 ( .A1(n954), .A2(G868), .ZN(n678) );
  NOR2_X1 U758 ( .A1(n679), .A2(n678), .ZN(G295) );
  NAND2_X1 U759 ( .A1(G2078), .A2(G2084), .ZN(n681) );
  XOR2_X1 U760 ( .A(KEYINPUT20), .B(KEYINPUT88), .Z(n680) );
  XNOR2_X1 U761 ( .A(n681), .B(n680), .ZN(n682) );
  NAND2_X1 U762 ( .A1(G2090), .A2(n682), .ZN(n683) );
  XNOR2_X1 U763 ( .A(KEYINPUT21), .B(n683), .ZN(n684) );
  NAND2_X1 U764 ( .A1(n684), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U765 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U766 ( .A1(G220), .A2(G219), .ZN(n685) );
  XOR2_X1 U767 ( .A(KEYINPUT22), .B(n685), .Z(n686) );
  NOR2_X1 U768 ( .A1(G218), .A2(n686), .ZN(n687) );
  XOR2_X1 U769 ( .A(KEYINPUT89), .B(n687), .Z(n688) );
  NAND2_X1 U770 ( .A1(G96), .A2(n688), .ZN(n959) );
  NAND2_X1 U771 ( .A1(G2106), .A2(n959), .ZN(n693) );
  NOR2_X1 U772 ( .A1(G236), .A2(G238), .ZN(n690) );
  NOR2_X1 U773 ( .A1(G235), .A2(G237), .ZN(n689) );
  NAND2_X1 U774 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U775 ( .A(KEYINPUT90), .B(n691), .ZN(n960) );
  NAND2_X1 U776 ( .A1(n960), .A2(G567), .ZN(n692) );
  NAND2_X1 U777 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U778 ( .A(KEYINPUT91), .B(n694), .ZN(G319) );
  INV_X1 U779 ( .A(G319), .ZN(n696) );
  NAND2_X1 U780 ( .A1(G661), .A2(G483), .ZN(n695) );
  NOR2_X1 U781 ( .A1(n696), .A2(n695), .ZN(n831) );
  NAND2_X1 U782 ( .A1(n831), .A2(G36), .ZN(G176) );
  INV_X1 U783 ( .A(G166), .ZN(G303) );
  NAND2_X1 U784 ( .A1(G40), .A2(G160), .ZN(n778) );
  INV_X1 U785 ( .A(n778), .ZN(n697) );
  NOR2_X1 U786 ( .A1(G164), .A2(G1384), .ZN(n779) );
  BUF_X2 U787 ( .A(n702), .Z(n739) );
  NAND2_X1 U788 ( .A1(G8), .A2(n739), .ZN(n769) );
  NOR2_X1 U789 ( .A1(G1981), .A2(G305), .ZN(n698) );
  XOR2_X1 U790 ( .A(n698), .B(KEYINPUT24), .Z(n699) );
  NOR2_X1 U791 ( .A1(n769), .A2(n699), .ZN(n777) );
  NAND2_X1 U792 ( .A1(G1348), .A2(n739), .ZN(n701) );
  INV_X1 U793 ( .A(n702), .ZN(n725) );
  NAND2_X1 U794 ( .A1(G2067), .A2(n725), .ZN(n700) );
  NAND2_X1 U795 ( .A1(n701), .A2(n700), .ZN(n709) );
  NOR2_X1 U796 ( .A1(n710), .A2(n709), .ZN(n708) );
  INV_X1 U797 ( .A(G1996), .ZN(n876) );
  NOR2_X1 U798 ( .A1(n702), .A2(n876), .ZN(n703) );
  XOR2_X1 U799 ( .A(n703), .B(KEYINPUT26), .Z(n706) );
  AND2_X1 U800 ( .A1(n739), .A2(G1341), .ZN(n704) );
  NOR2_X1 U801 ( .A1(n704), .A2(n1015), .ZN(n705) );
  AND2_X1 U802 ( .A1(n706), .A2(n705), .ZN(n707) );
  AND2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U804 ( .A1(n712), .A2(n711), .ZN(n717) );
  NAND2_X1 U805 ( .A1(n725), .A2(G2072), .ZN(n713) );
  XNOR2_X1 U806 ( .A(n713), .B(KEYINPUT27), .ZN(n715) );
  AND2_X1 U807 ( .A1(G1956), .A2(n739), .ZN(n714) );
  NOR2_X1 U808 ( .A1(G299), .A2(n719), .ZN(n716) );
  NOR2_X1 U809 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U810 ( .A(KEYINPUT97), .B(n718), .ZN(n722) );
  NAND2_X1 U811 ( .A1(G299), .A2(n719), .ZN(n720) );
  XNOR2_X1 U812 ( .A(KEYINPUT28), .B(n720), .ZN(n721) );
  AND2_X1 U813 ( .A1(n722), .A2(n721), .ZN(n724) );
  XNOR2_X1 U814 ( .A(KEYINPUT98), .B(KEYINPUT29), .ZN(n723) );
  XNOR2_X1 U815 ( .A(n724), .B(n723), .ZN(n729) );
  XOR2_X1 U816 ( .A(G1961), .B(KEYINPUT96), .Z(n921) );
  NAND2_X1 U817 ( .A1(n921), .A2(n739), .ZN(n727) );
  XNOR2_X1 U818 ( .A(G2078), .B(KEYINPUT25), .ZN(n882) );
  NAND2_X1 U819 ( .A1(n725), .A2(n882), .ZN(n726) );
  NAND2_X1 U820 ( .A1(n727), .A2(n726), .ZN(n733) );
  NAND2_X1 U821 ( .A1(G171), .A2(n733), .ZN(n728) );
  NAND2_X1 U822 ( .A1(n729), .A2(n728), .ZN(n738) );
  NOR2_X1 U823 ( .A1(G1966), .A2(n769), .ZN(n751) );
  NOR2_X1 U824 ( .A1(G2084), .A2(n739), .ZN(n748) );
  NOR2_X1 U825 ( .A1(n751), .A2(n748), .ZN(n730) );
  NAND2_X1 U826 ( .A1(G8), .A2(n730), .ZN(n731) );
  XNOR2_X1 U827 ( .A(KEYINPUT30), .B(n731), .ZN(n732) );
  NOR2_X1 U828 ( .A1(G168), .A2(n732), .ZN(n735) );
  NOR2_X1 U829 ( .A1(G171), .A2(n733), .ZN(n734) );
  NOR2_X1 U830 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U831 ( .A(KEYINPUT31), .B(n736), .Z(n737) );
  NAND2_X1 U832 ( .A1(n738), .A2(n737), .ZN(n749) );
  NAND2_X1 U833 ( .A1(n749), .A2(G286), .ZN(n744) );
  NOR2_X1 U834 ( .A1(G1971), .A2(n769), .ZN(n741) );
  NOR2_X1 U835 ( .A1(G2090), .A2(n739), .ZN(n740) );
  NOR2_X1 U836 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U837 ( .A1(n742), .A2(G303), .ZN(n743) );
  NAND2_X1 U838 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U839 ( .A1(n745), .A2(G8), .ZN(n747) );
  XOR2_X1 U840 ( .A(KEYINPUT32), .B(KEYINPUT99), .Z(n746) );
  XNOR2_X1 U841 ( .A(n747), .B(n746), .ZN(n755) );
  NAND2_X1 U842 ( .A1(G8), .A2(n748), .ZN(n753) );
  INV_X1 U843 ( .A(n749), .ZN(n750) );
  NOR2_X1 U844 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U845 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U846 ( .A1(n755), .A2(n754), .ZN(n766) );
  NOR2_X1 U847 ( .A1(G2090), .A2(G303), .ZN(n756) );
  NAND2_X1 U848 ( .A1(G8), .A2(n756), .ZN(n757) );
  NAND2_X1 U849 ( .A1(n766), .A2(n757), .ZN(n758) );
  XNOR2_X1 U850 ( .A(n758), .B(KEYINPUT102), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n759), .A2(n769), .ZN(n760) );
  XOR2_X1 U852 ( .A(KEYINPUT103), .B(n760), .Z(n775) );
  NOR2_X1 U853 ( .A1(G1976), .A2(G288), .ZN(n765) );
  NAND2_X1 U854 ( .A1(KEYINPUT33), .A2(n765), .ZN(n761) );
  NOR2_X1 U855 ( .A1(n769), .A2(n761), .ZN(n762) );
  XOR2_X1 U856 ( .A(KEYINPUT100), .B(n762), .Z(n773) );
  XOR2_X1 U857 ( .A(KEYINPUT101), .B(G1981), .Z(n763) );
  XNOR2_X1 U858 ( .A(G305), .B(n763), .ZN(n900) );
  NAND2_X1 U859 ( .A1(G1976), .A2(G288), .ZN(n903) );
  NOR2_X1 U860 ( .A1(G1971), .A2(G303), .ZN(n764) );
  NOR2_X1 U861 ( .A1(n765), .A2(n764), .ZN(n904) );
  NAND2_X1 U862 ( .A1(n904), .A2(n766), .ZN(n767) );
  NAND2_X1 U863 ( .A1(n903), .A2(n767), .ZN(n768) );
  NOR2_X1 U864 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U865 ( .A1(KEYINPUT33), .A2(n770), .ZN(n771) );
  NOR2_X1 U866 ( .A1(n900), .A2(n771), .ZN(n772) );
  NAND2_X1 U867 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U868 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U869 ( .A1(n777), .A2(n776), .ZN(n811) );
  NOR2_X1 U870 ( .A1(n779), .A2(n778), .ZN(n823) );
  NAND2_X1 U871 ( .A1(G140), .A2(n986), .ZN(n781) );
  NAND2_X1 U872 ( .A1(G104), .A2(n987), .ZN(n780) );
  NAND2_X1 U873 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U874 ( .A(KEYINPUT34), .B(n782), .ZN(n788) );
  NAND2_X1 U875 ( .A1(G116), .A2(n982), .ZN(n784) );
  NAND2_X1 U876 ( .A1(G128), .A2(n983), .ZN(n783) );
  NAND2_X1 U877 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U878 ( .A(KEYINPUT35), .B(n785), .Z(n786) );
  XNOR2_X1 U879 ( .A(KEYINPUT94), .B(n786), .ZN(n787) );
  NOR2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U881 ( .A(KEYINPUT36), .B(n789), .ZN(n1009) );
  XOR2_X1 U882 ( .A(G2067), .B(KEYINPUT37), .Z(n790) );
  XNOR2_X1 U883 ( .A(KEYINPUT93), .B(n790), .ZN(n821) );
  NOR2_X1 U884 ( .A1(n1009), .A2(n821), .ZN(n866) );
  NAND2_X1 U885 ( .A1(n823), .A2(n866), .ZN(n818) );
  NAND2_X1 U886 ( .A1(n986), .A2(G131), .ZN(n793) );
  NAND2_X1 U887 ( .A1(G95), .A2(n987), .ZN(n791) );
  XOR2_X1 U888 ( .A(KEYINPUT95), .B(n791), .Z(n792) );
  NAND2_X1 U889 ( .A1(n793), .A2(n792), .ZN(n797) );
  NAND2_X1 U890 ( .A1(G107), .A2(n982), .ZN(n795) );
  NAND2_X1 U891 ( .A1(G119), .A2(n983), .ZN(n794) );
  NAND2_X1 U892 ( .A1(n795), .A2(n794), .ZN(n796) );
  OR2_X1 U893 ( .A1(n797), .A2(n796), .ZN(n999) );
  AND2_X1 U894 ( .A1(n999), .A2(G1991), .ZN(n806) );
  NAND2_X1 U895 ( .A1(G141), .A2(n986), .ZN(n799) );
  NAND2_X1 U896 ( .A1(G129), .A2(n983), .ZN(n798) );
  NAND2_X1 U897 ( .A1(n799), .A2(n798), .ZN(n802) );
  NAND2_X1 U898 ( .A1(n987), .A2(G105), .ZN(n800) );
  XOR2_X1 U899 ( .A(KEYINPUT38), .B(n800), .Z(n801) );
  NOR2_X1 U900 ( .A1(n802), .A2(n801), .ZN(n804) );
  NAND2_X1 U901 ( .A1(n982), .A2(G117), .ZN(n803) );
  NAND2_X1 U902 ( .A1(n804), .A2(n803), .ZN(n1004) );
  AND2_X1 U903 ( .A1(n1004), .A2(G1996), .ZN(n805) );
  NOR2_X1 U904 ( .A1(n806), .A2(n805), .ZN(n855) );
  INV_X1 U905 ( .A(n823), .ZN(n807) );
  NOR2_X1 U906 ( .A1(n855), .A2(n807), .ZN(n814) );
  INV_X1 U907 ( .A(n814), .ZN(n808) );
  NAND2_X1 U908 ( .A1(n818), .A2(n808), .ZN(n809) );
  XNOR2_X1 U909 ( .A(G1986), .B(G290), .ZN(n912) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n1004), .ZN(n857) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n812) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n999), .ZN(n850) );
  NOR2_X1 U913 ( .A1(n812), .A2(n850), .ZN(n813) );
  NOR2_X1 U914 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U915 ( .A(n815), .B(KEYINPUT104), .ZN(n816) );
  NOR2_X1 U916 ( .A1(n857), .A2(n816), .ZN(n817) );
  XNOR2_X1 U917 ( .A(n817), .B(KEYINPUT39), .ZN(n819) );
  NAND2_X1 U918 ( .A1(n819), .A2(n818), .ZN(n820) );
  XOR2_X1 U919 ( .A(KEYINPUT105), .B(n820), .Z(n822) );
  NAND2_X1 U920 ( .A1(n1009), .A2(n821), .ZN(n863) );
  NAND2_X1 U921 ( .A1(n822), .A2(n863), .ZN(n824) );
  NAND2_X1 U922 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U923 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U924 ( .A(KEYINPUT40), .B(n827), .ZN(G329) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n828), .ZN(G217) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U927 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U929 ( .A1(n831), .A2(n830), .ZN(G188) );
  NAND2_X1 U931 ( .A1(G136), .A2(n986), .ZN(n833) );
  NAND2_X1 U932 ( .A1(G100), .A2(n987), .ZN(n832) );
  NAND2_X1 U933 ( .A1(n833), .A2(n832), .ZN(n838) );
  NAND2_X1 U934 ( .A1(G124), .A2(n983), .ZN(n834) );
  XNOR2_X1 U935 ( .A(n834), .B(KEYINPUT44), .ZN(n836) );
  NAND2_X1 U936 ( .A1(n982), .A2(G112), .ZN(n835) );
  NAND2_X1 U937 ( .A1(n836), .A2(n835), .ZN(n837) );
  NOR2_X1 U938 ( .A1(n838), .A2(n837), .ZN(G162) );
  NAND2_X1 U939 ( .A1(G139), .A2(n986), .ZN(n840) );
  NAND2_X1 U940 ( .A1(G103), .A2(n987), .ZN(n839) );
  NAND2_X1 U941 ( .A1(n840), .A2(n839), .ZN(n846) );
  NAND2_X1 U942 ( .A1(G115), .A2(n982), .ZN(n842) );
  NAND2_X1 U943 ( .A1(G127), .A2(n983), .ZN(n841) );
  NAND2_X1 U944 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U945 ( .A(KEYINPUT47), .B(n843), .ZN(n844) );
  XNOR2_X1 U946 ( .A(KEYINPUT111), .B(n844), .ZN(n845) );
  NOR2_X1 U947 ( .A1(n846), .A2(n845), .ZN(n998) );
  XOR2_X1 U948 ( .A(G2072), .B(n998), .Z(n848) );
  XOR2_X1 U949 ( .A(G164), .B(G2078), .Z(n847) );
  NOR2_X1 U950 ( .A1(n848), .A2(n847), .ZN(n849) );
  XOR2_X1 U951 ( .A(KEYINPUT50), .B(n849), .Z(n869) );
  NOR2_X1 U952 ( .A1(n850), .A2(n995), .ZN(n851) );
  XOR2_X1 U953 ( .A(KEYINPUT116), .B(n851), .Z(n853) );
  XOR2_X1 U954 ( .A(G2084), .B(G160), .Z(n852) );
  NOR2_X1 U955 ( .A1(n853), .A2(n852), .ZN(n854) );
  NAND2_X1 U956 ( .A1(n855), .A2(n854), .ZN(n862) );
  XOR2_X1 U957 ( .A(G2090), .B(G162), .Z(n856) );
  NOR2_X1 U958 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U959 ( .A(KEYINPUT51), .B(n858), .Z(n860) );
  XNOR2_X1 U960 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(n861) );
  NOR2_X1 U962 ( .A1(n862), .A2(n861), .ZN(n864) );
  NAND2_X1 U963 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U964 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U965 ( .A(KEYINPUT119), .B(n867), .ZN(n868) );
  NOR2_X1 U966 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U967 ( .A(KEYINPUT52), .B(n870), .ZN(n871) );
  INV_X1 U968 ( .A(KEYINPUT55), .ZN(n894) );
  NAND2_X1 U969 ( .A1(n871), .A2(n894), .ZN(n872) );
  NAND2_X1 U970 ( .A1(n872), .A2(G29), .ZN(n952) );
  XNOR2_X1 U971 ( .A(G1991), .B(G25), .ZN(n874) );
  XNOR2_X1 U972 ( .A(G33), .B(G2072), .ZN(n873) );
  NOR2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n881) );
  XOR2_X1 U974 ( .A(G2067), .B(G26), .Z(n875) );
  NAND2_X1 U975 ( .A1(n875), .A2(G28), .ZN(n879) );
  XOR2_X1 U976 ( .A(G32), .B(n876), .Z(n877) );
  XNOR2_X1 U977 ( .A(KEYINPUT120), .B(n877), .ZN(n878) );
  NOR2_X1 U978 ( .A1(n879), .A2(n878), .ZN(n880) );
  NAND2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n884) );
  XOR2_X1 U980 ( .A(G27), .B(n882), .Z(n883) );
  NOR2_X1 U981 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U982 ( .A(n885), .B(KEYINPUT121), .Z(n886) );
  XNOR2_X1 U983 ( .A(KEYINPUT53), .B(n886), .ZN(n888) );
  XNOR2_X1 U984 ( .A(G35), .B(G2090), .ZN(n887) );
  NOR2_X1 U985 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U986 ( .A(n889), .B(KEYINPUT122), .ZN(n892) );
  XOR2_X1 U987 ( .A(G2084), .B(KEYINPUT54), .Z(n890) );
  XNOR2_X1 U988 ( .A(G34), .B(n890), .ZN(n891) );
  NAND2_X1 U989 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U990 ( .A(n894), .B(n893), .ZN(n896) );
  INV_X1 U991 ( .A(G29), .ZN(n895) );
  NAND2_X1 U992 ( .A1(n896), .A2(n895), .ZN(n897) );
  NAND2_X1 U993 ( .A1(G11), .A2(n897), .ZN(n950) );
  INV_X1 U994 ( .A(G16), .ZN(n946) );
  XNOR2_X1 U995 ( .A(KEYINPUT56), .B(KEYINPUT123), .ZN(n898) );
  XNOR2_X1 U996 ( .A(n946), .B(n898), .ZN(n920) );
  XOR2_X1 U997 ( .A(G1966), .B(G168), .Z(n899) );
  NOR2_X1 U998 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U999 ( .A(KEYINPUT57), .B(n901), .Z(n918) );
  XNOR2_X1 U1000 ( .A(n1012), .B(G1348), .ZN(n914) );
  INV_X1 U1001 ( .A(G1971), .ZN(n902) );
  NOR2_X1 U1002 ( .A1(G166), .A2(n902), .ZN(n906) );
  NAND2_X1 U1003 ( .A1(n904), .A2(n903), .ZN(n905) );
  NOR2_X1 U1004 ( .A1(n906), .A2(n905), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(G301), .B(G1961), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n1015), .B(G1341), .ZN(n907) );
  NOR2_X1 U1007 ( .A1(n908), .A2(n907), .ZN(n909) );
  NAND2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(n911) );
  NOR2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(G1956), .B(G299), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1013 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1014 ( .A1(n920), .A2(n919), .ZN(n948) );
  XOR2_X1 U1015 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n944) );
  XOR2_X1 U1016 ( .A(G1966), .B(G21), .Z(n923) );
  XNOR2_X1 U1017 ( .A(n921), .B(G5), .ZN(n922) );
  NAND2_X1 U1018 ( .A1(n923), .A2(n922), .ZN(n930) );
  XNOR2_X1 U1019 ( .A(G1976), .B(G23), .ZN(n925) );
  XNOR2_X1 U1020 ( .A(G1971), .B(G22), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n927) );
  XOR2_X1 U1022 ( .A(G1986), .B(G24), .Z(n926) );
  NAND2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1024 ( .A(KEYINPUT58), .B(n928), .ZN(n929) );
  NOR2_X1 U1025 ( .A1(n930), .A2(n929), .ZN(n942) );
  XNOR2_X1 U1026 ( .A(G1348), .B(KEYINPUT59), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(n931), .B(G4), .ZN(n935) );
  XNOR2_X1 U1028 ( .A(G1981), .B(G6), .ZN(n933) );
  XNOR2_X1 U1029 ( .A(G19), .B(G1341), .ZN(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n938) );
  XNOR2_X1 U1032 ( .A(KEYINPUT124), .B(G1956), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(G20), .B(n936), .ZN(n937) );
  NOR2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1035 ( .A(n939), .B(KEYINPUT125), .Z(n940) );
  XNOR2_X1 U1036 ( .A(KEYINPUT60), .B(n940), .ZN(n941) );
  NAND2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(n944), .B(n943), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1040 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1041 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1042 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1043 ( .A(KEYINPUT62), .B(n953), .Z(G311) );
  XNOR2_X1 U1044 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  XOR2_X1 U1045 ( .A(n954), .B(KEYINPUT83), .Z(n958) );
  NAND2_X1 U1046 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1047 ( .A(n958), .B(n957), .ZN(G145) );
  INV_X1 U1048 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1049 ( .A1(n960), .A2(n959), .ZN(G325) );
  INV_X1 U1050 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1051 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n962) );
  XNOR2_X1 U1052 ( .A(G1986), .B(G1976), .ZN(n961) );
  XNOR2_X1 U1053 ( .A(n962), .B(n961), .ZN(n963) );
  XOR2_X1 U1054 ( .A(n963), .B(G1956), .Z(n965) );
  XNOR2_X1 U1055 ( .A(G1981), .B(G1961), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(n965), .B(n964), .ZN(n969) );
  XOR2_X1 U1057 ( .A(KEYINPUT41), .B(G2474), .Z(n967) );
  XNOR2_X1 U1058 ( .A(G1971), .B(G1966), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(n967), .B(n966), .ZN(n968) );
  XOR2_X1 U1060 ( .A(n969), .B(n968), .Z(n971) );
  XNOR2_X1 U1061 ( .A(G1996), .B(G1991), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(n971), .B(n970), .ZN(G229) );
  XOR2_X1 U1063 ( .A(KEYINPUT106), .B(G2678), .Z(n973) );
  XNOR2_X1 U1064 ( .A(G2072), .B(G2090), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(n973), .B(n972), .ZN(n977) );
  XOR2_X1 U1066 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n975) );
  XNOR2_X1 U1067 ( .A(G2067), .B(KEYINPUT42), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(n975), .B(n974), .ZN(n976) );
  XOR2_X1 U1069 ( .A(n977), .B(n976), .Z(n979) );
  XNOR2_X1 U1070 ( .A(G2096), .B(G2100), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(n979), .B(n978), .ZN(n981) );
  XOR2_X1 U1072 ( .A(G2078), .B(G2084), .Z(n980) );
  XNOR2_X1 U1073 ( .A(n981), .B(n980), .ZN(G227) );
  NAND2_X1 U1074 ( .A1(G118), .A2(n982), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(G130), .A2(n983), .ZN(n984) );
  NAND2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n993) );
  NAND2_X1 U1077 ( .A1(G142), .A2(n986), .ZN(n989) );
  NAND2_X1 U1078 ( .A1(G106), .A2(n987), .ZN(n988) );
  NAND2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1080 ( .A(KEYINPUT45), .B(n990), .Z(n991) );
  XNOR2_X1 U1081 ( .A(KEYINPUT110), .B(n991), .ZN(n992) );
  NOR2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(n995), .B(n994), .ZN(n1008) );
  XOR2_X1 U1084 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n997) );
  XNOR2_X1 U1085 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(n997), .B(n996), .ZN(n1003) );
  XOR2_X1 U1087 ( .A(G162), .B(n998), .Z(n1001) );
  XOR2_X1 U1088 ( .A(G164), .B(n999), .Z(n1000) );
  XNOR2_X1 U1089 ( .A(n1001), .B(n1000), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(n1003), .B(n1002), .ZN(n1006) );
  XOR2_X1 U1091 ( .A(G160), .B(n1004), .Z(n1005) );
  XNOR2_X1 U1092 ( .A(n1006), .B(n1005), .ZN(n1007) );
  XNOR2_X1 U1093 ( .A(n1008), .B(n1007), .ZN(n1010) );
  XOR2_X1 U1094 ( .A(n1010), .B(n1009), .Z(n1011) );
  NOR2_X1 U1095 ( .A1(G37), .A2(n1011), .ZN(G395) );
  XNOR2_X1 U1096 ( .A(n1012), .B(G286), .ZN(n1014) );
  XNOR2_X1 U1097 ( .A(n1014), .B(n1013), .ZN(n1017) );
  XOR2_X1 U1098 ( .A(n1015), .B(G171), .Z(n1016) );
  XNOR2_X1 U1099 ( .A(n1017), .B(n1016), .ZN(n1018) );
  NOR2_X1 U1100 ( .A1(G37), .A2(n1018), .ZN(G397) );
  NOR2_X1 U1101 ( .A1(G229), .A2(G227), .ZN(n1020) );
  XNOR2_X1 U1102 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n1019) );
  XNOR2_X1 U1103 ( .A(n1020), .B(n1019), .ZN(n1021) );
  NOR2_X1 U1104 ( .A1(G401), .A2(n1021), .ZN(n1022) );
  NAND2_X1 U1105 ( .A1(G319), .A2(n1022), .ZN(n1023) );
  XNOR2_X1 U1106 ( .A(KEYINPUT115), .B(n1023), .ZN(n1025) );
  NOR2_X1 U1107 ( .A1(G395), .A2(G397), .ZN(n1024) );
  NAND2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(G225) );
  INV_X1 U1109 ( .A(G225), .ZN(G308) );
endmodule

