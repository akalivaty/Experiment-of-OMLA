//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  NAND2_X1  g000(.A1(G234), .A2(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(G952), .A3(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT92), .ZN(new_n190));
  AND3_X1   g004(.A1(new_n187), .A2(G902), .A3(G953), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT21), .B(G898), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n190), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(G214), .B1(G237), .B2(G902), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n196), .B(KEYINPUT80), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT64), .B1(new_n198), .B2(G146), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(G146), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n205));
  AND4_X1   g019(.A1(new_n199), .A2(new_n202), .A3(new_n203), .A4(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n201), .A2(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(new_n203), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT67), .B(G128), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT1), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n210), .B1(G143), .B2(new_n201), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n208), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT68), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT68), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n208), .B(new_n214), .C1(new_n209), .C2(new_n211), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n206), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G125), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT0), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(new_n204), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n204), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n208), .A3(new_n222), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n199), .A2(new_n220), .A3(new_n202), .A4(new_n203), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G125), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n218), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G224), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(G953), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT7), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n233));
  INV_X1    g047(.A(G104), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n233), .B1(new_n234), .B2(G107), .ZN(new_n235));
  INV_X1    g049(.A(G107), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT3), .A3(G104), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(KEYINPUT75), .B1(new_n236), .B2(G104), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT75), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(new_n234), .A3(G107), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G101), .ZN(new_n243));
  INV_X1    g057(.A(G101), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n238), .A2(new_n244), .A3(new_n239), .A4(new_n241), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n243), .A2(KEYINPUT4), .A3(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(G116), .B(G119), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT2), .B(G113), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n247), .B(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n242), .A2(new_n251), .A3(G101), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n246), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n234), .A2(G107), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n236), .A2(G104), .ZN(new_n255));
  OAI21_X1  g069(.A(G101), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n245), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n247), .ZN(new_n258));
  OR2_X1    g072(.A1(new_n258), .A2(new_n248), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT81), .B(KEYINPUT5), .ZN(new_n260));
  INV_X1    g074(.A(G119), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(G116), .A3(new_n261), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n262), .B(G113), .C1(new_n258), .C2(new_n260), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n257), .A2(new_n259), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(G110), .B(G122), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n253), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n218), .A2(KEYINPUT7), .A3(new_n226), .A4(new_n230), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n232), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n265), .B(KEYINPUT8), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT84), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n262), .A2(new_n270), .A3(G113), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n270), .B1(new_n262), .B2(G113), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n247), .A2(KEYINPUT5), .ZN(new_n273));
  NOR3_X1   g087(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n257), .A2(new_n259), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT85), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n263), .A2(new_n259), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n245), .A2(new_n256), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NOR3_X1   g094(.A1(new_n274), .A2(new_n275), .A3(KEYINPUT85), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n269), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(G902), .B1(new_n268), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n227), .B(new_n229), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n253), .A2(new_n264), .ZN(new_n285));
  XOR2_X1   g099(.A(new_n265), .B(KEYINPUT82), .Z(new_n286));
  AND2_X1   g100(.A1(new_n286), .A2(KEYINPUT83), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n285), .A2(KEYINPUT6), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n266), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT6), .B1(new_n285), .B2(new_n287), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n284), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n283), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G210), .B1(G237), .B2(G902), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n283), .A2(new_n291), .A3(new_n293), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n197), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n195), .B1(new_n297), .B2(KEYINPUT86), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n298), .B1(KEYINPUT86), .B2(new_n297), .ZN(new_n299));
  INV_X1    g113(.A(G469), .ZN(new_n300));
  INV_X1    g114(.A(G902), .ZN(new_n301));
  XNOR2_X1  g115(.A(G110), .B(G140), .ZN(new_n302));
  INV_X1    g116(.A(G227), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n303), .A2(G953), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n302), .B(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n225), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n246), .A2(new_n307), .A3(new_n252), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT10), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n278), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n199), .A2(new_n202), .A3(new_n203), .A4(new_n205), .ZN(new_n311));
  INV_X1    g125(.A(new_n215), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT1), .B1(new_n198), .B2(G146), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT67), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(G128), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n204), .A2(KEYINPUT67), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n214), .B1(new_n317), .B2(new_n208), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n311), .B1(new_n312), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n310), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n199), .A2(new_n202), .A3(new_n203), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n313), .A2(G128), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(new_n311), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(new_n245), .A3(new_n256), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT76), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n325), .A2(new_n326), .A3(new_n309), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n326), .B1(new_n325), .B2(new_n309), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n308), .B(new_n320), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT79), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G137), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n332), .A2(G134), .B1(KEYINPUT65), .B2(KEYINPUT11), .ZN(new_n333));
  OR2_X1    g147(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n332), .A2(G134), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT66), .ZN(new_n338));
  AND2_X1   g152(.A1(KEYINPUT11), .A2(G134), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n338), .B1(new_n339), .B2(new_n332), .ZN(new_n340));
  NAND2_X1  g154(.A1(KEYINPUT11), .A2(G134), .ZN(new_n341));
  NOR3_X1   g155(.A1(new_n341), .A2(KEYINPUT66), .A3(G137), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n335), .B(new_n337), .C1(new_n340), .C2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G131), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n339), .A2(new_n338), .A3(new_n332), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT66), .B1(new_n341), .B2(G137), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n336), .A2(G131), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n335), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n320), .A2(new_n308), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n206), .B1(new_n321), .B2(new_n322), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n309), .B1(new_n352), .B2(new_n278), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT76), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n325), .A2(new_n326), .A3(new_n309), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n351), .A2(new_n356), .A3(KEYINPUT79), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n331), .A2(new_n350), .A3(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n350), .B(KEYINPUT77), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n351), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n306), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n306), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n345), .A2(new_n346), .B1(new_n333), .B2(new_n334), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n343), .A2(G131), .B1(new_n363), .B2(new_n348), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n278), .B(new_n311), .C1(new_n318), .C2(new_n312), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n364), .B1(new_n365), .B2(new_n325), .ZN(new_n366));
  NOR3_X1   g180(.A1(new_n366), .A2(KEYINPUT78), .A3(KEYINPUT12), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT12), .ZN(new_n369));
  AOI211_X1 g183(.A(new_n369), .B(new_n364), .C1(new_n365), .C2(new_n325), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n365), .A2(new_n325), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n350), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n369), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n370), .B1(new_n373), .B2(KEYINPUT78), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n362), .B1(new_n368), .B2(new_n374), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n300), .B(new_n301), .C1(new_n361), .C2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(G469), .A2(G902), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n356), .A2(new_n351), .A3(new_n359), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n364), .B1(new_n329), .B2(new_n330), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n378), .B1(new_n379), .B2(new_n357), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n306), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n366), .A2(KEYINPUT12), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n366), .A2(KEYINPUT12), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT78), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n360), .B1(new_n385), .B2(new_n367), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n305), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n381), .A2(G469), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n376), .A2(new_n377), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT20), .ZN(new_n390));
  INV_X1    g204(.A(G237), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(new_n188), .A3(G214), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n198), .ZN(new_n393));
  NOR2_X1   g207(.A1(G237), .A2(G953), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(G143), .A3(G214), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(KEYINPUT18), .A3(G131), .ZN(new_n397));
  XNOR2_X1  g211(.A(G125), .B(G140), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(new_n201), .ZN(new_n399));
  NAND2_X1  g213(.A1(KEYINPUT18), .A2(G131), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n393), .A2(new_n395), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT87), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n402), .B(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(G113), .B(G122), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(new_n234), .ZN(new_n406));
  INV_X1    g220(.A(G140), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G125), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n217), .A2(G140), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(KEYINPUT16), .ZN(new_n410));
  OR3_X1    g224(.A1(new_n217), .A2(KEYINPUT16), .A3(G140), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(G146), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT73), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT73), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n410), .A2(new_n411), .A3(new_n414), .A4(G146), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n410), .A2(new_n411), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n201), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n413), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n394), .A2(G143), .A3(G214), .ZN(new_n419));
  AOI21_X1  g233(.A(G143), .B1(new_n394), .B2(G214), .ZN(new_n420));
  OAI211_X1 g234(.A(KEYINPUT17), .B(G131), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT88), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT88), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n396), .A2(new_n423), .A3(KEYINPUT17), .A4(G131), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n418), .A2(KEYINPUT89), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G131), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n396), .B(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT17), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(KEYINPUT89), .B1(new_n418), .B2(new_n425), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n404), .B(new_n406), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n402), .A2(new_n403), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n402), .A2(new_n403), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n398), .B(KEYINPUT19), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n412), .B1(new_n437), .B2(G146), .ZN(new_n438));
  OAI22_X1  g252(.A1(new_n434), .A2(new_n435), .B1(new_n428), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n406), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n433), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(G475), .A2(G902), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n390), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n443), .ZN(new_n445));
  AOI211_X1 g259(.A(KEYINPUT20), .B(new_n445), .C1(new_n433), .C2(new_n441), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n404), .B1(new_n431), .B2(new_n432), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n440), .ZN(new_n448));
  AOI21_X1  g262(.A(G902), .B1(new_n448), .B2(new_n433), .ZN(new_n449));
  INV_X1    g263(.A(G475), .ZN(new_n450));
  OAI22_X1  g264(.A1(new_n444), .A2(new_n446), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT71), .B(G217), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT9), .B(G234), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n452), .A2(new_n453), .A3(G953), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n209), .A2(G143), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT91), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT91), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n209), .A2(new_n458), .A3(G143), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G134), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n198), .A2(G128), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G116), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n464), .A2(G122), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n464), .A2(KEYINPUT90), .A3(G122), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT90), .B1(new_n464), .B2(G122), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(G107), .ZN(new_n469));
  XOR2_X1   g283(.A(new_n462), .B(KEYINPUT13), .Z(new_n470));
  AOI21_X1  g284(.A(new_n470), .B1(new_n457), .B2(new_n459), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n463), .B(new_n469), .C1(new_n461), .C2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n236), .B1(new_n465), .B2(KEYINPUT14), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n468), .B(new_n474), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n209), .A2(new_n458), .A3(G143), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n458), .B1(new_n209), .B2(G143), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n462), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G134), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n475), .B1(new_n479), .B2(new_n463), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n455), .B1(new_n473), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n475), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n478), .A2(G134), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n461), .B1(new_n460), .B2(new_n462), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(new_n472), .A3(new_n454), .ZN(new_n486));
  AOI21_X1  g300(.A(G902), .B1(new_n481), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G478), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n487), .B(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n451), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(G221), .B1(new_n453), .B2(G902), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n389), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n299), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT30), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n461), .A2(G137), .ZN(new_n497));
  OAI21_X1  g311(.A(G131), .B1(new_n497), .B2(new_n336), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n349), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n213), .A2(new_n215), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n499), .B1(new_n500), .B2(new_n311), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n225), .B1(new_n344), .B2(new_n349), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n496), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n349), .A2(new_n498), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n319), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n427), .B1(new_n363), .B2(new_n337), .ZN(new_n506));
  INV_X1    g320(.A(new_n349), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n307), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n505), .A2(KEYINPUT30), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n503), .A2(new_n509), .A3(new_n250), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n505), .A2(new_n508), .A3(new_n249), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n394), .A2(G210), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT27), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT26), .B(G101), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  NOR3_X1   g332(.A1(new_n501), .A2(new_n502), .A3(new_n250), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n249), .B1(new_n505), .B2(new_n508), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT28), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT28), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n511), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n516), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT29), .B1(new_n518), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n516), .A2(KEYINPUT29), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n301), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(G472), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT32), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT30), .B1(new_n216), .B2(new_n499), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n250), .B1(new_n531), .B2(new_n502), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT30), .B1(new_n505), .B2(new_n508), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n511), .B(new_n516), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT69), .B1(new_n534), .B2(KEYINPUT31), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n519), .A2(new_n517), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT69), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT31), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n536), .A2(new_n510), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n524), .A2(new_n517), .B1(KEYINPUT31), .B2(new_n534), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(G472), .A2(G902), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n530), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n543), .ZN(new_n545));
  AOI211_X1 g359(.A(KEYINPUT32), .B(new_n545), .C1(new_n540), .C2(new_n541), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n529), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT70), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g363(.A(KEYINPUT70), .B(new_n529), .C1(new_n544), .C2(new_n546), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n452), .B1(G234), .B2(new_n301), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n413), .A2(new_n415), .A3(new_n417), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n209), .A2(G119), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n261), .A2(G128), .ZN(new_n555));
  XOR2_X1   g369(.A(KEYINPUT24), .B(G110), .Z(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT23), .B1(new_n204), .B2(G119), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n559), .B1(new_n261), .B2(G128), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT72), .B1(new_n561), .B2(G110), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT72), .ZN(new_n563));
  INV_X1    g377(.A(G110), .ZN(new_n564));
  AOI211_X1 g378(.A(new_n563), .B(new_n564), .C1(new_n558), .C2(new_n560), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n553), .B(new_n557), .C1(new_n562), .C2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n398), .A2(new_n201), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n561), .A2(G110), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n556), .B1(new_n554), .B2(new_n555), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n412), .B(new_n567), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT22), .B(G137), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n573));
  XOR2_X1   g387(.A(new_n572), .B(new_n573), .Z(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n566), .A2(new_n570), .A3(new_n574), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(new_n301), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT25), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n576), .A2(KEYINPUT25), .A3(new_n301), .A4(new_n577), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n552), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n577), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n574), .B1(new_n566), .B2(new_n570), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n551), .A2(G902), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n582), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n549), .A2(new_n550), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT74), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT74), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n549), .A2(new_n593), .A3(new_n550), .A4(new_n590), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n495), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(new_n244), .ZN(G3));
  INV_X1    g410(.A(G472), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n542), .B2(new_n301), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n542), .A2(new_n543), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n590), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n389), .A2(new_n493), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n283), .A2(new_n291), .A3(new_n293), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n293), .B1(new_n283), .B2(new_n291), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n196), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n485), .A2(new_n472), .A3(new_n454), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n454), .B1(new_n485), .B2(new_n472), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n488), .B(new_n301), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n488), .A2(new_n301), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(KEYINPUT33), .B1(new_n608), .B2(new_n609), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n481), .A2(new_n615), .A3(new_n486), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n613), .B1(new_n617), .B2(G478), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n451), .A2(new_n618), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n607), .A2(new_n619), .A3(new_n194), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n603), .A2(new_n604), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT34), .B(G104), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  NAND2_X1  g437(.A1(new_n442), .A2(new_n443), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT20), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n442), .A2(new_n390), .A3(new_n443), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(KEYINPUT93), .A3(new_n626), .ZN(new_n627));
  OR2_X1    g441(.A1(new_n626), .A2(KEYINPUT93), .ZN(new_n628));
  OR2_X1    g442(.A1(new_n449), .A2(new_n450), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n627), .A2(new_n628), .A3(new_n629), .A4(new_n491), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n630), .A2(new_n607), .A3(new_n194), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n603), .A2(new_n604), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NAND2_X1  g448(.A1(new_n580), .A2(new_n581), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n551), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n571), .A2(KEYINPUT94), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT94), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n566), .A2(new_n638), .A3(new_n570), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n575), .A2(KEYINPUT36), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n637), .A2(new_n641), .A3(new_n639), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n587), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n636), .A2(KEYINPUT95), .A3(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT95), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n588), .B1(new_n643), .B2(new_n644), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n648), .B1(new_n582), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g466(.A(KEYINPUT96), .B1(new_n601), .B2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT96), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n599), .A2(new_n651), .A3(new_n654), .A4(new_n600), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n299), .A2(new_n653), .A3(new_n655), .A4(new_n494), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT37), .B(G110), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G12));
  AND3_X1   g472(.A1(new_n389), .A2(new_n651), .A3(new_n493), .ZN(new_n659));
  INV_X1    g473(.A(G900), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n191), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n190), .A2(new_n661), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n630), .A2(new_n607), .A3(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n549), .A2(new_n659), .A3(new_n550), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT97), .B(G128), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G30));
  XOR2_X1   g480(.A(new_n662), .B(KEYINPUT39), .Z(new_n667));
  NAND2_X1  g481(.A1(new_n604), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT40), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n604), .A2(KEYINPUT40), .A3(new_n667), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n670), .A2(KEYINPUT100), .A3(new_n671), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n519), .A2(new_n520), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n516), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n677), .A2(KEYINPUT99), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n534), .B1(new_n677), .B2(KEYINPUT99), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n301), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(G472), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n681), .B1(new_n544), .B2(new_n546), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n605), .A2(new_n606), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n196), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n451), .A2(new_n491), .ZN(new_n688));
  NOR4_X1   g502(.A1(new_n686), .A2(new_n687), .A3(new_n651), .A4(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n674), .A2(new_n675), .A3(new_n682), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT101), .B(G143), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G45));
  NAND3_X1  g506(.A1(new_n614), .A2(new_n616), .A3(G478), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n610), .A3(new_n612), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n625), .A2(new_n626), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n694), .B1(new_n695), .B2(new_n629), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n687), .B1(new_n295), .B2(new_n296), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT102), .ZN(new_n698));
  INV_X1    g512(.A(new_n662), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n696), .A2(new_n697), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n451), .A2(new_n618), .A3(new_n699), .ZN(new_n701));
  OAI21_X1  g515(.A(KEYINPUT102), .B1(new_n701), .B2(new_n607), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n703), .A2(new_n549), .A3(new_n550), .A4(new_n659), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT103), .B(G146), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G48));
  OAI21_X1  g520(.A(new_n301), .B1(new_n361), .B2(new_n375), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(G469), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n493), .A3(new_n376), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n709), .A2(KEYINPUT104), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(KEYINPUT104), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n620), .A3(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n591), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT105), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n713), .B(new_n715), .ZN(G15));
  NAND3_X1  g530(.A1(new_n710), .A2(new_n631), .A3(new_n711), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n591), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n464), .ZN(G18));
  NOR2_X1   g533(.A1(new_n709), .A2(new_n607), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n651), .A2(new_n195), .A3(new_n492), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(new_n549), .A3(new_n550), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  NAND2_X1  g537(.A1(new_n600), .A2(KEYINPUT106), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n542), .A2(new_n725), .A3(new_n543), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n598), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n590), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n607), .A2(new_n688), .A3(new_n194), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n729), .A2(new_n711), .A3(new_n710), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  INV_X1    g546(.A(new_n701), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n720), .A2(new_n651), .A3(new_n733), .A4(new_n727), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G125), .ZN(G27));
  NAND4_X1  g549(.A1(new_n547), .A2(KEYINPUT42), .A3(new_n590), .A4(new_n733), .ZN(new_n736));
  XOR2_X1   g550(.A(new_n377), .B(KEYINPUT107), .Z(new_n737));
  AND2_X1   g551(.A1(new_n376), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n378), .B1(new_n374), .B2(new_n368), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n739), .B1(new_n740), .B2(new_n306), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n386), .A2(KEYINPUT108), .A3(new_n305), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n741), .A2(G469), .A3(new_n381), .A4(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n387), .A2(new_n739), .B1(new_n380), .B2(new_n306), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(KEYINPUT109), .A3(G469), .A4(new_n742), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n738), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n683), .A2(new_n196), .ZN(new_n749));
  INV_X1    g563(.A(new_n493), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n748), .A2(KEYINPUT110), .A3(new_n751), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n736), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n549), .A2(new_n550), .A3(new_n590), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT110), .B1(new_n748), .B2(new_n751), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n748), .A2(KEYINPUT110), .A3(new_n751), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n757), .B(new_n733), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(KEYINPUT111), .B(KEYINPUT42), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n756), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n427), .ZN(G33));
  NOR2_X1   g577(.A1(new_n630), .A2(new_n662), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n757), .B(new_n764), .C1(new_n758), .C2(new_n759), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G134), .ZN(G36));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n746), .A2(KEYINPUT45), .A3(new_n742), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n381), .A2(new_n387), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n300), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(KEYINPUT46), .A3(new_n737), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(KEYINPUT112), .A3(new_n376), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n737), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT46), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT112), .B1(new_n773), .B2(new_n376), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n493), .ZN(new_n781));
  INV_X1    g595(.A(new_n667), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n767), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n451), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n618), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n785), .B(KEYINPUT43), .Z(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n601), .A3(new_n651), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n789), .A2(new_n790), .A3(new_n749), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n780), .A2(KEYINPUT113), .A3(new_n493), .A4(new_n667), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n783), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  NAND2_X1  g608(.A1(new_n549), .A2(new_n550), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NOR4_X1   g610(.A1(new_n796), .A2(new_n590), .A3(new_n701), .A4(new_n749), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n780), .A2(KEYINPUT47), .A3(new_n493), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT47), .B1(new_n780), .B2(new_n493), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n797), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G140), .ZN(G42));
  NOR4_X1   g616(.A1(new_n785), .A2(new_n602), .A3(new_n197), .A4(new_n750), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT114), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n708), .A2(new_n376), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT49), .Z(new_n806));
  OR4_X1    g620(.A1(new_n682), .A2(new_n804), .A3(new_n685), .A4(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n190), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n786), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(new_n728), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n685), .A2(new_n196), .A3(new_n709), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT50), .ZN(new_n813));
  INV_X1    g627(.A(new_n749), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n805), .A2(new_n493), .A3(new_n814), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n815), .A2(new_n602), .A3(new_n190), .A4(new_n682), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n784), .A3(new_n694), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n809), .A2(new_n815), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n727), .A2(new_n651), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n818), .A2(KEYINPUT119), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT119), .B1(new_n818), .B2(new_n820), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n817), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n813), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n800), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n805), .A2(new_n750), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n825), .A2(new_n798), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n810), .A2(new_n814), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT117), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n827), .A2(new_n828), .ZN(new_n833));
  OAI211_X1 g647(.A(KEYINPUT51), .B(new_n824), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  XOR2_X1   g648(.A(new_n826), .B(KEYINPUT118), .Z(new_n835));
  NAND3_X1  g649(.A1(new_n825), .A2(new_n798), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n831), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT51), .B1(new_n837), .B2(new_n824), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n547), .A2(new_n590), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n818), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT48), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n810), .A2(new_n720), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n188), .A2(G952), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(new_n816), .B2(new_n696), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n841), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n838), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n834), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n299), .A2(new_n604), .A3(new_n603), .A4(new_n696), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n592), .A2(new_n594), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n848), .B(new_n849), .C1(new_n850), .C2(new_n495), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n784), .A2(new_n491), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n299), .A2(new_n604), .A3(new_n603), .A4(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n731), .A2(new_n656), .A3(new_n853), .A4(new_n722), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n591), .B1(new_n717), .B2(new_n712), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n849), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT115), .B1(new_n595), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n851), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n733), .B(new_n820), .C1(new_n759), .C2(new_n758), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n627), .A2(new_n629), .A3(new_n628), .ZN(new_n861));
  NOR4_X1   g675(.A1(new_n749), .A2(new_n861), .A3(new_n491), .A4(new_n662), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n796), .A2(new_n659), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n765), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n762), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n607), .A2(new_n688), .ZN(new_n867));
  NOR4_X1   g681(.A1(new_n582), .A2(new_n649), .A3(new_n750), .A4(new_n662), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n748), .A2(new_n867), .A3(new_n682), .A4(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n704), .A2(new_n664), .A3(new_n734), .A4(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT52), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT116), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n704), .A2(new_n664), .A3(new_n734), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(KEYINPUT52), .A3(new_n869), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n874), .A2(KEYINPUT116), .A3(KEYINPUT52), .A4(new_n869), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT53), .B1(new_n866), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n762), .A2(new_n864), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n880), .A2(new_n851), .A3(new_n858), .A4(new_n856), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT53), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n875), .A2(new_n872), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT54), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n882), .B1(new_n881), .B2(new_n883), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n851), .A2(new_n858), .A3(new_n856), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n887), .A2(new_n878), .A3(KEYINPUT53), .A4(new_n880), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n885), .B1(KEYINPUT54), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n847), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(G952), .A2(G953), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n807), .B1(new_n891), .B2(new_n892), .ZN(G75));
  INV_X1    g707(.A(KEYINPUT56), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n889), .A2(G902), .ZN(new_n895));
  INV_X1    g709(.A(G210), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n289), .A2(new_n290), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(new_n284), .Z(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT55), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n900), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n894), .B(new_n902), .C1(new_n895), .C2(new_n896), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n188), .A2(G952), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n901), .A2(new_n903), .A3(new_n905), .ZN(G51));
  XOR2_X1   g720(.A(new_n737), .B(KEYINPUT57), .Z(new_n907));
  NOR2_X1   g721(.A1(new_n889), .A2(KEYINPUT54), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT54), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(new_n886), .B2(new_n888), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n907), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n361), .A2(new_n375), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n895), .A2(new_n772), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n904), .B1(new_n913), .B2(new_n914), .ZN(G54));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n916));
  NAND2_X1  g730(.A1(KEYINPUT58), .A2(G475), .ZN(new_n917));
  AOI211_X1 g731(.A(new_n301), .B(new_n917), .C1(new_n886), .C2(new_n888), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n905), .B1(new_n918), .B2(new_n442), .ZN(new_n919));
  INV_X1    g733(.A(new_n917), .ZN(new_n920));
  AND4_X1   g734(.A1(G902), .A2(new_n889), .A3(new_n442), .A4(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n916), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n442), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n923), .B1(new_n895), .B2(new_n917), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n918), .A2(new_n442), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n924), .A2(new_n925), .A3(KEYINPUT121), .A4(new_n905), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n922), .A2(new_n926), .ZN(G60));
  NOR2_X1   g741(.A1(new_n908), .A2(new_n910), .ZN(new_n928));
  INV_X1    g742(.A(new_n617), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n611), .B(KEYINPUT59), .Z(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n905), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n929), .B1(new_n890), .B2(new_n930), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(G63));
  NAND2_X1  g748(.A1(G217), .A2(G902), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT60), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n889), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n904), .B1(new_n938), .B2(new_n586), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n936), .B1(new_n886), .B2(new_n888), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n645), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n939), .B(new_n941), .C1(new_n942), .C2(KEYINPUT61), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT61), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n942), .B(new_n905), .C1(new_n940), .C2(new_n585), .ZN(new_n945));
  INV_X1    g759(.A(new_n941), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n905), .B1(new_n940), .B2(new_n585), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n944), .B(new_n945), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n943), .A2(new_n948), .ZN(G66));
  NAND2_X1  g763(.A1(new_n859), .A2(new_n188), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(G953), .B1(new_n192), .B2(new_n228), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(KEYINPUT124), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n188), .A2(G898), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n289), .A2(new_n290), .A3(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT124), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n952), .A2(new_n958), .A3(new_n953), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n955), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n957), .B1(new_n955), .B2(new_n959), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n960), .A2(new_n961), .ZN(G69));
  OAI21_X1  g776(.A(G953), .B1(new_n303), .B2(new_n660), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n503), .A2(new_n509), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT125), .Z(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(new_n436), .ZN(new_n966));
  NAND2_X1  g780(.A1(G900), .A2(G953), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n783), .A2(new_n867), .A3(new_n839), .A4(new_n792), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n874), .A2(new_n765), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n762), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n968), .A2(new_n793), .A3(new_n801), .A4(new_n970), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n966), .B(new_n967), .C1(new_n971), .C2(G953), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT126), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n690), .A2(new_n874), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n974), .B1(new_n975), .B2(KEYINPUT62), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT62), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n690), .A2(KEYINPUT126), .A3(new_n977), .A4(new_n874), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n814), .B1(new_n852), .B2(new_n696), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n850), .A2(new_n668), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n975), .B2(KEYINPUT62), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n979), .A2(new_n793), .A3(new_n801), .A4(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n966), .B1(new_n983), .B2(new_n188), .ZN(new_n984));
  OAI211_X1 g798(.A(KEYINPUT127), .B(new_n963), .C1(new_n973), .C2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n984), .ZN(new_n986));
  OR2_X1    g800(.A1(new_n963), .A2(KEYINPUT127), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n963), .A2(KEYINPUT127), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n986), .A2(new_n972), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n985), .A2(new_n989), .ZN(G72));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT63), .Z(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n983), .B2(new_n859), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n512), .A2(new_n517), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n992), .B1(new_n971), .B2(new_n859), .ZN(new_n996));
  INV_X1    g810(.A(new_n518), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n992), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n997), .A2(new_n999), .A3(new_n994), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n1000), .B1(new_n879), .B2(new_n884), .ZN(new_n1001));
  AND4_X1   g815(.A1(new_n905), .A2(new_n995), .A3(new_n998), .A4(new_n1001), .ZN(G57));
endmodule


