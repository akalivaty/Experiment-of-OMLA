//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 0 1 1 0 0 0 1 1 1 0 1 1 0 0 1 0 1 0 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1230, new_n1231,
    new_n1232, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G50), .ZN(new_n203));
  INV_X1    g0003(.A(G77), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n202), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(new_n213), .A2(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  INV_X1    g0022(.A(G97), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  INV_X1    g0026(.A(G50), .ZN(new_n227));
  INV_X1    g0027(.A(G226), .ZN(new_n228));
  INV_X1    g0028(.A(G244), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n204), .C2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n211), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n219), .B1(new_n214), .B2(new_n213), .C1(new_n231), .C2(KEYINPUT1), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT65), .ZN(new_n243));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  OAI21_X1  g0049(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n250));
  INV_X1    g0050(.A(G274), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  OAI211_X1 g0055(.A(G1), .B(G13), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n250), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n253), .B1(new_n257), .B2(new_n228), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT3), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n254), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G223), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(new_n262), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G222), .A3(new_n259), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n264), .B(new_n266), .C1(new_n204), .C2(new_n265), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n258), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G200), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n271), .B(KEYINPUT69), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n208), .A2(G13), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(new_n209), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G50), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n210), .A2(G33), .B1(G1), .B2(G13), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n276), .B1(G1), .B2(new_n209), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n275), .B1(new_n277), .B2(G50), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n203), .A2(new_n209), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n280), .B1(G150), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT8), .B(G58), .ZN(new_n283));
  OR2_X1    g0083(.A1(new_n283), .A2(KEYINPUT66), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(KEYINPUT66), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n284), .A2(new_n209), .A3(G33), .A4(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g0087(.A(KEYINPUT9), .B(new_n279), .C1(new_n287), .C2(new_n276), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT9), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n276), .B1(new_n282), .B2(new_n286), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n289), .B1(new_n290), .B2(new_n278), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n269), .A2(G190), .ZN(new_n292));
  AND2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n272), .A2(new_n288), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT70), .B1(new_n294), .B2(KEYINPUT10), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT69), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n271), .B(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n288), .A2(new_n292), .A3(new_n291), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT70), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT10), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n295), .A2(new_n302), .B1(KEYINPUT10), .B2(new_n294), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n269), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(G179), .B2(new_n269), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n279), .B1(new_n287), .B2(new_n276), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G232), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n253), .B1(new_n257), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n263), .A2(G226), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n265), .A2(G223), .A3(new_n259), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n313), .B(new_n314), .C1(new_n254), .C2(new_n221), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n312), .B1(new_n315), .B2(new_n268), .ZN(new_n316));
  INV_X1    g0116(.A(G179), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n316), .A2(G169), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G68), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT7), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n265), .B2(G20), .ZN(new_n323));
  AND2_X1   g0123(.A1(KEYINPUT3), .A2(G33), .ZN(new_n324));
  NOR2_X1   g0124(.A1(KEYINPUT3), .A2(G33), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n321), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G58), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(new_n321), .ZN(new_n330));
  OAI21_X1  g0130(.A(G20), .B1(new_n330), .B2(new_n201), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n281), .A2(G159), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT16), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n333), .B2(KEYINPUT75), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n336), .B1(new_n328), .B2(new_n333), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n276), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n284), .A2(new_n285), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n341), .A2(new_n274), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(new_n277), .B2(new_n341), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n320), .B(KEYINPUT18), .C1(new_n340), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT76), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n338), .A2(new_n339), .ZN(new_n346));
  INV_X1    g0146(.A(new_n276), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n343), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT76), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n350), .A2(new_n351), .A3(KEYINPUT18), .A4(new_n320), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT18), .ZN(new_n353));
  INV_X1    g0153(.A(new_n320), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n340), .A2(new_n343), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n345), .A2(new_n352), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G190), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n316), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(G200), .B2(new_n316), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n348), .A2(new_n349), .A3(new_n360), .ZN(new_n361));
  XNOR2_X1  g0161(.A(new_n361), .B(KEYINPUT17), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n263), .A2(G238), .ZN(new_n364));
  INV_X1    g0164(.A(G107), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n265), .A2(new_n259), .ZN(new_n366));
  OAI221_X1 g0166(.A(new_n364), .B1(new_n365), .B2(new_n265), .C1(new_n311), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n268), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n368), .B(new_n253), .C1(new_n229), .C2(new_n257), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n369), .A2(G190), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n370), .B1(new_n270), .B2(new_n369), .ZN(new_n371));
  XNOR2_X1  g0171(.A(KEYINPUT15), .B(G87), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n209), .A2(G33), .ZN(new_n373));
  OAI22_X1  g0173(.A1(new_n372), .A2(new_n373), .B1(new_n209), .B2(new_n204), .ZN(new_n374));
  INV_X1    g0174(.A(new_n281), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n283), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n347), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT67), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n274), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n204), .ZN(new_n381));
  INV_X1    g0181(.A(new_n277), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n381), .B1(new_n382), .B2(new_n204), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT68), .ZN(new_n385));
  XNOR2_X1  g0185(.A(new_n384), .B(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n371), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n369), .A2(G169), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n317), .B2(new_n369), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n363), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  NOR3_X1   g0191(.A1(new_n273), .A2(new_n209), .A3(G68), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n392), .B(KEYINPUT12), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n382), .B2(G68), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n281), .A2(G50), .B1(G20), .B2(new_n321), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n204), .B2(new_n373), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n347), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT11), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n399), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n395), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n263), .A2(G232), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G97), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n405), .B(new_n406), .C1(new_n228), .C2(new_n366), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n268), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n257), .A2(KEYINPUT71), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n257), .A2(KEYINPUT71), .ZN(new_n410));
  OAI21_X1  g0210(.A(G238), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(new_n411), .A3(new_n253), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT13), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n413), .A2(KEYINPUT72), .ZN(new_n414));
  XOR2_X1   g0214(.A(new_n412), .B(new_n414), .Z(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G179), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n412), .A2(new_n413), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT14), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n408), .A2(new_n411), .A3(KEYINPUT13), .A4(new_n253), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n417), .A2(new_n418), .A3(G169), .A4(new_n419), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n420), .A2(KEYINPUT74), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(KEYINPUT74), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n416), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n417), .A2(G169), .A3(new_n419), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT73), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n424), .A2(new_n425), .A3(KEYINPUT14), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(new_n424), .B2(KEYINPUT14), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n404), .B1(new_n423), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n415), .A2(G190), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n417), .A2(G200), .A3(new_n419), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n430), .A2(new_n403), .A3(new_n431), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n310), .A2(new_n391), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n273), .A2(new_n209), .A3(G107), .ZN(new_n436));
  XOR2_X1   g0236(.A(KEYINPUT84), .B(KEYINPUT25), .Z(new_n437));
  NOR2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n437), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n438), .B1(KEYINPUT85), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(KEYINPUT85), .B2(new_n439), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n208), .A2(G33), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n276), .A2(new_n380), .A3(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n441), .B1(new_n365), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n209), .A2(G107), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT23), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G116), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n209), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n265), .A2(new_n209), .A3(G87), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n451), .A2(KEYINPUT22), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(KEYINPUT22), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n454), .A2(KEYINPUT24), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n276), .B1(new_n454), .B2(KEYINPUT24), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n444), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT88), .ZN(new_n459));
  OAI211_X1 g0259(.A(G257), .B(G1698), .C1(new_n324), .C2(new_n325), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT86), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT86), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n265), .A2(new_n462), .A3(G257), .A4(G1698), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n222), .A2(G1698), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(new_n324), .B2(new_n325), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT87), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n265), .A2(KEYINPUT87), .A3(new_n465), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G294), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n268), .B1(new_n464), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G45), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(G1), .ZN(new_n474));
  AND2_X1   g0274(.A1(KEYINPUT5), .A2(G41), .ZN(new_n475));
  NOR2_X1   g0275(.A1(KEYINPUT5), .A2(G41), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n477), .A2(new_n256), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G264), .ZN(new_n479));
  OR2_X1    g0279(.A1(new_n477), .A2(new_n251), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n472), .A2(G179), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n472), .A2(new_n479), .A3(new_n480), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n459), .A2(new_n481), .B1(new_n482), .B2(G169), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n482), .A2(new_n459), .A3(G169), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT89), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n481), .A2(new_n459), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n482), .A2(G169), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n482), .A2(new_n459), .A3(G169), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT89), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n458), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT90), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n263), .A2(KEYINPUT83), .A3(G264), .ZN(new_n494));
  INV_X1    g0294(.A(G303), .ZN(new_n495));
  OAI221_X1 g0295(.A(new_n494), .B1(new_n495), .B2(new_n265), .C1(new_n224), .C2(new_n366), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT83), .B1(new_n263), .B2(G264), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n268), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT82), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n499), .B1(new_n478), .B2(G270), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n477), .A2(new_n499), .A3(G270), .A4(new_n256), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n480), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n443), .A2(G116), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(G116), .B2(new_n274), .ZN(new_n506));
  INV_X1    g0306(.A(G116), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n209), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G283), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n223), .B2(G33), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n508), .B1(new_n510), .B2(new_n209), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT20), .ZN(new_n512));
  OR3_X1    g0312(.A1(new_n511), .A2(new_n276), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n511), .B2(new_n276), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n304), .B1(new_n506), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n504), .A2(KEYINPUT21), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n506), .A2(new_n515), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n518), .A2(new_n498), .A3(G179), .A4(new_n503), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n498), .A2(new_n358), .A3(new_n503), .ZN(new_n522));
  AOI21_X1  g0322(.A(G200), .B1(new_n498), .B2(new_n503), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n515), .B(new_n506), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(KEYINPUT21), .B1(new_n504), .B2(new_n516), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n265), .A2(new_n209), .A3(G68), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT19), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n209), .B1(new_n406), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(G87), .A2(G97), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n365), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT80), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n528), .B1(new_n406), .B2(G20), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n527), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n529), .B2(new_n531), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n347), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OR2_X1    g0337(.A1(new_n443), .A2(new_n221), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n274), .A2(new_n372), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(G250), .B1(new_n473), .B2(G1), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n474), .A2(G274), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n268), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n265), .A2(G238), .A3(new_n259), .ZN(new_n544));
  OAI211_X1 g0344(.A(G244), .B(G1698), .C1(new_n324), .C2(new_n325), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(new_n447), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n543), .B1(new_n546), .B2(new_n268), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n540), .B1(G190), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n268), .ZN(new_n549));
  INV_X1    g0349(.A(new_n543), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G200), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n547), .A2(G179), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n304), .B2(new_n547), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT81), .ZN(new_n555));
  XNOR2_X1  g0355(.A(new_n372), .B(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n556), .A2(new_n276), .A3(new_n380), .A4(new_n442), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n537), .A2(new_n557), .A3(new_n539), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n548), .A2(new_n552), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n521), .A2(new_n524), .A3(new_n526), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n263), .A2(G250), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT4), .ZN(new_n562));
  AOI21_X1  g0362(.A(G1698), .B1(new_n562), .B2(KEYINPUT78), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(KEYINPUT78), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n265), .A2(G244), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n561), .A2(new_n565), .A3(new_n509), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n229), .B1(new_n261), .B2(new_n262), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n564), .B1(new_n567), .B2(new_n563), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n268), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT79), .ZN(new_n570));
  INV_X1    g0370(.A(new_n480), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n571), .B1(G257), .B2(new_n478), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT79), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n573), .B(new_n268), .C1(new_n566), .C2(new_n568), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n570), .A2(new_n317), .A3(new_n572), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n572), .A2(new_n569), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n304), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OR2_X1    g0379(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n580));
  NAND2_X1  g0380(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n580), .B(new_n581), .C1(new_n223), .C2(G107), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n580), .A2(new_n581), .ZN(new_n583));
  XNOR2_X1  g0383(.A(G97), .B(G107), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n582), .B(G20), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n204), .B2(new_n375), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n365), .B1(new_n323), .B2(new_n327), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n347), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n443), .A2(G97), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(G97), .B2(new_n274), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n579), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n576), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n591), .B1(new_n593), .B2(G190), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n570), .A2(new_n572), .A3(new_n574), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G200), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n560), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n485), .B1(new_n483), .B2(new_n484), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n489), .A2(KEYINPUT89), .A3(new_n490), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n457), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT90), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n482), .A2(new_n270), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n482), .A2(G190), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n457), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n493), .A2(new_n599), .A3(new_n604), .A4(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n435), .A2(new_n608), .ZN(G372));
  INV_X1    g0409(.A(new_n429), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n432), .A2(new_n390), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n362), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n356), .A2(new_n344), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n300), .B1(new_n299), .B2(new_n301), .ZN(new_n615));
  NOR4_X1   g0415(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT70), .A4(KEYINPUT10), .ZN(new_n616));
  OAI22_X1  g0416(.A1(new_n615), .A2(new_n616), .B1(new_n301), .B2(new_n299), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n309), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n448), .B1(new_n567), .B2(G1698), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n256), .B1(new_n619), .B2(new_n544), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n620), .A2(new_n317), .A3(new_n543), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n304), .B1(new_n549), .B2(new_n550), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n558), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT91), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(new_n547), .B2(new_n270), .ZN(new_n625));
  OAI211_X1 g0425(.A(KEYINPUT91), .B(G200), .C1(new_n620), .C2(new_n543), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n547), .A2(G190), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n628), .A2(new_n539), .A3(new_n537), .A4(new_n538), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n623), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT92), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n623), .B(KEYINPUT92), .C1(new_n627), .C2(new_n629), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n578), .A2(KEYINPUT94), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT94), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n575), .A2(new_n577), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n634), .A2(new_n638), .A3(new_n639), .A4(new_n591), .ZN(new_n640));
  INV_X1    g0440(.A(new_n623), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n559), .A2(new_n579), .A3(new_n591), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n641), .B1(new_n642), .B2(KEYINPUT26), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT95), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT95), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n640), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n634), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n592), .A2(new_n597), .A3(new_n607), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT93), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n520), .B2(new_n525), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n526), .A2(KEYINPUT93), .A3(new_n517), .A4(new_n519), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n458), .B1(new_n484), .B2(new_n483), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n645), .A2(new_n647), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n618), .B1(new_n435), .B2(new_n659), .ZN(G369));
  OR3_X1    g0460(.A1(new_n273), .A2(KEYINPUT27), .A3(G20), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT27), .B1(new_n273), .B2(G20), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G213), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(G343), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n458), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n493), .A2(new_n604), .A3(new_n607), .A4(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n602), .A2(new_n665), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n654), .A2(new_n518), .A3(new_n665), .ZN(new_n670));
  INV_X1    g0470(.A(G330), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n520), .A2(new_n525), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n672), .A2(new_n524), .B1(new_n518), .B2(new_n665), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n670), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n655), .A2(new_n665), .ZN(new_n676));
  INV_X1    g0476(.A(new_n665), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n520), .B2(new_n525), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n667), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n675), .A2(new_n676), .A3(new_n679), .ZN(G399));
  INV_X1    g0480(.A(new_n212), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(G41), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n530), .A2(new_n365), .A3(new_n507), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(G1), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n217), .B2(new_n683), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n623), .B1(new_n642), .B2(KEYINPUT26), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n634), .A2(new_n591), .A3(new_n638), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n689), .B1(new_n690), .B2(KEYINPUT26), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT97), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n602), .A2(new_n603), .ZN(new_n693));
  AOI211_X1 g0493(.A(KEYINPUT90), .B(new_n457), .C1(new_n600), .C2(new_n601), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n692), .B1(new_n695), .B2(new_n672), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n493), .A2(new_n692), .A3(new_n604), .A4(new_n672), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n650), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n691), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(KEYINPUT29), .A3(new_n677), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n659), .B2(new_n665), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT31), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n472), .A2(new_n479), .A3(new_n547), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n593), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n498), .A2(G179), .A3(new_n503), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n705), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n708), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(KEYINPUT30), .A3(new_n593), .A4(new_n706), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  AOI211_X1 g0512(.A(G179), .B(new_n547), .C1(new_n498), .C2(new_n503), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(new_n482), .A3(new_n595), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT96), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n714), .A2(KEYINPUT96), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n712), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n704), .B1(new_n719), .B2(new_n677), .ZN(new_n720));
  OAI211_X1 g0520(.A(KEYINPUT31), .B(new_n665), .C1(new_n712), .C2(new_n715), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n720), .B(new_n721), .C1(new_n608), .C2(new_n665), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n722), .A2(G330), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n703), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n688), .B1(new_n724), .B2(G1), .ZN(G364));
  NOR2_X1   g0525(.A1(G13), .A2(G33), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G20), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(new_n670), .B2(new_n673), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n209), .A2(G13), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G45), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n683), .A2(G1), .A3(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT98), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n209), .A2(new_n358), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n270), .A2(G179), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n209), .A2(G190), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G179), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI22_X1  g0545(.A1(G303), .A2(new_n741), .B1(new_n745), .B2(G329), .ZN(new_n746));
  INV_X1    g0546(.A(G283), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n739), .A2(new_n742), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n746), .B(new_n326), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n209), .B1(new_n743), .B2(G190), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n749), .B1(G294), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n317), .A2(new_n270), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n738), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G326), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n317), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n738), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G322), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n754), .A2(new_n755), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  XOR2_X1   g0559(.A(KEYINPUT33), .B(G317), .Z(new_n760));
  NAND2_X1  g0560(.A1(new_n753), .A2(new_n742), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n756), .A2(new_n742), .ZN(new_n762));
  INV_X1    g0562(.A(G311), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n760), .A2(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n762), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G77), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n767), .B1(new_n227), .B2(new_n754), .C1(new_n321), .C2(new_n761), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT32), .ZN(new_n769));
  INV_X1    g0569(.A(G159), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n769), .B1(new_n744), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n745), .A2(KEYINPUT32), .A3(G159), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n768), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n265), .B1(new_n740), .B2(new_n221), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n757), .A2(new_n329), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n748), .A2(new_n365), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n750), .A2(new_n223), .ZN(new_n777));
  NOR4_X1   g0577(.A1(new_n774), .A2(new_n775), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n752), .A2(new_n765), .B1(new_n773), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n215), .B1(G20), .B2(new_n304), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n737), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n728), .A2(new_n780), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n681), .A2(new_n265), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n245), .A2(new_n473), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n218), .A2(G45), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n681), .A2(new_n326), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n789), .A2(G355), .B1(new_n507), .B2(new_n681), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n784), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n782), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n729), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT99), .Z(new_n794));
  NOR2_X1   g0594(.A1(new_n674), .A2(new_n737), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n671), .B1(new_n670), .B2(new_n673), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(G396));
  NOR2_X1   g0599(.A1(new_n780), .A2(new_n726), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n736), .B1(new_n204), .B2(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G107), .A2(new_n741), .B1(new_n745), .B2(G311), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n802), .B(new_n326), .C1(new_n221), .C2(new_n748), .ZN(new_n803));
  INV_X1    g0603(.A(G294), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n757), .A2(new_n804), .B1(new_n762), .B2(new_n507), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n754), .A2(new_n495), .B1(new_n761), .B2(new_n747), .ZN(new_n806));
  NOR4_X1   g0606(.A1(new_n803), .A2(new_n777), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n754), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n808), .A2(G137), .B1(new_n766), .B2(G159), .ZN(new_n809));
  INV_X1    g0609(.A(G143), .ZN(new_n810));
  INV_X1    g0610(.A(G150), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n809), .B1(new_n810), .B2(new_n757), .C1(new_n811), .C2(new_n761), .ZN(new_n812));
  XOR2_X1   g0612(.A(KEYINPUT100), .B(KEYINPUT34), .Z(new_n813));
  XNOR2_X1  g0613(.A(new_n812), .B(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n265), .B1(new_n740), .B2(new_n227), .ZN(new_n815));
  INV_X1    g0615(.A(G132), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n748), .A2(new_n321), .B1(new_n744), .B2(new_n816), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n815), .B(new_n817), .C1(G58), .C2(new_n751), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n807), .B1(new_n814), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n390), .A2(new_n387), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n386), .A2(new_n665), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n386), .A2(new_n389), .ZN(new_n822));
  OAI21_X1  g0622(.A(KEYINPUT101), .B1(new_n822), .B2(new_n677), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT101), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n386), .A2(new_n824), .A3(new_n389), .A4(new_n665), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n820), .A2(new_n821), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n801), .B1(new_n781), .B2(new_n819), .C1(new_n827), .C2(new_n727), .ZN(new_n828));
  AOI22_X1  g0628(.A1(KEYINPUT95), .A2(new_n644), .B1(new_n650), .B2(new_n656), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n665), .B1(new_n829), .B2(new_n647), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(new_n826), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n723), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n832), .A2(KEYINPUT102), .A3(new_n736), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n723), .B2(new_n831), .ZN(new_n834));
  AOI21_X1  g0634(.A(KEYINPUT102), .B1(new_n832), .B2(new_n736), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n828), .B1(new_n834), .B2(new_n835), .ZN(G384));
  NAND3_X1  g0636(.A1(new_n700), .A2(new_n434), .A3(new_n702), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n618), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT105), .ZN(new_n839));
  INV_X1    g0639(.A(new_n663), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n613), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n334), .B(new_n335), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n347), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n349), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n840), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n363), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT103), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n355), .B1(new_n354), .B2(new_n663), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n361), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n848), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n350), .B1(new_n320), .B2(new_n840), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n853), .A2(new_n361), .A3(KEYINPUT103), .A4(new_n850), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n844), .B1(new_n320), .B2(new_n840), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n361), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT37), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n847), .A2(new_n859), .A3(KEYINPUT38), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n852), .A2(new_n854), .B1(new_n857), .B2(KEYINPUT37), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n845), .B1(new_n357), .B2(new_n362), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT39), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT104), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n361), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n355), .A2(KEYINPUT104), .A3(new_n360), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n853), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n852), .A2(new_n854), .B1(new_n870), .B2(KEYINPUT37), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n350), .A2(new_n840), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n362), .B2(new_n613), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n861), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT39), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n860), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n866), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n429), .A2(new_n665), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n841), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n404), .A2(new_n665), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n429), .A2(new_n432), .A3(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n404), .B(new_n665), .C1(new_n423), .C2(new_n428), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n658), .A2(new_n677), .A3(new_n827), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n822), .A2(new_n665), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n884), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n865), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n879), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n839), .B(new_n891), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n714), .B(new_n716), .ZN(new_n893));
  OAI211_X1 g0693(.A(KEYINPUT31), .B(new_n665), .C1(new_n893), .C2(new_n712), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n894), .B(new_n720), .C1(new_n608), .C2(new_n665), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n826), .B1(new_n881), .B2(new_n882), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT40), .B1(new_n860), .B2(new_n864), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n860), .A2(new_n874), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n899), .A2(new_n895), .A3(new_n896), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n897), .A2(new_n898), .B1(new_n900), .B2(KEYINPUT40), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n434), .A2(new_n895), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n901), .B(new_n902), .Z(new_n903));
  NOR2_X1   g0703(.A1(new_n903), .A2(new_n671), .ZN(new_n904));
  OAI22_X1  g0704(.A1(new_n892), .A2(new_n904), .B1(new_n208), .B2(new_n730), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n892), .B2(new_n904), .ZN(new_n906));
  OR3_X1    g0706(.A1(new_n217), .A2(new_n204), .A3(new_n330), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n227), .A2(G68), .ZN(new_n908));
  AOI211_X1 g0708(.A(new_n208), .B(G13), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n583), .A2(new_n584), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n910), .A2(new_n582), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n911), .A2(KEYINPUT35), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(KEYINPUT35), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n912), .A2(G116), .A3(new_n216), .A4(new_n913), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT36), .Z(new_n915));
  OR3_X1    g0715(.A1(new_n906), .A2(new_n909), .A3(new_n915), .ZN(G367));
  NAND2_X1  g0716(.A1(new_n591), .A2(new_n665), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n592), .A2(new_n597), .A3(new_n917), .ZN(new_n918));
  OR3_X1    g0718(.A1(new_n679), .A2(KEYINPUT42), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT42), .B1(new_n679), .B2(new_n918), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n638), .A2(new_n591), .A3(new_n665), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n695), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n592), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n677), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n919), .A2(new_n920), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n540), .A2(new_n665), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n648), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n641), .B2(new_n926), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n925), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT106), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n934), .A2(new_n935), .B1(new_n925), .B2(new_n930), .ZN(new_n936));
  INV_X1    g0736(.A(new_n675), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n921), .A2(new_n918), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n936), .B(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n682), .B(KEYINPUT41), .Z(new_n942));
  NAND3_X1  g0742(.A1(new_n679), .A2(new_n676), .A3(new_n938), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT45), .Z(new_n944));
  AOI21_X1  g0744(.A(new_n938), .B1(new_n679), .B2(new_n676), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT44), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(new_n675), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n669), .A2(new_n674), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n937), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(new_n678), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n724), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT107), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n952), .A2(KEYINPUT107), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n948), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n942), .B1(new_n956), .B2(new_n724), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n731), .A2(G1), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n941), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NOR3_X1   g0759(.A1(new_n240), .A2(new_n681), .A3(new_n265), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n783), .B1(new_n212), .B2(new_n372), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n804), .A2(new_n761), .B1(new_n757), .B2(new_n495), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n265), .B(new_n962), .C1(G317), .C2(new_n745), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n751), .A2(G107), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n741), .A2(G116), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT46), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n754), .A2(new_n763), .B1(new_n762), .B2(new_n747), .ZN(new_n967));
  INV_X1    g0767(.A(new_n748), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n967), .B1(G97), .B2(new_n968), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n963), .A2(new_n964), .A3(new_n966), .A4(new_n969), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n754), .A2(new_n810), .B1(new_n757), .B2(new_n811), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n761), .A2(new_n770), .B1(new_n762), .B2(new_n227), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n751), .A2(G68), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n326), .B1(new_n741), .B2(G58), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n748), .A2(new_n204), .ZN(new_n976));
  XNOR2_X1  g0776(.A(KEYINPUT108), .B(G137), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n976), .B1(new_n745), .B2(new_n978), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n973), .A2(new_n974), .A3(new_n975), .A4(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n970), .A2(KEYINPUT47), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n780), .ZN(new_n982));
  AOI21_X1  g0782(.A(KEYINPUT47), .B1(new_n970), .B2(new_n980), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n737), .B1(new_n960), .B2(new_n961), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT109), .Z(new_n985));
  INV_X1    g0785(.A(new_n728), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n985), .B1(new_n929), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n959), .A2(new_n987), .ZN(G387));
  NAND2_X1  g0788(.A1(new_n951), .A2(new_n958), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n283), .A2(G50), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT50), .Z(new_n991));
  OAI211_X1 g0791(.A(new_n685), .B(new_n473), .C1(new_n321), .C2(new_n204), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n785), .B1(new_n991), .B2(new_n992), .C1(new_n237), .C2(new_n473), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n789), .A2(new_n684), .B1(new_n365), .B2(new_n681), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n556), .A2(new_n751), .ZN(new_n996));
  INV_X1    g0796(.A(new_n341), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n996), .B1(new_n997), .B2(new_n761), .ZN(new_n998));
  INV_X1    g0798(.A(new_n757), .ZN(new_n999));
  AOI22_X1  g0799(.A1(G50), .A2(new_n999), .B1(new_n766), .B2(G68), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n770), .B2(new_n754), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(G77), .A2(new_n741), .B1(new_n745), .B2(G150), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1002), .B(new_n265), .C1(new_n223), .C2(new_n748), .ZN(new_n1003));
  NOR3_X1   g0803(.A1(new_n998), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT110), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n741), .A2(G294), .B1(new_n751), .B2(G283), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n808), .A2(G322), .B1(new_n766), .B2(G303), .ZN(new_n1007));
  INV_X1    g0807(.A(G317), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1007), .B1(new_n763), .B2(new_n761), .C1(new_n1008), .C2(new_n757), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT48), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1006), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT111), .Z(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n1010), .B2(new_n1009), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1013), .A2(KEYINPUT49), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n326), .B1(new_n744), .B2(new_n755), .C1(new_n507), .C2(new_n748), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n1013), .B2(KEYINPUT49), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1005), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n737), .B1(new_n784), .B2(new_n995), .C1(new_n1017), .C2(new_n781), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT112), .Z(new_n1019));
  NOR2_X1   g0819(.A1(new_n669), .A2(new_n986), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n952), .A2(new_n682), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n724), .A2(new_n951), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n989), .B1(new_n1019), .B2(new_n1020), .C1(new_n1021), .C2(new_n1022), .ZN(G393));
  XNOR2_X1  g0823(.A(new_n947), .B(new_n937), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n683), .B1(new_n1024), .B2(new_n952), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n956), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n948), .A2(new_n958), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n754), .A2(new_n811), .B1(new_n757), .B2(new_n770), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT51), .Z(new_n1029));
  OAI22_X1  g0829(.A1(new_n761), .A2(new_n227), .B1(new_n744), .B2(new_n810), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n740), .A2(new_n321), .B1(new_n762), .B2(new_n283), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n265), .B1(new_n750), .B2(new_n204), .C1(new_n221), .C2(new_n748), .ZN(new_n1032));
  OR4_X1    g0832(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n754), .A2(new_n1008), .B1(new_n757), .B2(new_n763), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT52), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n740), .A2(new_n747), .B1(new_n762), .B2(new_n804), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n761), .A2(new_n495), .B1(new_n744), .B2(new_n758), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n265), .B(new_n776), .C1(G116), .C2(new_n751), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1035), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n781), .B1(new_n1033), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n783), .B1(new_n223), .B2(new_n212), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n785), .B2(new_n248), .ZN(new_n1043));
  NOR3_X1   g0843(.A1(new_n1041), .A2(new_n736), .A3(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n938), .B2(new_n986), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1026), .A2(new_n1027), .A3(new_n1045), .ZN(G390));
  OAI211_X1 g0846(.A(new_n866), .B(new_n876), .C1(new_n888), .C2(new_n878), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n722), .A2(new_n883), .A3(G330), .A4(new_n827), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n699), .A2(new_n677), .A3(new_n827), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n884), .B1(new_n1049), .B2(new_n887), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n878), .B1(new_n860), .B2(new_n874), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1047), .B(new_n1048), .C1(new_n1050), .C2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n885), .A2(new_n887), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n883), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n878), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n877), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1049), .A2(new_n887), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n883), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1057), .B1(new_n1059), .B2(new_n1051), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n895), .A2(new_n896), .A3(G330), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1053), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT114), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n886), .B1(new_n830), .B2(new_n827), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n722), .A2(G330), .A3(new_n827), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n884), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1064), .B1(new_n1066), .B2(new_n1061), .ZN(new_n1067));
  AND3_X1   g0867(.A1(new_n1049), .A2(new_n887), .A3(new_n1048), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n895), .A2(KEYINPUT113), .A3(G330), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n827), .ZN(new_n1070));
  AOI21_X1  g0870(.A(KEYINPUT113), .B1(new_n895), .B2(G330), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n884), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1067), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n902), .A2(G330), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n837), .A2(new_n618), .A3(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1063), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n837), .A2(new_n618), .A3(new_n1074), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1049), .A2(new_n887), .A3(new_n1048), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1071), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1079), .A2(new_n827), .A3(new_n1069), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1078), .B1(new_n884), .B2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1077), .B(KEYINPUT114), .C1(new_n1081), .C2(new_n1067), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1062), .A2(new_n1076), .A3(new_n1082), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1083), .A2(new_n682), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1076), .A2(new_n1082), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1053), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n493), .A2(new_n604), .A3(new_n672), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(KEYINPUT97), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1088), .A2(new_n650), .A3(new_n697), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n665), .B1(new_n1089), .B2(new_n691), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n886), .B1(new_n1090), .B2(new_n827), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1051), .B1(new_n1091), .B2(new_n884), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1061), .B1(new_n1092), .B2(new_n1047), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1086), .A2(new_n1093), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n1085), .A2(KEYINPUT115), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(KEYINPUT115), .B1(new_n1085), .B2(new_n1094), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1084), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n866), .A2(new_n726), .A3(new_n876), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n800), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n761), .A2(new_n977), .B1(new_n748), .B2(new_n227), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n741), .A2(G150), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT53), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1100), .B(new_n1102), .C1(G125), .C2(new_n745), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n265), .B1(new_n757), .B2(new_n816), .ZN(new_n1104));
  INV_X1    g0904(.A(G128), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(KEYINPUT54), .B(G143), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n754), .A2(new_n1105), .B1(new_n762), .B2(new_n1106), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1104), .B(new_n1107), .C1(G159), .C2(new_n751), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n748), .A2(new_n321), .B1(new_n744), .B2(new_n804), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT116), .Z(new_n1110));
  OAI221_X1 g0910(.A(new_n326), .B1(new_n750), .B2(new_n204), .C1(new_n221), .C2(new_n740), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n761), .A2(new_n365), .B1(new_n762), .B2(new_n223), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n754), .A2(new_n747), .B1(new_n757), .B2(new_n507), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1103), .A2(new_n1108), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n737), .B1(new_n341), .B2(new_n1099), .C1(new_n1115), .C2(new_n781), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT117), .Z(new_n1117));
  AOI22_X1  g0917(.A1(new_n1094), .A2(new_n958), .B1(new_n1098), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1097), .A2(new_n1118), .ZN(G378));
  XOR2_X1   g0919(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1120));
  INV_X1    g0920(.A(KEYINPUT119), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n303), .B2(new_n309), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n308), .A2(new_n663), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n309), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n617), .A2(KEYINPUT119), .A3(new_n1124), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1122), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1123), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1120), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1123), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1122), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1120), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1128), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n726), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n737), .B1(G50), .B2(new_n1099), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n265), .A2(G41), .ZN(new_n1138));
  AOI211_X1 g0938(.A(G50), .B(new_n1138), .C1(new_n254), .C2(new_n255), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G107), .A2(new_n999), .B1(new_n745), .B2(G283), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n223), .B2(new_n761), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(G116), .A2(new_n808), .B1(new_n741), .B2(G77), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n968), .A2(G58), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1142), .A2(new_n974), .A3(new_n1138), .A4(new_n1143), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1141), .B(new_n1144), .C1(new_n556), .C2(new_n766), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1139), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(G125), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n754), .A2(new_n1148), .B1(new_n761), .B2(new_n816), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n766), .A2(G137), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1150), .B1(new_n1105), .B2(new_n757), .C1(new_n740), .C2(new_n1106), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1149), .B(new_n1151), .C1(G150), .C2(new_n751), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1153), .A2(KEYINPUT59), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n254), .B(new_n255), .C1(new_n748), .C2(new_n770), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G124), .B2(new_n745), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT59), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1156), .B1(new_n1152), .B2(new_n1157), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1147), .B1(new_n1146), .B2(new_n1145), .C1(new_n1154), .C2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1137), .B1(new_n1159), .B2(new_n780), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1136), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT120), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n900), .A2(KEYINPUT40), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n898), .A2(new_n895), .A3(new_n896), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n671), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1128), .A2(new_n1134), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1162), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1135), .B(KEYINPUT120), .C1(new_n901), .C2(new_n671), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1167), .A2(new_n1168), .B1(new_n1166), .B2(new_n1165), .ZN(new_n1169));
  OAI21_X1  g0969(.A(KEYINPUT121), .B1(new_n1169), .B2(new_n891), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1171), .A2(new_n891), .A3(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1170), .B(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n958), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1161), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT57), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1068), .A2(new_n1072), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1067), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(KEYINPUT114), .B1(new_n1180), .B2(new_n1077), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1073), .A2(new_n1063), .A3(new_n1075), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1094), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT115), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1085), .A2(KEYINPUT115), .A3(new_n1094), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1075), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1177), .B1(new_n1187), .B2(new_n1174), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1077), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n891), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT122), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1190), .B1(new_n1173), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1169), .A2(new_n891), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(KEYINPUT122), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1177), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n683), .B1(new_n1189), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1176), .B1(new_n1188), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(G375));
  NOR2_X1   g0998(.A1(new_n1180), .A2(new_n1077), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT123), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n942), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1200), .A2(new_n1201), .A3(new_n1076), .A4(new_n1082), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n736), .B1(new_n321), .B2(new_n800), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G97), .A2(new_n741), .B1(new_n745), .B2(G303), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n507), .B2(new_n761), .C1(new_n747), .C2(new_n757), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n754), .A2(new_n804), .B1(new_n762), .B2(new_n365), .ZN(new_n1206));
  NOR4_X1   g1006(.A1(new_n1205), .A2(new_n265), .A3(new_n976), .A4(new_n1206), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n770), .A2(new_n740), .B1(new_n761), .B2(new_n1106), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n762), .A2(new_n811), .B1(new_n744), .B2(new_n1105), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n754), .A2(new_n816), .B1(new_n757), .B2(new_n977), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1143), .A2(new_n265), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(G50), .C2(new_n751), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1207), .A2(new_n996), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1203), .B1(new_n781), .B2(new_n1214), .C1(new_n883), .C2(new_n727), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1073), .B2(new_n1175), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1202), .A2(new_n1217), .ZN(G381));
  NOR2_X1   g1018(.A1(G393), .A2(G396), .ZN(new_n1219));
  INV_X1    g1019(.A(G384), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT124), .ZN(new_n1222));
  INV_X1    g1022(.A(G390), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n959), .A2(new_n1223), .A3(new_n987), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1222), .A2(new_n1202), .A3(new_n1217), .A4(new_n1224), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1225), .A2(KEYINPUT125), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(G375), .A2(G378), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(KEYINPUT125), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .ZN(G407));
  NAND2_X1  g1029(.A1(new_n664), .A2(G213), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT126), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1227), .A2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(G407), .A2(G213), .A3(new_n1232), .ZN(G409));
  INV_X1    g1033(.A(KEYINPUT127), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1223), .B1(new_n959), .B2(new_n987), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(G393), .B(new_n798), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1224), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1236), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G387), .A2(G390), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n959), .A2(new_n1223), .A3(new_n987), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1238), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1234), .B1(new_n1237), .B2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1236), .B1(new_n1224), .B2(new_n1235), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1239), .A2(new_n1240), .A3(new_n1238), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n1244), .A3(KEYINPUT127), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1199), .A2(KEYINPUT60), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n682), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1076), .A2(new_n1082), .A3(KEYINPUT60), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1248), .B1(new_n1200), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1220), .B1(new_n1250), .B2(new_n1216), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT123), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1199), .B(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1249), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(G384), .B(new_n1217), .C1(new_n1255), .C2(new_n1248), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1231), .A2(G2897), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1251), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1257), .B1(new_n1251), .B2(new_n1256), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1170), .B(new_n1193), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1189), .A2(new_n1201), .A3(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1161), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1264), .B1(new_n1265), .B2(new_n958), .ZN(new_n1266));
  AOI21_X1  g1066(.A(G378), .B1(new_n1263), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(new_n1197), .B2(G378), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1261), .B1(new_n1268), .B2(new_n1231), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1264), .B1(new_n1262), .B2(new_n958), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n890), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1193), .B2(KEYINPUT122), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1173), .A2(new_n1191), .ZN(new_n1274));
  OAI21_X1  g1074(.A(KEYINPUT57), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n682), .B1(new_n1187), .B2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT57), .B1(new_n1189), .B2(new_n1262), .ZN(new_n1277));
  OAI211_X1 g1077(.A(G378), .B(new_n1270), .C1(new_n1276), .C2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1263), .A2(new_n1266), .ZN(new_n1279));
  INV_X1    g1079(.A(G378), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1278), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT62), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1231), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1251), .A2(new_n1256), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .A4(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT61), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1269), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  AOI211_X1 g1089(.A(new_n1231), .B(new_n1285), .C1(new_n1278), .C2(new_n1281), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1290), .A2(new_n1283), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1246), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1231), .B1(new_n1278), .B2(new_n1281), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1286), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1260), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1258), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1293), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT63), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1294), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1243), .A2(new_n1244), .A3(new_n1288), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1300), .B1(KEYINPUT63), .B2(new_n1290), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1292), .A2(new_n1302), .ZN(G405));
  OAI21_X1  g1103(.A(new_n1285), .B1(new_n1237), .B2(new_n1241), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1243), .A2(new_n1244), .A3(new_n1286), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1197), .A2(new_n1280), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1306), .B1(new_n1227), .B2(new_n1307), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1227), .A2(new_n1307), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1309), .A2(new_n1304), .A3(new_n1305), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1308), .A2(new_n1310), .ZN(G402));
endmodule


