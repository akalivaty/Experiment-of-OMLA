

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580;

  INV_X1 U321 ( .A(n560), .ZN(n499) );
  XNOR2_X1 U322 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U323 ( .A(n429), .B(n428), .Z(n289) );
  XOR2_X1 U324 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n290) );
  XOR2_X1 U325 ( .A(n434), .B(n433), .Z(n291) );
  NOR2_X1 U326 ( .A1(n500), .A2(n499), .ZN(n503) );
  XNOR2_X1 U327 ( .A(n435), .B(n291), .ZN(n436) );
  NOR2_X1 U328 ( .A1(n560), .A2(n559), .ZN(n562) );
  XNOR2_X1 U329 ( .A(n570), .B(KEYINPUT41), .ZN(n552) );
  XOR2_X1 U330 ( .A(KEYINPUT28), .B(n545), .Z(n513) );
  XOR2_X1 U331 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n293) );
  XNOR2_X1 U332 ( .A(KEYINPUT14), .B(KEYINPUT79), .ZN(n292) );
  XNOR2_X1 U333 ( .A(n293), .B(n292), .ZN(n306) );
  XOR2_X1 U334 ( .A(G57GAT), .B(KEYINPUT13), .Z(n295) );
  XNOR2_X1 U335 ( .A(G71GAT), .B(KEYINPUT71), .ZN(n294) );
  XNOR2_X1 U336 ( .A(n295), .B(n294), .ZN(n438) );
  XNOR2_X1 U337 ( .A(G8GAT), .B(G183GAT), .ZN(n296) );
  XNOR2_X1 U338 ( .A(n296), .B(G211GAT), .ZN(n362) );
  XOR2_X1 U339 ( .A(n362), .B(KEYINPUT12), .Z(n298) );
  NAND2_X1 U340 ( .A1(G231GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U342 ( .A(n438), .B(n299), .Z(n301) );
  XOR2_X1 U343 ( .A(G15GAT), .B(G127GAT), .Z(n337) );
  XOR2_X1 U344 ( .A(G22GAT), .B(G155GAT), .Z(n355) );
  XNOR2_X1 U345 ( .A(n337), .B(n355), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U347 ( .A(n302), .B(G64GAT), .Z(n304) );
  XOR2_X1 U348 ( .A(KEYINPUT68), .B(G1GAT), .Z(n410) );
  XNOR2_X1 U349 ( .A(n410), .B(G78GAT), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U351 ( .A(n306), .B(n305), .Z(n501) );
  XOR2_X1 U352 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n308) );
  XNOR2_X1 U353 ( .A(G43GAT), .B(G29GAT), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U355 ( .A(KEYINPUT67), .B(n309), .Z(n424) );
  XOR2_X1 U356 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n311) );
  XNOR2_X1 U357 ( .A(G134GAT), .B(G106GAT), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U359 ( .A(n424), .B(n312), .ZN(n321) );
  XOR2_X1 U360 ( .A(G85GAT), .B(KEYINPUT74), .Z(n314) );
  XNOR2_X1 U361 ( .A(G99GAT), .B(G92GAT), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n314), .B(n313), .ZN(n432) );
  XOR2_X1 U363 ( .A(G36GAT), .B(G190GAT), .Z(n366) );
  XOR2_X1 U364 ( .A(n432), .B(n366), .Z(n316) );
  NAND2_X1 U365 ( .A1(G232GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U367 ( .A(n317), .B(KEYINPUT9), .Z(n319) );
  XOR2_X1 U368 ( .A(G50GAT), .B(G162GAT), .Z(n354) );
  XNOR2_X1 U369 ( .A(G218GAT), .B(n354), .ZN(n318) );
  XNOR2_X1 U370 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n321), .B(n320), .ZN(n560) );
  NAND2_X1 U372 ( .A1(n501), .A2(n560), .ZN(n323) );
  XNOR2_X1 U373 ( .A(KEYINPUT81), .B(KEYINPUT16), .ZN(n322) );
  XNOR2_X1 U374 ( .A(n323), .B(n322), .ZN(n407) );
  XOR2_X1 U375 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n325) );
  XNOR2_X1 U376 ( .A(G71GAT), .B(G183GAT), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U378 ( .A(G176GAT), .B(G190GAT), .Z(n327) );
  XNOR2_X1 U379 ( .A(G43GAT), .B(G99GAT), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U381 ( .A(n329), .B(n328), .Z(n335) );
  XOR2_X1 U382 ( .A(G120GAT), .B(KEYINPUT0), .Z(n331) );
  XNOR2_X1 U383 ( .A(G113GAT), .B(G134GAT), .ZN(n330) );
  XNOR2_X1 U384 ( .A(n331), .B(n330), .ZN(n385) );
  XOR2_X1 U385 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n333) );
  XNOR2_X1 U386 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n370) );
  XNOR2_X1 U388 ( .A(n385), .B(n370), .ZN(n334) );
  XNOR2_X1 U389 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U390 ( .A(n337), .B(n336), .Z(n339) );
  NAND2_X1 U391 ( .A1(G227GAT), .A2(G233GAT), .ZN(n338) );
  XOR2_X1 U392 ( .A(n339), .B(n338), .Z(n510) );
  INV_X1 U393 ( .A(n510), .ZN(n547) );
  XOR2_X1 U394 ( .A(KEYINPUT86), .B(KEYINPUT2), .Z(n341) );
  XNOR2_X1 U395 ( .A(KEYINPUT3), .B(KEYINPUT85), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U397 ( .A(G141GAT), .B(n342), .Z(n389) );
  XOR2_X1 U398 ( .A(KEYINPUT83), .B(KEYINPUT87), .Z(n344) );
  XNOR2_X1 U399 ( .A(KEYINPUT24), .B(KEYINPUT88), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U401 ( .A(G211GAT), .B(KEYINPUT22), .Z(n346) );
  XNOR2_X1 U402 ( .A(KEYINPUT89), .B(KEYINPUT84), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U404 ( .A(n348), .B(n347), .Z(n360) );
  XOR2_X1 U405 ( .A(G204GAT), .B(KEYINPUT21), .Z(n350) );
  XNOR2_X1 U406 ( .A(G197GAT), .B(G218GAT), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n350), .B(n349), .ZN(n369) );
  XOR2_X1 U408 ( .A(n369), .B(KEYINPUT23), .Z(n352) );
  NAND2_X1 U409 ( .A1(G228GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n352), .B(n351), .ZN(n358) );
  XNOR2_X1 U411 ( .A(G106GAT), .B(G78GAT), .ZN(n353) );
  XNOR2_X1 U412 ( .A(n353), .B(G148GAT), .ZN(n439) );
  XNOR2_X1 U413 ( .A(n354), .B(n439), .ZN(n356) );
  XNOR2_X1 U414 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U416 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U417 ( .A(n389), .B(n361), .ZN(n545) );
  NOR2_X1 U418 ( .A1(n547), .A2(n513), .ZN(n395) );
  XOR2_X1 U419 ( .A(G176GAT), .B(G64GAT), .Z(n429) );
  XOR2_X1 U420 ( .A(n429), .B(KEYINPUT95), .Z(n364) );
  XNOR2_X1 U421 ( .A(n362), .B(G92GAT), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U423 ( .A(n366), .B(n365), .Z(n368) );
  NAND2_X1 U424 ( .A1(G226GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U425 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U426 ( .A(n370), .B(n369), .Z(n371) );
  XNOR2_X1 U427 ( .A(n372), .B(n371), .ZN(n539) );
  XNOR2_X1 U428 ( .A(KEYINPUT27), .B(n539), .ZN(n400) );
  XOR2_X1 U429 ( .A(G57GAT), .B(G155GAT), .Z(n374) );
  XNOR2_X1 U430 ( .A(G1GAT), .B(G148GAT), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U432 ( .A(G85GAT), .B(G162GAT), .Z(n376) );
  XNOR2_X1 U433 ( .A(G29GAT), .B(G127GAT), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U435 ( .A(n378), .B(n377), .ZN(n393) );
  XOR2_X1 U436 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n380) );
  XNOR2_X1 U437 ( .A(KEYINPUT4), .B(KEYINPUT94), .ZN(n379) );
  XNOR2_X1 U438 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U439 ( .A(KEYINPUT90), .B(KEYINPUT6), .Z(n382) );
  XNOR2_X1 U440 ( .A(KEYINPUT92), .B(KEYINPUT91), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U442 ( .A(n384), .B(n383), .Z(n391) );
  XOR2_X1 U443 ( .A(n385), .B(KEYINPUT1), .Z(n387) );
  NAND2_X1 U444 ( .A1(G225GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U446 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U448 ( .A(n393), .B(n392), .Z(n404) );
  INV_X1 U449 ( .A(n404), .ZN(n543) );
  NAND2_X1 U450 ( .A1(n400), .A2(n543), .ZN(n394) );
  XOR2_X1 U451 ( .A(KEYINPUT96), .B(n394), .Z(n509) );
  NAND2_X1 U452 ( .A1(n395), .A2(n509), .ZN(n406) );
  NAND2_X1 U453 ( .A1(n547), .A2(n539), .ZN(n396) );
  NAND2_X1 U454 ( .A1(n545), .A2(n396), .ZN(n397) );
  XOR2_X1 U455 ( .A(KEYINPUT25), .B(n397), .Z(n402) );
  NOR2_X1 U456 ( .A1(n547), .A2(n545), .ZN(n398) );
  XOR2_X1 U457 ( .A(KEYINPUT97), .B(n398), .Z(n399) );
  XOR2_X1 U458 ( .A(KEYINPUT26), .B(n399), .Z(n528) );
  INV_X1 U459 ( .A(n528), .ZN(n564) );
  NAND2_X1 U460 ( .A1(n400), .A2(n564), .ZN(n401) );
  NAND2_X1 U461 ( .A1(n402), .A2(n401), .ZN(n403) );
  NAND2_X1 U462 ( .A1(n404), .A2(n403), .ZN(n405) );
  NAND2_X1 U463 ( .A1(n406), .A2(n405), .ZN(n456) );
  NAND2_X1 U464 ( .A1(n407), .A2(n456), .ZN(n472) );
  XOR2_X1 U465 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n409) );
  XNOR2_X1 U466 ( .A(KEYINPUT69), .B(KEYINPUT29), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n409), .B(n408), .ZN(n414) );
  XOR2_X1 U468 ( .A(G50GAT), .B(G36GAT), .Z(n412) );
  XNOR2_X1 U469 ( .A(n410), .B(KEYINPUT66), .ZN(n411) );
  XNOR2_X1 U470 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U471 ( .A(n414), .B(n413), .Z(n416) );
  NAND2_X1 U472 ( .A1(G229GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U474 ( .A(G197GAT), .B(G15GAT), .Z(n418) );
  XNOR2_X1 U475 ( .A(G169GAT), .B(G113GAT), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U477 ( .A(n420), .B(n419), .Z(n426) );
  XOR2_X1 U478 ( .A(KEYINPUT70), .B(G8GAT), .Z(n422) );
  XNOR2_X1 U479 ( .A(G141GAT), .B(G22GAT), .ZN(n421) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U482 ( .A(n426), .B(n425), .Z(n470) );
  INV_X1 U483 ( .A(n470), .ZN(n566) );
  XNOR2_X1 U484 ( .A(G120GAT), .B(G204GAT), .ZN(n427) );
  XNOR2_X1 U485 ( .A(n290), .B(n427), .ZN(n428) );
  NAND2_X1 U486 ( .A1(G230GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n289), .B(n430), .ZN(n431) );
  XOR2_X1 U488 ( .A(n431), .B(KEYINPUT76), .Z(n437) );
  XNOR2_X1 U489 ( .A(n432), .B(KEYINPUT72), .ZN(n435) );
  XOR2_X1 U490 ( .A(KEYINPUT77), .B(KEYINPUT73), .Z(n434) );
  XNOR2_X1 U491 ( .A(KEYINPUT31), .B(KEYINPUT75), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n570) );
  NOR2_X1 U494 ( .A1(n566), .A2(n570), .ZN(n442) );
  XOR2_X1 U495 ( .A(KEYINPUT78), .B(n442), .Z(n460) );
  NOR2_X1 U496 ( .A1(n472), .A2(n460), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n443), .B(KEYINPUT98), .ZN(n452) );
  NAND2_X1 U498 ( .A1(n452), .A2(n543), .ZN(n447) );
  XOR2_X1 U499 ( .A(KEYINPUT100), .B(KEYINPUT34), .Z(n445) );
  XNOR2_X1 U500 ( .A(G1GAT), .B(KEYINPUT99), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(G1324GAT) );
  NAND2_X1 U503 ( .A1(n452), .A2(n539), .ZN(n448) );
  XNOR2_X1 U504 ( .A(n448), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U505 ( .A(KEYINPUT35), .B(KEYINPUT101), .Z(n450) );
  NAND2_X1 U506 ( .A1(n547), .A2(n452), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U508 ( .A(G15GAT), .B(n451), .Z(G1326GAT) );
  NAND2_X1 U509 ( .A1(n452), .A2(n513), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n453), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U511 ( .A(KEYINPUT102), .B(KEYINPUT105), .Z(n455) );
  XNOR2_X1 U512 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n454) );
  XNOR2_X1 U513 ( .A(n455), .B(n454), .ZN(n464) );
  XNOR2_X1 U514 ( .A(KEYINPUT36), .B(n560), .ZN(n577) );
  INV_X1 U515 ( .A(n501), .ZN(n574) );
  NAND2_X1 U516 ( .A1(n574), .A2(n456), .ZN(n457) );
  NOR2_X1 U517 ( .A1(n577), .A2(n457), .ZN(n458) );
  XOR2_X1 U518 ( .A(n458), .B(KEYINPUT37), .Z(n459) );
  XNOR2_X1 U519 ( .A(KEYINPUT103), .B(n459), .ZN(n482) );
  NOR2_X1 U520 ( .A1(n460), .A2(n482), .ZN(n462) );
  XNOR2_X1 U521 ( .A(KEYINPUT104), .B(KEYINPUT38), .ZN(n461) );
  XNOR2_X1 U522 ( .A(n462), .B(n461), .ZN(n468) );
  NAND2_X1 U523 ( .A1(n543), .A2(n468), .ZN(n463) );
  XOR2_X1 U524 ( .A(n464), .B(n463), .Z(G1328GAT) );
  NAND2_X1 U525 ( .A1(n539), .A2(n468), .ZN(n465) );
  XNOR2_X1 U526 ( .A(n465), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U527 ( .A1(n468), .A2(n547), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n466), .B(KEYINPUT40), .ZN(n467) );
  XNOR2_X1 U529 ( .A(G43GAT), .B(n467), .ZN(G1330GAT) );
  NAND2_X1 U530 ( .A1(n513), .A2(n468), .ZN(n469) );
  XNOR2_X1 U531 ( .A(n469), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U532 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n474) );
  NOR2_X1 U533 ( .A1(n470), .A2(n552), .ZN(n471) );
  XOR2_X1 U534 ( .A(KEYINPUT106), .B(n471), .Z(n483) );
  NOR2_X1 U535 ( .A1(n483), .A2(n472), .ZN(n477) );
  NAND2_X1 U536 ( .A1(n543), .A2(n477), .ZN(n473) );
  XNOR2_X1 U537 ( .A(n474), .B(n473), .ZN(G1332GAT) );
  NAND2_X1 U538 ( .A1(n539), .A2(n477), .ZN(n475) );
  XNOR2_X1 U539 ( .A(n475), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U540 ( .A1(n477), .A2(n547), .ZN(n476) );
  XNOR2_X1 U541 ( .A(n476), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n479) );
  NAND2_X1 U543 ( .A1(n477), .A2(n513), .ZN(n478) );
  XNOR2_X1 U544 ( .A(n479), .B(n478), .ZN(n481) );
  XOR2_X1 U545 ( .A(G78GAT), .B(KEYINPUT108), .Z(n480) );
  XNOR2_X1 U546 ( .A(n481), .B(n480), .ZN(G1335GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n485) );
  NOR2_X1 U548 ( .A1(n483), .A2(n482), .ZN(n491) );
  NAND2_X1 U549 ( .A1(n491), .A2(n543), .ZN(n484) );
  XNOR2_X1 U550 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U551 ( .A(G85GAT), .B(n486), .ZN(G1336GAT) );
  XOR2_X1 U552 ( .A(G92GAT), .B(KEYINPUT111), .Z(n488) );
  NAND2_X1 U553 ( .A1(n491), .A2(n539), .ZN(n487) );
  XNOR2_X1 U554 ( .A(n488), .B(n487), .ZN(G1337GAT) );
  NAND2_X1 U555 ( .A1(n491), .A2(n547), .ZN(n489) );
  XNOR2_X1 U556 ( .A(n489), .B(KEYINPUT112), .ZN(n490) );
  XNOR2_X1 U557 ( .A(G99GAT), .B(n490), .ZN(G1338GAT) );
  NAND2_X1 U558 ( .A1(n513), .A2(n491), .ZN(n492) );
  XNOR2_X1 U559 ( .A(n492), .B(KEYINPUT44), .ZN(n493) );
  XNOR2_X1 U560 ( .A(G106GAT), .B(n493), .ZN(G1339GAT) );
  XNOR2_X1 U561 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n495) );
  NOR2_X1 U562 ( .A1(n574), .A2(n577), .ZN(n494) );
  XOR2_X1 U563 ( .A(n495), .B(n494), .Z(n496) );
  NOR2_X1 U564 ( .A1(n570), .A2(n496), .ZN(n497) );
  NAND2_X1 U565 ( .A1(n497), .A2(n566), .ZN(n507) );
  XOR2_X1 U566 ( .A(KEYINPUT47), .B(KEYINPUT114), .Z(n505) );
  NOR2_X1 U567 ( .A1(n566), .A2(n552), .ZN(n498) );
  XNOR2_X1 U568 ( .A(n498), .B(KEYINPUT46), .ZN(n500) );
  XOR2_X1 U569 ( .A(KEYINPUT113), .B(n501), .Z(n555) );
  INV_X1 U570 ( .A(n555), .ZN(n502) );
  NAND2_X1 U571 ( .A1(n503), .A2(n502), .ZN(n504) );
  XNOR2_X1 U572 ( .A(n505), .B(n504), .ZN(n506) );
  NAND2_X1 U573 ( .A1(n507), .A2(n506), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n508), .B(KEYINPUT48), .ZN(n540) );
  NAND2_X1 U575 ( .A1(n540), .A2(n509), .ZN(n527) );
  NOR2_X1 U576 ( .A1(n510), .A2(n527), .ZN(n511) );
  XNOR2_X1 U577 ( .A(KEYINPUT115), .B(n511), .ZN(n512) );
  NOR2_X1 U578 ( .A1(n513), .A2(n512), .ZN(n519) );
  INV_X1 U579 ( .A(n519), .ZN(n523) );
  NOR2_X1 U580 ( .A1(n566), .A2(n523), .ZN(n514) );
  XOR2_X1 U581 ( .A(G113GAT), .B(n514), .Z(G1340GAT) );
  NOR2_X1 U582 ( .A1(n523), .A2(n552), .ZN(n518) );
  XOR2_X1 U583 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n516) );
  XNOR2_X1 U584 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n515) );
  XNOR2_X1 U585 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U586 ( .A(n518), .B(n517), .ZN(G1341GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n521) );
  NAND2_X1 U588 ( .A1(n519), .A2(n555), .ZN(n520) );
  XNOR2_X1 U589 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U590 ( .A(G127GAT), .B(n522), .Z(G1342GAT) );
  NOR2_X1 U591 ( .A1(n560), .A2(n523), .ZN(n525) );
  XNOR2_X1 U592 ( .A(KEYINPUT119), .B(KEYINPUT51), .ZN(n524) );
  XNOR2_X1 U593 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U594 ( .A(G134GAT), .B(n526), .Z(G1343GAT) );
  NOR2_X1 U595 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U596 ( .A(KEYINPUT120), .B(n529), .Z(n537) );
  NOR2_X1 U597 ( .A1(n566), .A2(n537), .ZN(n530) );
  XOR2_X1 U598 ( .A(G141GAT), .B(n530), .Z(G1344GAT) );
  NOR2_X1 U599 ( .A1(n552), .A2(n537), .ZN(n534) );
  XOR2_X1 U600 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n532) );
  XNOR2_X1 U601 ( .A(G148GAT), .B(KEYINPUT121), .ZN(n531) );
  XNOR2_X1 U602 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U603 ( .A(n534), .B(n533), .ZN(G1345GAT) );
  NOR2_X1 U604 ( .A1(n537), .A2(n574), .ZN(n535) );
  XOR2_X1 U605 ( .A(KEYINPUT122), .B(n535), .Z(n536) );
  XNOR2_X1 U606 ( .A(G155GAT), .B(n536), .ZN(G1346GAT) );
  NOR2_X1 U607 ( .A1(n560), .A2(n537), .ZN(n538) );
  XOR2_X1 U608 ( .A(G162GAT), .B(n538), .Z(G1347GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT123), .B(KEYINPUT54), .Z(n542) );
  NAND2_X1 U610 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U611 ( .A(n542), .B(n541), .ZN(n544) );
  NOR2_X2 U612 ( .A1(n544), .A2(n543), .ZN(n565) );
  NAND2_X1 U613 ( .A1(n565), .A2(n545), .ZN(n546) );
  XNOR2_X1 U614 ( .A(KEYINPUT55), .B(n546), .ZN(n548) );
  NAND2_X1 U615 ( .A1(n548), .A2(n547), .ZN(n559) );
  NOR2_X1 U616 ( .A1(n566), .A2(n559), .ZN(n549) );
  XOR2_X1 U617 ( .A(G169GAT), .B(n549), .Z(G1348GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT56), .B(KEYINPUT124), .Z(n551) );
  XNOR2_X1 U619 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n550) );
  XNOR2_X1 U620 ( .A(n551), .B(n550), .ZN(n554) );
  NOR2_X1 U621 ( .A1(n552), .A2(n559), .ZN(n553) );
  XOR2_X1 U622 ( .A(n554), .B(n553), .Z(G1349GAT) );
  XOR2_X1 U623 ( .A(G183GAT), .B(KEYINPUT125), .Z(n558) );
  INV_X1 U624 ( .A(n559), .ZN(n556) );
  NAND2_X1 U625 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(G1350GAT) );
  XNOR2_X1 U627 ( .A(KEYINPUT126), .B(KEYINPUT58), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n563) );
  XOR2_X1 U629 ( .A(G190GAT), .B(n563), .Z(G1351GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n576) );
  NOR2_X1 U631 ( .A1(n566), .A2(n576), .ZN(n568) );
  XNOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .Z(n573) );
  INV_X1 U636 ( .A(n576), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n576), .ZN(n575) );
  XOR2_X1 U640 ( .A(G211GAT), .B(n575), .Z(G1354GAT) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n579) );
  XNOR2_X1 U642 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

