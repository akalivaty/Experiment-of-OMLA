//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n830, new_n832, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(KEYINPUT41), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT97), .ZN(new_n205));
  XNOR2_X1  g004(.A(G134gat), .B(G162gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT14), .B(G29gat), .ZN(new_n210));
  INV_X1    g009(.A(G36gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G29gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT88), .ZN(new_n216));
  XNOR2_X1  g015(.A(G43gat), .B(G50gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT15), .ZN(new_n218));
  OR3_X1    g017(.A1(new_n215), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n216), .B1(new_n215), .B2(new_n218), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(new_n217), .B(KEYINPUT15), .Z(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(new_n215), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT17), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT89), .ZN(new_n227));
  AOI22_X1  g026(.A1(new_n219), .A2(new_n220), .B1(new_n215), .B2(new_n222), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n227), .B1(new_n228), .B2(KEYINPUT17), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n224), .A2(KEYINPUT89), .A3(new_n225), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n226), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(KEYINPUT99), .A2(G85gat), .A3(G92gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n232), .B(KEYINPUT7), .ZN(new_n233));
  NAND2_X1  g032(.A1(G99gat), .A2(G106gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT8), .ZN(new_n235));
  XOR2_X1   g034(.A(KEYINPUT100), .B(G92gat), .Z(new_n236));
  OAI211_X1 g035(.A(new_n233), .B(new_n235), .C1(G85gat), .C2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G99gat), .B(G106gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n231), .A2(new_n240), .ZN(new_n241));
  AOI22_X1  g040(.A1(new_n224), .A2(new_n239), .B1(KEYINPUT41), .B2(new_n203), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT101), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT101), .ZN(new_n244));
  INV_X1    g043(.A(new_n242), .ZN(new_n245));
  AOI211_X1 g044(.A(new_n244), .B(new_n245), .C1(new_n231), .C2(new_n240), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n209), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n229), .ZN(new_n248));
  INV_X1    g047(.A(new_n226), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n248), .A2(new_n249), .A3(new_n240), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n244), .B1(new_n250), .B2(new_n245), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n241), .A2(KEYINPUT101), .A3(new_n242), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(G190gat), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n247), .A2(new_n253), .A3(G218gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT98), .ZN(new_n255));
  AOI21_X1  g054(.A(G218gat), .B1(new_n247), .B2(new_n253), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n208), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n256), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n258), .A2(KEYINPUT98), .A3(new_n254), .A4(new_n207), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT94), .B(G57gat), .Z(new_n261));
  INV_X1    g060(.A(KEYINPUT95), .ZN(new_n262));
  INV_X1    g061(.A(G64gat), .ZN(new_n263));
  OR3_X1    g062(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n262), .B1(new_n261), .B2(new_n263), .ZN(new_n265));
  INV_X1    g064(.A(G57gat), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT96), .B1(new_n266), .B2(G64gat), .ZN(new_n267));
  OR3_X1    g066(.A1(new_n266), .A2(KEYINPUT96), .A3(G64gat), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n264), .A2(new_n265), .A3(new_n267), .A4(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n270), .B(KEYINPUT93), .Z(new_n271));
  XOR2_X1   g070(.A(G71gat), .B(G78gat), .Z(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  XOR2_X1   g074(.A(G57gat), .B(G64gat), .Z(new_n276));
  NAND2_X1  g075(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(new_n272), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT21), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G231gat), .A2(G233gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(G127gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(G15gat), .B(G22gat), .ZN(new_n285));
  OR2_X1    g084(.A1(new_n285), .A2(G1gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT90), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT16), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n285), .B1(new_n288), .B2(G1gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n286), .A2(KEYINPUT90), .ZN(new_n291));
  OAI21_X1  g090(.A(G8gat), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT91), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G8gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n289), .A2(new_n293), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n294), .A2(new_n295), .A3(new_n286), .A4(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(new_n279), .B2(new_n280), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n284), .B(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n301), .B(G155gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(G183gat), .B(G211gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n300), .B(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n260), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G230gat), .A2(G233gat), .ZN(new_n308));
  XOR2_X1   g107(.A(new_n308), .B(KEYINPUT103), .Z(new_n309));
  INV_X1    g108(.A(KEYINPUT102), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n238), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n275), .A2(new_n278), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n240), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT10), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n239), .A2(new_n278), .A3(new_n275), .A4(new_n311), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n239), .A2(KEYINPUT10), .A3(new_n275), .A4(new_n278), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n309), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  XOR2_X1   g118(.A(G120gat), .B(G148gat), .Z(new_n320));
  XNOR2_X1  g119(.A(new_n320), .B(KEYINPUT104), .ZN(new_n321));
  XNOR2_X1  g120(.A(G176gat), .B(G204gat), .ZN(new_n322));
  XOR2_X1   g121(.A(new_n321), .B(new_n322), .Z(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n309), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n313), .A2(new_n315), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n319), .B(new_n324), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n325), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n323), .B1(new_n328), .B2(new_n318), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(KEYINPUT105), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT105), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n331), .B(new_n323), .C1(new_n328), .C2(new_n318), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n307), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n248), .A2(new_n298), .A3(new_n249), .ZN(new_n335));
  NAND2_X1  g134(.A1(G229gat), .A2(G233gat), .ZN(new_n336));
  OR2_X1    g135(.A1(new_n298), .A2(new_n228), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT18), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n336), .B(KEYINPUT13), .Z(new_n340));
  NAND2_X1  g139(.A1(new_n298), .A2(new_n228), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT92), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n298), .A2(KEYINPUT92), .A3(new_n228), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(new_n337), .A3(new_n344), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n338), .A2(new_n339), .B1(new_n340), .B2(new_n345), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n335), .A2(new_n337), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(KEYINPUT18), .A3(new_n336), .ZN(new_n348));
  XNOR2_X1  g147(.A(G113gat), .B(G141gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(G169gat), .B(G197gat), .Z(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT12), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n346), .A2(new_n348), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n354), .B1(new_n346), .B2(new_n348), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT78), .B(KEYINPUT5), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362));
  OR2_X1    g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n362), .B1(new_n363), .B2(KEYINPUT2), .ZN(new_n364));
  INV_X1    g163(.A(G141gat), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT77), .B1(new_n365), .B2(G148gat), .ZN(new_n366));
  INV_X1    g165(.A(G148gat), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n366), .B1(G141gat), .B2(new_n367), .ZN(new_n368));
  NOR3_X1   g167(.A1(new_n365), .A2(KEYINPUT77), .A3(G148gat), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n364), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G141gat), .B(G148gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT76), .B(KEYINPUT2), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n362), .B(new_n363), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT3), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n370), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n374), .B1(new_n370), .B2(new_n373), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  XOR2_X1   g176(.A(G127gat), .B(G134gat), .Z(new_n378));
  NOR2_X1   g177(.A1(G113gat), .A2(G120gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G113gat), .A2(G120gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NOR3_X1   g181(.A1(new_n378), .A2(new_n382), .A3(KEYINPUT1), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT69), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n380), .A2(new_n385), .A3(new_n381), .ZN(new_n386));
  AND2_X1   g185(.A1(G113gat), .A2(G120gat), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT69), .B1(new_n387), .B2(new_n379), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT1), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT70), .ZN(new_n391));
  NOR2_X1   g190(.A1(G127gat), .A2(G134gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(KEYINPUT68), .B(G127gat), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n392), .B1(new_n393), .B2(G134gat), .ZN(new_n394));
  AND3_X1   g193(.A1(new_n390), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n391), .B1(new_n390), .B2(new_n394), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n384), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI211_X1 g196(.A(new_n359), .B(new_n361), .C1(new_n377), .C2(new_n397), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n370), .A2(new_n373), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n399), .B(new_n384), .C1(new_n395), .C2(new_n396), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT4), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n390), .A2(new_n394), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT70), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n390), .A2(new_n391), .A3(new_n394), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT4), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n405), .A2(new_n406), .A3(new_n384), .A4(new_n399), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT80), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n401), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n383), .B1(new_n403), .B2(new_n404), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n410), .A2(KEYINPUT80), .A3(new_n406), .A4(new_n399), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n398), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT81), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n398), .A2(new_n409), .A3(KEYINPUT81), .A4(new_n411), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n399), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n397), .A2(new_n417), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n418), .A2(new_n400), .ZN(new_n419));
  OAI211_X1 g218(.A(KEYINPUT79), .B(new_n359), .C1(new_n419), .C2(new_n360), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT79), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n360), .B1(new_n418), .B2(new_n400), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(new_n358), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n377), .A2(new_n397), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n360), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n401), .A2(new_n407), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n420), .B(new_n423), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n416), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G1gat), .B(G29gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT0), .ZN(new_n430));
  XNOR2_X1  g229(.A(G57gat), .B(G85gat), .ZN(new_n431));
  XOR2_X1   g230(.A(new_n430), .B(new_n431), .Z(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT6), .ZN(new_n433));
  INV_X1    g232(.A(new_n432), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n428), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n416), .A2(new_n427), .A3(new_n435), .A4(new_n434), .ZN(new_n438));
  NAND2_X1  g237(.A1(G226gat), .A2(G233gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(G169gat), .A2(G176gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT64), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT64), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(G169gat), .A3(G176gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n445));
  OR3_X1    g244(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(G183gat), .A2(G190gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OR2_X1    g248(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(KEYINPUT27), .B(G183gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT28), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n452), .A2(KEYINPUT28), .A3(new_n453), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n449), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT24), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n448), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n461));
  INV_X1    g260(.A(G183gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n209), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT23), .ZN(new_n465));
  INV_X1    g264(.A(G169gat), .ZN(new_n466));
  INV_X1    g265(.A(G176gat), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n464), .A2(new_n470), .A3(new_n444), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT25), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(new_n444), .A3(KEYINPUT25), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n450), .A2(new_n462), .A3(new_n451), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT66), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT66), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n476), .A2(new_n478), .A3(new_n461), .A4(new_n480), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n473), .A2(KEYINPUT65), .B1(new_n475), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT65), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n471), .A2(new_n483), .A3(new_n472), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n458), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n439), .B1(new_n485), .B2(KEYINPUT29), .ZN(new_n486));
  XNOR2_X1  g285(.A(G197gat), .B(G204gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT74), .B(G211gat), .ZN(new_n488));
  INV_X1    g287(.A(G218gat), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(KEYINPUT73), .B(KEYINPUT22), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G211gat), .B(G218gat), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n493), .B(new_n487), .C1(new_n490), .C2(new_n491), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n473), .A2(KEYINPUT65), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n475), .A2(new_n481), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n484), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n456), .A2(new_n457), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n501), .A2(new_n448), .A3(new_n447), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n439), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n486), .A2(new_n497), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT29), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n504), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT75), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n509), .B1(new_n485), .B2(new_n439), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n503), .A2(KEYINPUT75), .A3(new_n504), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n508), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n506), .B1(new_n512), .B2(new_n497), .ZN(new_n513));
  XNOR2_X1  g312(.A(G8gat), .B(G36gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(G64gat), .B(G92gat), .ZN(new_n515));
  XOR2_X1   g314(.A(new_n514), .B(new_n515), .Z(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  OR3_X1    g316(.A1(new_n513), .A2(KEYINPUT30), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n510), .A2(new_n511), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n497), .B1(new_n519), .B2(new_n486), .ZN(new_n520));
  INV_X1    g319(.A(new_n506), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n506), .B(new_n516), .C1(new_n512), .C2(new_n497), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(KEYINPUT30), .A3(new_n523), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n437), .A2(new_n438), .B1(new_n518), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n497), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(KEYINPUT29), .B2(new_n375), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n527), .A2(KEYINPUT83), .B1(G228gat), .B2(G233gat), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT83), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n526), .B(new_n529), .C1(KEYINPUT29), .C2(new_n375), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n495), .A2(KEYINPUT82), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT82), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n532), .B1(new_n492), .B2(new_n494), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n496), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT3), .B1(new_n534), .B2(new_n507), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n528), .B(new_n530), .C1(new_n535), .C2(new_n399), .ZN(new_n536));
  INV_X1    g335(.A(new_n527), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n497), .A2(new_n507), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n399), .B1(new_n538), .B2(new_n374), .ZN(new_n539));
  OAI211_X1 g338(.A(G228gat), .B(G233gat), .C1(new_n537), .C2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT31), .B(G50gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G78gat), .B(G106gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(G22gat), .ZN(new_n545));
  INV_X1    g344(.A(new_n542), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n535), .A2(new_n399), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n527), .A2(KEYINPUT83), .ZN(new_n548));
  NAND2_X1  g347(.A1(G228gat), .A2(G233gat), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(new_n530), .A3(new_n549), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n540), .B(new_n546), .C1(new_n547), .C2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n543), .A2(new_n545), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n545), .ZN(new_n553));
  INV_X1    g352(.A(new_n551), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n546), .B1(new_n536), .B2(new_n540), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n525), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n484), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n476), .A2(new_n461), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n479), .B(new_n477), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n474), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n483), .B1(new_n471), .B2(new_n472), .ZN(new_n563));
  NOR3_X1   g362(.A1(new_n559), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n410), .B1(new_n564), .B2(new_n458), .ZN(new_n565));
  INV_X1    g364(.A(G227gat), .ZN(new_n566));
  INV_X1    g365(.A(G233gat), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n397), .A2(new_n500), .A3(new_n502), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n565), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT32), .ZN(new_n571));
  XNOR2_X1  g370(.A(G15gat), .B(G43gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(G71gat), .B(G99gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n571), .B1(KEYINPUT33), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT72), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n571), .A2(new_n575), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT71), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT33), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n580), .B1(new_n570), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n570), .A2(new_n580), .A3(new_n581), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n578), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n581), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT71), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n574), .B1(new_n570), .B2(KEYINPUT32), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n587), .A2(new_n578), .A3(new_n584), .A4(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n577), .B1(new_n585), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n565), .A2(new_n569), .ZN(new_n592));
  INV_X1    g391(.A(new_n568), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT34), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n587), .A2(new_n584), .A3(new_n588), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT72), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(new_n589), .ZN(new_n599));
  INV_X1    g398(.A(new_n595), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n600), .A3(new_n577), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n596), .A2(KEYINPUT36), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT36), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n600), .B1(new_n599), .B2(new_n577), .ZN(new_n604));
  AOI211_X1 g403(.A(new_n595), .B(new_n576), .C1(new_n598), .C2(new_n589), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n558), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n552), .A2(new_n556), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT38), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n517), .A2(KEYINPUT37), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n522), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n513), .A2(KEYINPUT37), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n517), .B1(new_n513), .B2(KEYINPUT37), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n512), .A2(new_n526), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n486), .A2(new_n526), .A3(new_n505), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT37), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n609), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n523), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n437), .A2(new_n438), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n608), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n428), .A2(new_n434), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n623), .A2(new_n518), .A3(new_n524), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n409), .A2(new_n411), .A3(new_n424), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n361), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n627), .B1(new_n419), .B2(new_n360), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n625), .A2(new_n627), .A3(new_n361), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n630), .A2(KEYINPUT84), .A3(new_n432), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT84), .B1(new_n630), .B2(new_n432), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT40), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n634), .B1(new_n626), .B2(new_n628), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n636), .B1(new_n631), .B2(new_n632), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n624), .A2(KEYINPUT85), .A3(new_n635), .A4(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT85), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n637), .A2(new_n518), .A3(new_n623), .A4(new_n524), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n630), .A2(new_n432), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT84), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n630), .A2(KEYINPUT84), .A3(new_n432), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT40), .B1(new_n645), .B2(new_n629), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n639), .B1(new_n640), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n622), .A2(new_n638), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n607), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n596), .A2(new_n557), .A3(new_n525), .A4(new_n601), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT86), .B(KEYINPUT35), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n604), .A2(new_n605), .ZN(new_n653));
  NAND2_X1  g452(.A1(KEYINPUT86), .A2(KEYINPUT35), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n653), .A2(new_n557), .A3(new_n525), .A4(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n357), .B1(new_n649), .B2(new_n656), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n334), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n621), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g459(.A1(new_n518), .A2(new_n524), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT16), .B(G8gat), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT42), .Z(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(G8gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT106), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(G1325gat));
  INV_X1    g468(.A(new_n658), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n602), .A2(new_n606), .ZN(new_n671));
  OAI21_X1  g470(.A(G15gat), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n653), .ZN(new_n673));
  OR2_X1    g472(.A1(new_n673), .A2(G15gat), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n672), .B1(new_n670), .B2(new_n674), .ZN(G1326gat));
  NAND3_X1  g474(.A1(new_n334), .A2(new_n657), .A3(new_n608), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT107), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT43), .B(G22gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  NOR2_X1   g478(.A1(new_n306), .A2(new_n333), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(new_n357), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n260), .B1(new_n649), .B2(new_n656), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n621), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n684), .A2(G29gat), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT45), .Z(new_n687));
  INV_X1    g486(.A(KEYINPUT108), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n649), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n607), .A2(new_n648), .A3(KEYINPUT108), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n652), .A2(KEYINPUT109), .A3(new_n655), .ZN(new_n692));
  AOI21_X1  g491(.A(KEYINPUT109), .B1(new_n652), .B2(new_n655), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  AND2_X1   g494(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n257), .A2(new_n259), .ZN(new_n697));
  NOR2_X1   g496(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700));
  OAI22_X1  g499(.A1(new_n695), .A2(new_n699), .B1(new_n700), .B2(new_n683), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n682), .ZN(new_n702));
  OAI21_X1  g501(.A(G29gat), .B1(new_n702), .B2(new_n685), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n703), .ZN(G1328gat));
  NOR3_X1   g503(.A1(new_n684), .A2(G36gat), .A3(new_n661), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT46), .ZN(new_n706));
  OAI21_X1  g505(.A(G36gat), .B1(new_n702), .B2(new_n661), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(G1329gat));
  INV_X1    g507(.A(new_n671), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G43gat), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n684), .A2(new_n673), .ZN(new_n711));
  OAI22_X1  g510(.A1(new_n702), .A2(new_n710), .B1(G43gat), .B2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g512(.A1(new_n657), .A2(new_n608), .ZN(new_n714));
  NOR4_X1   g513(.A1(new_n714), .A2(G50gat), .A3(new_n260), .A4(new_n681), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n701), .A2(new_n608), .A3(new_n682), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n715), .B1(new_n716), .B2(G50gat), .ZN(new_n717));
  XNOR2_X1  g516(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n717), .B(new_n719), .ZN(G1331gat));
  OR2_X1    g519(.A1(new_n355), .A2(new_n356), .ZN(new_n721));
  INV_X1    g520(.A(new_n333), .ZN(new_n722));
  NOR4_X1   g521(.A1(new_n695), .A2(new_n721), .A3(new_n307), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n621), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(new_n261), .ZN(G1332gat));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n662), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n727));
  XOR2_X1   g526(.A(KEYINPUT49), .B(G64gat), .Z(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n726), .B2(new_n728), .ZN(G1333gat));
  INV_X1    g528(.A(G71gat), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n723), .A2(new_n730), .A3(new_n653), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n730), .B1(new_n723), .B2(new_n709), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT50), .ZN(new_n733));
  OR3_X1    g532(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n731), .B2(new_n732), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(G1334gat));
  NAND2_X1  g535(.A1(new_n723), .A2(new_n608), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g537(.A1(new_n722), .A2(new_n685), .A3(G85gat), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT114), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n607), .A2(KEYINPUT108), .A3(new_n648), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT108), .B1(new_n607), .B2(new_n648), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n656), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n652), .A2(new_n655), .A3(KEYINPUT109), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n305), .A2(new_n357), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n260), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n748), .A2(KEYINPUT51), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT51), .B1(new_n748), .B2(new_n750), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n752), .A2(new_n753), .A3(KEYINPUT113), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT113), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n750), .B1(new_n691), .B2(new_n694), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n755), .B1(new_n758), .B2(new_n751), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n740), .B1(new_n754), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n749), .A2(new_n722), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT112), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n701), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(G85gat), .B1(new_n763), .B2(new_n685), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n760), .A2(new_n764), .ZN(G1336gat));
  NOR2_X1   g564(.A1(new_n661), .A2(G92gat), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  AOI211_X1 g566(.A(new_n722), .B(new_n767), .C1(new_n758), .C2(new_n751), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n699), .B1(new_n743), .B2(new_n747), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n683), .A2(new_n700), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n662), .B(new_n762), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n236), .ZN(new_n773));
  XNOR2_X1  g572(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n769), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n772), .A2(new_n776), .A3(new_n236), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n772), .B2(new_n236), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n777), .A2(new_n768), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n775), .B1(new_n779), .B2(new_n780), .ZN(G1337gat));
  NOR3_X1   g580(.A1(new_n673), .A2(new_n722), .A3(G99gat), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n782), .B1(new_n754), .B2(new_n759), .ZN(new_n783));
  OAI21_X1  g582(.A(G99gat), .B1(new_n763), .B2(new_n671), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1338gat));
  NAND3_X1  g584(.A1(new_n701), .A2(new_n608), .A3(new_n762), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G106gat), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n557), .A2(G106gat), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n333), .B(new_n788), .C1(new_n752), .C2(new_n753), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n787), .A2(KEYINPUT117), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT53), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n787), .A2(new_n789), .A3(KEYINPUT117), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(G1339gat));
  NOR4_X1   g593(.A1(new_n697), .A2(new_n305), .A3(new_n721), .A4(new_n333), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n316), .A2(new_n309), .A3(new_n317), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n319), .A2(KEYINPUT54), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n324), .B1(new_n318), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n797), .A2(KEYINPUT55), .A3(new_n799), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n802), .A2(new_n327), .A3(new_n803), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n357), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n347), .A2(new_n336), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n345), .A2(new_n340), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n353), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n346), .A2(new_n348), .A3(new_n354), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n808), .A2(new_n809), .A3(new_n330), .A4(new_n332), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n810), .A2(KEYINPUT118), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(KEYINPUT118), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n805), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n260), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n808), .A2(new_n809), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n803), .A2(new_n327), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(new_n802), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n697), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n795), .B1(new_n820), .B2(new_n305), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n653), .A2(new_n557), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n685), .A2(new_n662), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n721), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n333), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g628(.A1(new_n825), .A2(new_n306), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(new_n393), .ZN(G1342gat));
  INV_X1    g630(.A(KEYINPUT56), .ZN(new_n832));
  INV_X1    g631(.A(G134gat), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n825), .B(new_n697), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n834), .B(new_n835), .ZN(G1343gat));
  NOR2_X1   g635(.A1(new_n709), .A2(new_n824), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(new_n821), .B2(new_n557), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n557), .A2(new_n839), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n810), .B1(new_n357), .B2(new_n804), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(new_n257), .A3(new_n259), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n306), .B1(new_n819), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n841), .B1(new_n844), .B2(new_n795), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n838), .B1(new_n840), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(G141gat), .A3(new_n721), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT58), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n848), .A2(KEYINPUT119), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n709), .A2(new_n557), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n823), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n821), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n721), .ZN(new_n853));
  AOI22_X1  g652(.A1(new_n853), .A2(new_n365), .B1(KEYINPUT119), .B2(new_n848), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n847), .A2(new_n849), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n849), .B1(new_n847), .B2(new_n854), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(G1344gat));
  NAND2_X1  g656(.A1(new_n852), .A2(new_n333), .ZN(new_n858));
  AOI21_X1  g657(.A(G148gat), .B1(new_n858), .B2(KEYINPUT59), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n722), .A2(KEYINPUT59), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n859), .B1(new_n846), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n843), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n817), .B1(new_n257), .B2(new_n259), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT120), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n819), .A2(new_n865), .A3(new_n843), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n305), .A3(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n260), .A2(new_n357), .A3(new_n306), .A4(new_n722), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n557), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n841), .ZN(new_n870));
  OAI22_X1  g669(.A1(new_n869), .A2(KEYINPUT57), .B1(new_n821), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n333), .A3(new_n837), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n861), .A2(new_n873), .ZN(G1345gat));
  INV_X1    g673(.A(G155gat), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n852), .A2(new_n875), .A3(new_n306), .ZN(new_n876));
  AOI211_X1 g675(.A(new_n305), .B(new_n838), .C1(new_n840), .C2(new_n845), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(new_n875), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT121), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n880), .B(new_n876), .C1(new_n877), .C2(new_n875), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(G1346gat));
  AOI21_X1  g681(.A(G162gat), .B1(new_n852), .B2(new_n697), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n697), .A2(G162gat), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n883), .B1(new_n846), .B2(new_n884), .ZN(G1347gat));
  AOI21_X1  g684(.A(new_n863), .B1(new_n813), .B2(new_n260), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n868), .B1(new_n886), .B2(new_n306), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n822), .A2(new_n661), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n887), .A2(new_n685), .A3(new_n888), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n889), .A2(new_n466), .A3(new_n357), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n891), .B1(new_n821), .B2(new_n621), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n887), .A2(KEYINPUT122), .A3(new_n685), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n721), .A3(new_n888), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n890), .B1(new_n895), .B2(new_n466), .ZN(G1348gat));
  OAI21_X1  g695(.A(G176gat), .B1(new_n889), .B2(new_n722), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n894), .A2(new_n888), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n333), .A2(new_n467), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(G1349gat));
  OR3_X1    g699(.A1(new_n889), .A2(KEYINPUT123), .A3(new_n305), .ZN(new_n901));
  OAI21_X1  g700(.A(KEYINPUT123), .B1(new_n889), .B2(new_n305), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n901), .A2(G183gat), .A3(new_n902), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n894), .A2(new_n453), .A3(new_n306), .A4(new_n888), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g704(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1350gat));
  OAI21_X1  g709(.A(G190gat), .B1(new_n889), .B2(new_n260), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT61), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n697), .A2(new_n452), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n898), .B2(new_n913), .ZN(G1351gat));
  NAND2_X1  g713(.A1(new_n850), .A2(new_n662), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n894), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(KEYINPUT125), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n915), .B1(new_n892), .B2(new_n893), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT125), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n918), .A2(new_n721), .A3(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(G197gat), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n709), .A2(new_n621), .A3(new_n661), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n871), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n357), .A2(new_n923), .ZN(new_n926));
  AOI22_X1  g725(.A1(new_n922), .A2(new_n923), .B1(new_n925), .B2(new_n926), .ZN(G1352gat));
  NAND3_X1  g726(.A1(new_n871), .A2(new_n333), .A3(new_n924), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n871), .A2(KEYINPUT126), .A3(new_n333), .A4(new_n924), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n930), .A2(G204gat), .A3(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n722), .A2(G204gat), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n919), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n933), .B1(new_n919), .B2(new_n934), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n932), .A2(new_n937), .ZN(G1353gat));
  NAND4_X1  g737(.A1(new_n918), .A2(new_n921), .A3(new_n488), .A4(new_n306), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n871), .A2(new_n306), .A3(new_n924), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n940), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT63), .B1(new_n940), .B2(G211gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(G1354gat));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n867), .A2(new_n868), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT57), .B1(new_n945), .B2(new_n608), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n821), .A2(new_n870), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n944), .B(new_n924), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n697), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n944), .B1(new_n871), .B2(new_n924), .ZN(new_n950));
  OAI21_X1  g749(.A(G218gat), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n918), .A2(new_n921), .A3(new_n489), .A4(new_n697), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1355gat));
endmodule


