//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n555, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1133, new_n1134, new_n1135, new_n1136;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(KEYINPUT65), .A3(G125), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n475));
  NAND2_X1  g050(.A1(G101), .A2(G2104), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n476), .B1(new_n467), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G2105), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n473), .A2(new_n475), .A3(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(G160));
  OR2_X1    g058(.A1(new_n471), .A2(KEYINPUT67), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n471), .A2(KEYINPUT67), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n484), .A2(new_n485), .A3(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n484), .A2(new_n485), .A3(new_n479), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  OR2_X1    g066(.A1(G100), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G112), .C2(new_n479), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n488), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n497), .A2(new_n464), .A3(new_n466), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n471), .A2(new_n500), .A3(new_n497), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n464), .A2(new_n466), .A3(G126), .ZN(new_n503));
  NAND2_X1  g078(.A1(G114), .A2(G2104), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G2105), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n463), .A2(G2105), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G102), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n502), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT68), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G50), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n513), .B(new_n515), .C1(new_n521), .C2(new_n522), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G88), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n520), .A2(new_n526), .A3(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NAND2_X1  g106(.A1(new_n525), .A2(G51), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n528), .A2(G89), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n513), .A2(new_n515), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n534), .A2(G63), .A3(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n532), .A2(new_n533), .A3(new_n535), .A4(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  XOR2_X1   g114(.A(KEYINPUT69), .B(G52), .Z(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n524), .A2(new_n541), .B1(new_n542), .B2(new_n527), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n534), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n543), .B1(G651), .B2(new_n545), .ZN(G171));
  AOI22_X1  g121(.A1(new_n534), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G651), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n524), .A2(new_n550), .B1(new_n551), .B2(new_n527), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G188));
  INV_X1    g134(.A(G78), .ZN(new_n560));
  OR3_X1    g135(.A1(new_n560), .A2(new_n512), .A3(KEYINPUT71), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT71), .B1(new_n560), .B2(new_n512), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI211_X1 g138(.A(new_n561), .B(new_n562), .C1(new_n563), .C2(new_n516), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n564), .A2(G651), .B1(G91), .B2(new_n528), .ZN(new_n565));
  XOR2_X1   g140(.A(KEYINPUT70), .B(KEYINPUT9), .Z(new_n566));
  NAND3_X1  g141(.A1(new_n525), .A2(G53), .A3(new_n566), .ZN(new_n567));
  NOR2_X1   g142(.A1(KEYINPUT70), .A2(KEYINPUT9), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n524), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n565), .A2(new_n567), .A3(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  NAND2_X1  g147(.A1(new_n525), .A2(G49), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n534), .B2(G74), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n528), .A2(G87), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT72), .B1(new_n516), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT72), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n513), .A2(new_n515), .A3(new_n580), .A4(G61), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(G86), .B2(new_n528), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n525), .A2(G48), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G305));
  AOI22_X1  g160(.A1(new_n534), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n548), .ZN(new_n587));
  INV_X1    g162(.A(G47), .ZN(new_n588));
  INV_X1    g163(.A(G85), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n524), .A2(new_n588), .B1(new_n589), .B2(new_n527), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n528), .A2(G92), .ZN(new_n594));
  XOR2_X1   g169(.A(KEYINPUT73), .B(KEYINPUT10), .Z(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n516), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n525), .A2(G54), .B1(new_n599), .B2(G651), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n593), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n593), .B1(new_n602), .B2(G868), .ZN(G321));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(G299), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n605), .B2(G168), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(new_n605), .B2(G168), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n602), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT75), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n617), .B(new_n618), .C1(G111), .C2(new_n479), .ZN(new_n619));
  INV_X1    g194(.A(G123), .ZN(new_n620));
  INV_X1    g195(.A(G135), .ZN(new_n621));
  OAI221_X1 g196(.A(new_n619), .B1(new_n486), .B2(new_n620), .C1(new_n621), .C2(new_n489), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(G2096), .Z(new_n623));
  NAND2_X1  g198(.A1(new_n471), .A2(new_n507), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT74), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n627), .A2(G2100), .ZN(new_n628));
  AND2_X1   g203(.A1(new_n627), .A2(G2100), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n623), .B(new_n630), .C1(new_n628), .C2(new_n626), .ZN(G156));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT76), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  XOR2_X1   g209(.A(G2443), .B(G2446), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT77), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2427), .B(G2430), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(KEYINPUT14), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n638), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(G14), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT78), .Z(G401));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT79), .Z(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(G2072), .B(G2078), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT18), .Z(new_n653));
  XOR2_X1   g228(.A(new_n649), .B(KEYINPUT80), .Z(new_n654));
  OAI21_X1  g229(.A(KEYINPUT17), .B1(new_n654), .B2(new_n650), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(new_n651), .Z(new_n656));
  AND2_X1   g231(.A1(new_n654), .A2(new_n650), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n653), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2096), .B(G2100), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(G227));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n661));
  XOR2_X1   g236(.A(G1961), .B(G1966), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT81), .ZN(new_n663));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n661), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n663), .A2(new_n664), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n670), .A2(new_n667), .A3(new_n665), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n665), .A2(new_n661), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n672), .A2(new_n669), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n668), .B(new_n671), .C1(new_n673), .C2(new_n667), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G1986), .ZN(new_n675));
  INV_X1    g250(.A(G1981), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT82), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n677), .B(new_n681), .Z(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(G229));
  INV_X1    g258(.A(G29), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G26), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT90), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT28), .ZN(new_n687));
  OR2_X1    g262(.A1(G104), .A2(G2105), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n688), .B(G2104), .C1(G116), .C2(new_n479), .ZN(new_n689));
  INV_X1    g264(.A(G128), .ZN(new_n690));
  INV_X1    g265(.A(G140), .ZN(new_n691));
  OAI221_X1 g266(.A(new_n689), .B1(new_n486), .B2(new_n690), .C1(new_n691), .C2(new_n489), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT89), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n687), .B1(new_n694), .B2(G29), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT91), .ZN(new_n696));
  INV_X1    g271(.A(G2067), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(G29), .A2(G33), .ZN(new_n699));
  AOI22_X1  g274(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n700), .A2(new_n479), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n507), .A2(G103), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT92), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT25), .ZN(new_n704));
  AOI211_X1 g279(.A(new_n701), .B(new_n704), .C1(G139), .C2(new_n490), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT93), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n699), .B1(new_n706), .B2(G29), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(G2072), .Z(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G21), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G168), .B2(new_n709), .ZN(new_n711));
  INV_X1    g286(.A(G1966), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(G5), .A2(G16), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G171), .B2(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G1961), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n622), .A2(new_n684), .ZN(new_n717));
  INV_X1    g292(.A(G28), .ZN(new_n718));
  AOI21_X1  g293(.A(G29), .B1(new_n718), .B2(KEYINPUT30), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(KEYINPUT30), .B2(new_n718), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n713), .A2(new_n716), .A3(new_n717), .A4(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT31), .B(G11), .Z(new_n722));
  OAI21_X1  g297(.A(KEYINPUT96), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(G29), .A2(G32), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n490), .A2(G141), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n487), .A2(G129), .ZN(new_n726));
  NAND3_X1  g301(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT26), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n507), .A2(G105), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n725), .A2(new_n726), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n724), .B1(new_n730), .B2(new_n684), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT27), .B(G1996), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  INV_X1    g309(.A(new_n715), .ZN(new_n735));
  INV_X1    g310(.A(G1961), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n709), .A2(G19), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n553), .B2(new_n709), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n735), .A2(new_n736), .B1(G1341), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n733), .A2(new_n734), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n709), .A2(G4), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n602), .B2(new_n709), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1348), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n738), .A2(G1341), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n684), .A2(G27), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G164), .B2(new_n684), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2078), .ZN(new_n747));
  NOR4_X1   g322(.A1(new_n740), .A2(new_n743), .A3(new_n744), .A4(new_n747), .ZN(new_n748));
  OR3_X1    g323(.A1(new_n721), .A2(KEYINPUT96), .A3(new_n722), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n708), .A2(new_n723), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT23), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n709), .A2(G20), .ZN(new_n752));
  AOI211_X1 g327(.A(new_n751), .B(new_n752), .C1(G299), .C2(G16), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n751), .B2(new_n752), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT98), .B(G1956), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n684), .A2(G35), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G162), .B2(new_n684), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n756), .B1(G2090), .B2(new_n760), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT99), .Z(new_n762));
  NAND2_X1  g337(.A1(G160), .A2(G29), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT24), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n684), .B1(new_n764), .B2(G34), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT94), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n764), .A2(G34), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n765), .A2(new_n766), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n763), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT95), .ZN(new_n772));
  INV_X1    g347(.A(G2084), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G2090), .B2(new_n760), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n750), .A2(new_n762), .A3(new_n775), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n709), .A2(G6), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G305), .B2(G16), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT86), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT32), .B(G1981), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n709), .A2(G23), .ZN(new_n782));
  INV_X1    g357(.A(G288), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n709), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT33), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1976), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n709), .A2(G22), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G166), .B2(new_n709), .ZN(new_n788));
  INV_X1    g363(.A(G1971), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n781), .A2(new_n786), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT87), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT34), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n791), .A2(KEYINPUT87), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n791), .A2(KEYINPUT87), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n795), .A2(KEYINPUT34), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n709), .A2(G24), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n591), .B2(new_n709), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT85), .B(G1986), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(G25), .A2(G29), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n487), .A2(G119), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n490), .A2(G131), .ZN(new_n804));
  OR2_X1    g379(.A1(G95), .A2(G2105), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n805), .B(G2104), .C1(G107), .C2(new_n479), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT83), .Z(new_n807));
  NAND3_X1  g382(.A1(new_n803), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n802), .B1(new_n809), .B2(G29), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT84), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT35), .B(G1991), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n811), .B(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n794), .A2(new_n797), .A3(new_n801), .A4(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(KEYINPUT88), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(KEYINPUT88), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT36), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(KEYINPUT36), .B1(new_n816), .B2(new_n817), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n698), .B(new_n776), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(G311));
  XNOR2_X1  g398(.A(new_n818), .B(new_n819), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT100), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n824), .A2(new_n825), .A3(new_n698), .A4(new_n776), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n822), .A2(KEYINPUT100), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(G150));
  NAND2_X1  g403(.A1(new_n528), .A2(G93), .ZN(new_n829));
  INV_X1    g404(.A(G55), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n534), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n831));
  OAI221_X1 g406(.A(new_n829), .B1(new_n524), .B2(new_n830), .C1(new_n831), .C2(new_n548), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G860), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT101), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT37), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n602), .A2(G559), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT38), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n553), .B(new_n832), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT39), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n837), .B(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n835), .B1(new_n840), .B2(G860), .ZN(G145));
  XNOR2_X1  g416(.A(new_n693), .B(new_n730), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G164), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n843), .A2(new_n706), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n705), .B2(new_n843), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n808), .B(new_n625), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n487), .A2(G130), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n490), .A2(G142), .ZN(new_n848));
  NOR2_X1   g423(.A1(G106), .A2(G2105), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(new_n479), .B2(G118), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n847), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n846), .B(new_n851), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n845), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n853), .A2(KEYINPUT102), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n494), .B(new_n622), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(G160), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n845), .A2(new_n852), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n853), .A2(KEYINPUT102), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(G37), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT103), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n845), .A2(KEYINPUT103), .A3(new_n852), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n863), .A2(new_n853), .A3(new_n864), .A4(new_n856), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n860), .A2(new_n861), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g442(.A1(new_n832), .A2(G868), .ZN(new_n868));
  XNOR2_X1  g443(.A(G303), .B(G305), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n591), .B(G288), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT104), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n870), .A2(KEYINPUT104), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(new_n869), .B2(new_n872), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT105), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(new_n876), .B2(KEYINPUT42), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(KEYINPUT42), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n877), .B(new_n878), .Z(new_n879));
  INV_X1    g454(.A(KEYINPUT106), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n601), .B(G299), .Z(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(KEYINPUT41), .Z(new_n882));
  XNOR2_X1  g457(.A(new_n611), .B(new_n838), .ZN(new_n883));
  MUX2_X1   g458(.A(new_n881), .B(new_n882), .S(new_n883), .Z(new_n884));
  OAI21_X1  g459(.A(new_n879), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n880), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n885), .B(new_n886), .Z(new_n887));
  AOI21_X1  g462(.A(new_n868), .B1(new_n887), .B2(G868), .ZN(G295));
  AOI21_X1  g463(.A(new_n868), .B1(new_n887), .B2(G868), .ZN(G331));
  XNOR2_X1  g464(.A(new_n838), .B(G171), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(G286), .ZN(new_n891));
  MUX2_X1   g466(.A(new_n881), .B(new_n882), .S(new_n891), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n875), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n861), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT43), .ZN(new_n895));
  NAND2_X1  g470(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n897), .B(new_n898), .ZN(G397));
  AOI22_X1  g474(.A1(new_n471), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT66), .B1(new_n900), .B2(G2105), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n901), .B1(G2105), .B2(new_n473), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n473), .A2(new_n475), .A3(G2105), .ZN(new_n903));
  OAI21_X1  g478(.A(G40), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(G1384), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n509), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT45), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n693), .B(new_n697), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n909), .B1(new_n910), .B2(new_n730), .ZN(new_n911));
  INV_X1    g486(.A(G1996), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(KEYINPUT122), .A2(KEYINPUT46), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n913), .B(new_n914), .Z(new_n915));
  OAI211_X1 g490(.A(new_n911), .B(new_n915), .C1(KEYINPUT122), .C2(KEYINPUT46), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT123), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT47), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(G290), .A2(G1986), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n909), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT48), .ZN(new_n922));
  INV_X1    g497(.A(new_n910), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n730), .B(new_n912), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n809), .A2(new_n813), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n927), .B1(new_n812), .B2(new_n808), .ZN(new_n928));
  INV_X1    g503(.A(new_n909), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n922), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n917), .A2(new_n918), .ZN(new_n931));
  INV_X1    g506(.A(new_n925), .ZN(new_n932));
  OAI22_X1  g507(.A1(new_n932), .A2(new_n926), .B1(G2067), .B2(new_n694), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n909), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n919), .A2(new_n930), .A3(new_n931), .A4(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT124), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n935), .B(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT63), .ZN(new_n938));
  XOR2_X1   g513(.A(KEYINPUT110), .B(G8), .Z(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n906), .A2(KEYINPUT108), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n509), .A2(new_n942), .A3(new_n905), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G40), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n945), .B1(new_n481), .B2(new_n482), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n940), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n783), .A2(G1976), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT52), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G1976), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT52), .B1(G288), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n947), .A2(new_n948), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n904), .B1(new_n941), .B2(new_n943), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n582), .A2(G651), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n676), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(G305), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT111), .B1(new_n582), .B2(G651), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n583), .B(new_n584), .C1(new_n961), .C2(new_n676), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT49), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n956), .A2(new_n963), .A3(new_n940), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n960), .A2(KEYINPUT49), .A3(new_n962), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT112), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n960), .A2(new_n967), .A3(new_n962), .A4(KEYINPUT49), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n964), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT113), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n964), .A2(new_n972), .A3(new_n969), .ZN(new_n973));
  AOI211_X1 g548(.A(new_n951), .B(new_n955), .C1(new_n971), .C2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n509), .A2(KEYINPUT45), .A3(new_n905), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n946), .A2(new_n975), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n509), .A2(new_n942), .A3(new_n905), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n942), .B1(new_n509), .B2(new_n905), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n977), .A2(new_n978), .A3(KEYINPUT45), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n712), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(new_n977), .B2(new_n978), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n906), .A2(KEYINPUT50), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n982), .A2(new_n773), .A3(new_n946), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n985), .A2(G168), .A3(new_n939), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n946), .A2(new_n908), .A3(new_n975), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n789), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n982), .A2(new_n946), .A3(new_n983), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n988), .B1(new_n989), .B2(G2090), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT109), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n988), .B(new_n992), .C1(new_n989), .C2(G2090), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(G8), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(G303), .A2(G8), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n995), .A2(KEYINPUT55), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(KEYINPUT55), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n986), .B1(new_n994), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n938), .B1(new_n974), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n973), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n972), .B1(new_n964), .B2(new_n969), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n950), .B(new_n954), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n986), .A2(KEYINPUT63), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n977), .A2(new_n978), .A3(new_n981), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT114), .B1(new_n1006), .B2(new_n904), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1008), .B(new_n946), .C1(new_n944), .C2(new_n981), .ZN(new_n1009));
  INV_X1    g584(.A(G2090), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n509), .A2(new_n981), .A3(new_n905), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n940), .B1(new_n1012), .B2(new_n988), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1005), .B1(new_n998), .B2(new_n1013), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n991), .A2(G8), .A3(new_n998), .A4(new_n993), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1004), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n947), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n952), .B(new_n783), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n583), .A2(new_n676), .A3(new_n584), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1001), .A2(new_n1016), .A3(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT56), .B(G2072), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n987), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1007), .A2(new_n1011), .A3(new_n1009), .ZN(new_n1025));
  INV_X1    g600(.A(G1956), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1024), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(G299), .B(KEYINPUT57), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1348), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n989), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n956), .A2(new_n697), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n904), .B1(new_n944), .B2(new_n981), .ZN(new_n1036));
  AOI21_X1  g611(.A(G1348), .B1(new_n1036), .B2(new_n983), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n944), .A2(new_n697), .A3(new_n946), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT115), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1030), .A2(new_n602), .A3(new_n1035), .A4(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1028), .B1(new_n1041), .B2(new_n1024), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT61), .B1(new_n1042), .B2(new_n1030), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1045));
  AOI211_X1 g620(.A(new_n1028), .B(new_n1024), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT61), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1032), .A2(new_n1034), .A3(new_n1033), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1034), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT60), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT60), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1039), .A2(new_n1053), .A3(new_n1035), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(new_n1054), .A3(new_n602), .ZN(new_n1055));
  OAI211_X1 g630(.A(KEYINPUT60), .B(new_n601), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT58), .B(G1341), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n956), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n987), .A2(G1996), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n553), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1060), .B1(new_n1061), .B2(KEYINPUT59), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(KEYINPUT59), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1061), .A2(KEYINPUT59), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n553), .B(new_n1064), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1062), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1055), .A2(new_n1056), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1043), .B1(new_n1049), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G2078), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n946), .A2(new_n1069), .A3(new_n908), .A4(new_n975), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT118), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n989), .A2(new_n736), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1070), .A2(new_n1075), .A3(new_n1071), .ZN(new_n1076));
  INV_X1    g651(.A(new_n975), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(G2078), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n474), .A2(KEYINPUT53), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1079), .B1(new_n479), .B2(new_n478), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1078), .A2(G40), .A3(new_n908), .A4(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .A4(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(G171), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n904), .A2(new_n1077), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n941), .A2(new_n907), .A3(new_n943), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1085), .A2(KEYINPUT53), .A3(new_n1069), .A4(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .A4(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT54), .B1(new_n1088), .B2(G171), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT119), .B1(new_n1084), .B2(new_n1089), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1088), .A2(G171), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT119), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1091), .A2(new_n1092), .A3(KEYINPUT54), .A4(new_n1083), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(G168), .A2(new_n940), .ZN(new_n1095));
  AOI211_X1 g670(.A(KEYINPUT51), .B(new_n1095), .C1(new_n985), .C2(new_n939), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n980), .A2(KEYINPUT117), .A3(new_n984), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT117), .B1(new_n980), .B2(new_n984), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1095), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1097), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(G8), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1096), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1015), .B1(new_n998), .B2(new_n1013), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1106), .A2(new_n1004), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1088), .A2(G171), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1082), .A2(G171), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1108), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1094), .A2(new_n1105), .A3(new_n1107), .A4(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1021), .B1(new_n1068), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1105), .A2(KEYINPUT62), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1105), .A2(KEYINPUT62), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1116), .A2(new_n1109), .A3(new_n1117), .A4(new_n1107), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1021), .B(KEYINPUT120), .C1(new_n1068), .C2(new_n1112), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1115), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n1121));
  INV_X1    g696(.A(G1986), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n928), .B1(new_n1122), .B2(new_n591), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n909), .B1(new_n1123), .B2(new_n920), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1120), .A2(new_n1121), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1121), .B1(new_n1120), .B2(new_n1124), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n937), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g704(.A(KEYINPUT125), .B(new_n937), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g706(.A1(G227), .A2(new_n460), .ZN(new_n1133));
  AOI21_X1  g707(.A(G401), .B1(KEYINPUT126), .B2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g708(.A(new_n1134), .B(new_n682), .C1(KEYINPUT126), .C2(new_n1133), .ZN(new_n1135));
  XOR2_X1   g709(.A(new_n1135), .B(KEYINPUT127), .Z(new_n1136));
  NAND3_X1  g710(.A1(new_n1136), .A2(new_n895), .A3(new_n866), .ZN(G225));
  INV_X1    g711(.A(G225), .ZN(G308));
endmodule


