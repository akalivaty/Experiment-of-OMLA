//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G469), .ZN(new_n191));
  INV_X1    g005(.A(G902), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT80), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT79), .ZN(new_n195));
  INV_X1    g009(.A(G104), .ZN(new_n196));
  AOI22_X1  g010(.A1(new_n195), .A2(KEYINPUT3), .B1(new_n196), .B2(G107), .ZN(new_n197));
  OAI22_X1  g011(.A1(new_n195), .A2(KEYINPUT3), .B1(new_n196), .B2(G107), .ZN(new_n198));
  INV_X1    g012(.A(G101), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n200));
  INV_X1    g014(.A(G107), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n200), .A2(new_n201), .A3(KEYINPUT79), .A4(G104), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n197), .A2(new_n198), .A3(new_n199), .A4(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n201), .A2(G104), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n196), .A2(G107), .ZN(new_n205));
  OAI21_X1  g019(.A(G101), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(G146), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT64), .A3(G143), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n210), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT1), .B1(new_n209), .B2(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G128), .ZN(new_n216));
  XNOR2_X1  g030(.A(G143), .B(G146), .ZN(new_n217));
  INV_X1    g031(.A(G128), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n214), .A2(new_n216), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n207), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n212), .A2(G143), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n222), .A3(new_n211), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n218), .B1(new_n222), .B2(KEYINPUT1), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n223), .B1(new_n224), .B2(new_n217), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(new_n203), .A3(new_n206), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT66), .B(G131), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n228));
  INV_X1    g042(.A(G134), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n228), .A2(KEYINPUT11), .B1(new_n229), .B2(G137), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT11), .ZN(new_n231));
  INV_X1    g045(.A(G137), .ZN(new_n232));
  AND4_X1   g046(.A1(KEYINPUT65), .A2(new_n231), .A3(new_n232), .A4(G134), .ZN(new_n233));
  AOI22_X1  g047(.A1(KEYINPUT65), .A2(new_n231), .B1(new_n232), .B2(G134), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n227), .B(new_n230), .C1(new_n233), .C2(new_n234), .ZN(new_n235));
  OAI22_X1  g049(.A1(new_n228), .A2(KEYINPUT11), .B1(new_n229), .B2(G137), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n231), .A2(new_n232), .A3(KEYINPUT65), .A4(G134), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n230), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G131), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n221), .A2(new_n226), .B1(new_n235), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n194), .B1(new_n241), .B2(KEYINPUT12), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n221), .A2(new_n226), .ZN(new_n243));
  OAI22_X1  g057(.A1(KEYINPUT65), .A2(new_n231), .B1(new_n232), .B2(G134), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n244), .B1(new_n236), .B2(new_n237), .ZN(new_n245));
  INV_X1    g059(.A(G131), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n235), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT12), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n242), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n197), .A2(new_n198), .A3(new_n202), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G101), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT4), .A3(new_n203), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n252), .A2(new_n255), .A3(G101), .ZN(new_n256));
  AND2_X1   g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n214), .A2(new_n259), .B1(new_n217), .B2(new_n257), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n254), .A2(new_n256), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n247), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT10), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n226), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n214), .A2(new_n216), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n223), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n266), .A2(KEYINPUT10), .A3(new_n203), .A4(new_n206), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n261), .A2(new_n262), .A3(new_n264), .A4(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(G110), .B(G140), .ZN(new_n269));
  INV_X1    g083(.A(G227), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(G953), .ZN(new_n271));
  XOR2_X1   g085(.A(new_n269), .B(new_n271), .Z(new_n272));
  NAND3_X1  g086(.A1(new_n248), .A2(new_n194), .A3(new_n249), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n251), .A2(new_n268), .A3(new_n272), .A4(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n261), .A2(new_n264), .A3(new_n267), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n247), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n268), .ZN(new_n277));
  INV_X1    g091(.A(new_n272), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(G902), .B1(new_n274), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n193), .B1(new_n280), .B2(new_n191), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n251), .A2(new_n268), .A3(new_n273), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n278), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n276), .A2(new_n268), .A3(new_n272), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(G469), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n190), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(G214), .B1(G237), .B2(G902), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT69), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT2), .ZN(new_n289));
  INV_X1    g103(.A(G113), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT69), .B1(KEYINPUT2), .B2(G113), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(KEYINPUT2), .A2(G113), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(G116), .B(G119), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n293), .A2(new_n294), .A3(new_n296), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n254), .A2(new_n300), .A3(new_n256), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT81), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT5), .ZN(new_n304));
  INV_X1    g118(.A(G119), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(G116), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n306), .B1(new_n297), .B2(new_n304), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n299), .B1(new_n307), .B2(new_n290), .ZN(new_n308));
  OR2_X1    g122(.A1(new_n308), .A2(new_n207), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n254), .A2(new_n300), .A3(KEYINPUT81), .A4(new_n256), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n303), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(G110), .B(G122), .ZN(new_n312));
  XOR2_X1   g126(.A(new_n312), .B(KEYINPUT82), .Z(new_n313));
  AND2_X1   g127(.A1(new_n313), .A2(KEYINPUT83), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT6), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n303), .A2(new_n312), .A3(new_n309), .A4(new_n310), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n311), .A2(KEYINPUT6), .A3(new_n314), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n260), .A2(G125), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(G125), .B2(new_n220), .ZN(new_n322));
  INV_X1    g136(.A(G224), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(G953), .ZN(new_n324));
  XOR2_X1   g138(.A(new_n322), .B(new_n324), .Z(new_n325));
  AOI21_X1  g139(.A(G902), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(G210), .B1(G237), .B2(G902), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n325), .B1(KEYINPUT7), .B2(new_n324), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n308), .B(new_n207), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n312), .B(KEYINPUT8), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OR3_X1    g145(.A1(new_n322), .A2(KEYINPUT7), .A3(new_n324), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n328), .A2(new_n318), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n326), .A2(new_n327), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n327), .B1(new_n326), .B2(new_n333), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n286), .B(new_n287), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G478), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(KEYINPUT15), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT88), .ZN(new_n340));
  XOR2_X1   g154(.A(KEYINPUT86), .B(KEYINPUT13), .Z(new_n341));
  NOR2_X1   g155(.A1(new_n218), .A2(G143), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT87), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n209), .A2(G128), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n344), .B1(new_n341), .B2(new_n342), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT86), .B(KEYINPUT13), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT87), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n346), .B(new_n347), .C1(new_n218), .C2(G143), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n343), .A2(new_n345), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G134), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n342), .A2(new_n344), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n229), .ZN(new_n352));
  XNOR2_X1  g166(.A(G116), .B(G122), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT85), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT85), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n201), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n355), .A2(new_n357), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(G107), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n350), .B(new_n352), .C1(new_n358), .C2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n351), .B(new_n229), .ZN(new_n362));
  INV_X1    g176(.A(G116), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(KEYINPUT14), .A3(G122), .ZN(new_n364));
  OAI211_X1 g178(.A(G107), .B(new_n364), .C1(new_n354), .C2(KEYINPUT14), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n362), .B(new_n365), .C1(G107), .C2(new_n359), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G217), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n188), .A2(new_n368), .A3(G953), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n361), .A2(new_n366), .A3(new_n369), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n340), .B1(new_n373), .B2(new_n192), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n361), .A2(new_n366), .A3(new_n369), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n369), .B1(new_n361), .B2(new_n366), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n340), .B(new_n192), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n339), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n192), .B1(new_n375), .B2(new_n376), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n339), .B1(new_n380), .B2(KEYINPUT88), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G953), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G952), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n385), .B1(G234), .B2(G237), .ZN(new_n386));
  XOR2_X1   g200(.A(KEYINPUT21), .B(G898), .Z(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(G234), .A2(G237), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(G902), .A3(G953), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n386), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G475), .ZN(new_n393));
  XOR2_X1   g207(.A(G125), .B(G140), .Z(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT19), .ZN(new_n395));
  XNOR2_X1  g209(.A(G125), .B(G140), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT19), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n395), .A2(new_n212), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G125), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n400), .A2(KEYINPUT16), .A3(G140), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT16), .ZN(new_n403));
  OAI211_X1 g217(.A(G146), .B(new_n402), .C1(new_n394), .C2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G237), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(new_n384), .A3(G214), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n209), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n405), .A2(new_n384), .A3(G143), .A4(G214), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n227), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n407), .A2(new_n227), .A3(new_n408), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n399), .B(new_n404), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT84), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n407), .A2(new_n408), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(KEYINPUT18), .A3(G131), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n394), .A2(G146), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n396), .A2(new_n212), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(KEYINPUT18), .A2(G131), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n407), .A2(new_n408), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n414), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n411), .A2(new_n412), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n412), .B1(new_n411), .B2(new_n420), .ZN(new_n423));
  XNOR2_X1  g237(.A(G113), .B(G122), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(new_n196), .ZN(new_n425));
  NOR3_X1   g239(.A1(new_n422), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n402), .B1(new_n394), .B2(new_n403), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n212), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n428), .A2(new_n404), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n409), .A2(KEYINPUT17), .ZN(new_n430));
  OR2_X1    g244(.A1(new_n410), .A2(new_n409), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n429), .B(new_n430), .C1(new_n431), .C2(KEYINPUT17), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n432), .A2(new_n425), .A3(new_n420), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n393), .B(new_n192), .C1(new_n426), .C2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT20), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n425), .B1(new_n432), .B2(new_n420), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n192), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G475), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n423), .A2(new_n425), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n421), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n432), .A2(new_n425), .A3(new_n420), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n443), .A2(KEYINPUT20), .A3(new_n393), .A4(new_n192), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n436), .A2(new_n439), .A3(new_n444), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n383), .A2(new_n392), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n337), .A2(new_n446), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n238), .A2(new_n227), .A3(new_n230), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n246), .B1(new_n238), .B2(new_n230), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n260), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n232), .A2(G134), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n229), .A2(G137), .ZN(new_n452));
  OAI21_X1  g266(.A(G131), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n266), .A2(new_n235), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(new_n300), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(KEYINPUT72), .ZN(new_n457));
  INV_X1    g271(.A(new_n300), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n450), .A2(new_n454), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n455), .A2(KEYINPUT72), .A3(new_n300), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(KEYINPUT28), .A3(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n456), .A2(KEYINPUT28), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  XOR2_X1   g278(.A(KEYINPUT26), .B(G101), .Z(new_n465));
  NAND3_X1  g279(.A1(new_n405), .A2(new_n384), .A3(G210), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n468));
  XOR2_X1   g282(.A(new_n467), .B(new_n468), .Z(new_n469));
  NAND4_X1  g283(.A1(new_n462), .A2(KEYINPUT29), .A3(new_n464), .A4(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n469), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT67), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n450), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n247), .A2(KEYINPUT67), .A3(new_n260), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT68), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n454), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n266), .A2(KEYINPUT68), .A3(new_n235), .A4(new_n453), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n473), .A2(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT71), .B1(new_n478), .B2(new_n458), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT67), .B1(new_n247), .B2(new_n260), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n247), .A2(KEYINPUT67), .A3(new_n260), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n265), .A2(new_n223), .B1(new_n245), .B2(new_n227), .ZN(new_n482));
  AOI21_X1  g296(.A(KEYINPUT68), .B1(new_n482), .B2(new_n453), .ZN(new_n483));
  AND4_X1   g297(.A1(KEYINPUT68), .A2(new_n266), .A3(new_n235), .A4(new_n453), .ZN(new_n484));
  OAI22_X1  g298(.A1(new_n480), .A2(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT71), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n486), .A3(new_n300), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n459), .A2(new_n458), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n479), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI211_X1 g303(.A(new_n463), .B(new_n471), .C1(new_n489), .C2(KEYINPUT28), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT30), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n455), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n493), .B(new_n300), .C1(new_n478), .C2(KEYINPUT30), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n488), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n471), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT29), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n192), .B(new_n470), .C1(new_n490), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(G472), .ZN(new_n500));
  NOR2_X1   g314(.A1(G472), .A2(G902), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT28), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n485), .A2(new_n300), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n456), .B1(new_n504), .B2(KEYINPUT71), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n503), .B1(new_n505), .B2(new_n487), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n471), .B1(new_n506), .B2(new_n463), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n494), .A2(new_n488), .A3(new_n469), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT31), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n494), .A2(KEYINPUT31), .A3(new_n488), .A4(new_n469), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI211_X1 g326(.A(KEYINPUT32), .B(new_n502), .C1(new_n507), .C2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT32), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n492), .B1(new_n485), .B2(new_n491), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n456), .B1(new_n515), .B2(new_n300), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT31), .B1(new_n516), .B2(new_n469), .ZN(new_n517));
  INV_X1    g331(.A(new_n511), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n463), .B1(new_n489), .B2(KEYINPUT28), .ZN(new_n519));
  OAI22_X1  g333(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n469), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n514), .B1(new_n520), .B2(new_n501), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n500), .B1(new_n513), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT73), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n305), .A2(G128), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n523), .B(KEYINPUT23), .C1(new_n524), .C2(KEYINPUT74), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n305), .A2(G128), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT23), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n218), .A2(G119), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n527), .B1(new_n528), .B2(KEYINPUT73), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT74), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT73), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n525), .B(new_n526), .C1(new_n529), .C2(new_n531), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n526), .A2(new_n528), .ZN(new_n533));
  XOR2_X1   g347(.A(KEYINPUT24), .B(G110), .Z(new_n534));
  OAI22_X1  g348(.A1(new_n532), .A2(G110), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(new_n416), .A3(new_n404), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT76), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n532), .A2(KEYINPUT75), .A3(G110), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT75), .B1(new_n532), .B2(G110), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n428), .A2(new_n404), .B1(new_n533), .B2(new_n534), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n537), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n532), .A2(G110), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT75), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n532), .A2(KEYINPUT75), .A3(G110), .ZN(new_n546));
  AND4_X1   g360(.A1(new_n537), .A2(new_n541), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n536), .B1(new_n542), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n384), .A2(G221), .A3(G234), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(KEYINPUT22), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(G137), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n536), .B(new_n551), .C1(new_n542), .C2(new_n547), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(new_n192), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT77), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT25), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n368), .B1(G234), .B2(new_n192), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT25), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n560), .A2(G902), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n553), .A2(new_n554), .A3(new_n563), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n522), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT78), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n562), .A2(new_n564), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n473), .A2(new_n474), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n476), .A2(new_n477), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n458), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n488), .B1(new_n571), .B2(new_n486), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n478), .A2(KEYINPUT71), .A3(new_n458), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT28), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n464), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n575), .A2(new_n471), .B1(new_n510), .B2(new_n511), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT32), .B1(new_n576), .B2(new_n502), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n520), .A2(new_n514), .A3(new_n501), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n568), .B1(new_n579), .B2(new_n500), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT78), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n447), .B1(new_n567), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(new_n199), .ZN(G3));
  INV_X1    g398(.A(new_n392), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n287), .B(new_n585), .C1(new_n334), .C2(new_n335), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT89), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT33), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(KEYINPUT89), .A2(KEYINPUT33), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n373), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n371), .A2(new_n587), .A3(new_n588), .A4(new_n372), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(G478), .A3(new_n192), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n380), .A2(new_n338), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n445), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT90), .B1(new_n586), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n597), .ZN(new_n599));
  INV_X1    g413(.A(new_n287), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n320), .A2(new_n325), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n601), .A2(new_n192), .A3(new_n333), .ZN(new_n602));
  INV_X1    g416(.A(new_n327), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n326), .A2(new_n327), .A3(new_n333), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n600), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT90), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n599), .A2(new_n606), .A3(new_n607), .A4(new_n585), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n598), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n507), .B2(new_n512), .ZN(new_n610));
  INV_X1    g424(.A(G472), .ZN(new_n611));
  OAI22_X1  g425(.A1(new_n610), .A2(new_n611), .B1(new_n576), .B2(new_n502), .ZN(new_n612));
  INV_X1    g426(.A(new_n286), .ZN(new_n613));
  OR3_X1    g427(.A1(new_n612), .A2(new_n613), .A3(new_n568), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT34), .B(G104), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT91), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n615), .B(new_n617), .ZN(G6));
  NAND2_X1  g432(.A1(new_n380), .A2(KEYINPUT88), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n377), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n381), .B1(new_n620), .B2(new_n339), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n586), .A2(new_n621), .A3(new_n445), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n614), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT35), .B(G107), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  NOR2_X1   g440(.A1(new_n552), .A2(KEYINPUT36), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n548), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n563), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT25), .ZN(new_n631));
  AOI21_X1  g445(.A(KEYINPUT25), .B1(new_n555), .B2(new_n556), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n630), .B1(new_n633), .B2(new_n560), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n447), .A2(new_n612), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G110), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT92), .B(KEYINPUT37), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G12));
  NAND2_X1  g452(.A1(new_n562), .A2(new_n629), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT93), .B(G900), .Z(new_n640));
  AOI21_X1  g454(.A(new_n386), .B1(new_n391), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n436), .A2(new_n439), .A3(new_n444), .A4(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT94), .B1(new_n644), .B2(new_n383), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT94), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n621), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n522), .A2(new_n337), .A3(new_n639), .A4(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT95), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n634), .B1(new_n579), .B2(new_n500), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n652), .A2(KEYINPUT95), .A3(new_n337), .A4(new_n648), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G128), .ZN(G30));
  INV_X1    g469(.A(new_n445), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(new_n621), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n641), .B(KEYINPUT39), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n613), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n662), .B(new_n287), .C1(new_n661), .C2(new_n660), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n460), .A2(new_n461), .ZN(new_n664));
  AOI21_X1  g478(.A(G902), .B1(new_n664), .B2(new_n471), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n495), .A2(new_n469), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n611), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n667), .B1(new_n577), .B2(new_n578), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n334), .A2(new_n335), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT38), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n604), .A2(new_n605), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT38), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  NOR4_X1   g488(.A1(new_n663), .A2(new_n639), .A3(new_n668), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(new_n209), .ZN(G45));
  AND3_X1   g490(.A1(new_n522), .A2(new_n337), .A3(new_n639), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n597), .A2(new_n641), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT96), .B(G146), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G48));
  NAND2_X1  g495(.A1(new_n274), .A2(new_n279), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(G469), .B1(new_n683), .B2(G902), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n280), .A2(new_n191), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n684), .A2(new_n189), .A3(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n580), .A2(new_n608), .A3(new_n598), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT41), .B(G113), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G15));
  NAND3_X1  g503(.A1(new_n580), .A2(new_n622), .A3(new_n686), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G116), .ZN(G18));
  NAND2_X1  g505(.A1(new_n606), .A2(new_n686), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n652), .A2(new_n446), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G119), .ZN(G21));
  AND2_X1   g509(.A1(new_n462), .A2(new_n464), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n512), .B1(new_n696), .B2(new_n469), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n501), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n698), .B1(new_n610), .B2(new_n611), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n568), .ZN(new_n700));
  INV_X1    g514(.A(new_n586), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n700), .A2(new_n701), .A3(new_n657), .A4(new_n686), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G122), .ZN(G24));
  INV_X1    g517(.A(KEYINPUT97), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n704), .B1(new_n699), .B2(new_n634), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n520), .A2(new_n192), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(G472), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n639), .A2(KEYINPUT97), .A3(new_n707), .A4(new_n698), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(new_n678), .A3(new_n693), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  INV_X1    g525(.A(KEYINPUT98), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n283), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n282), .A2(KEYINPUT98), .A3(new_n278), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n713), .A2(G469), .A3(new_n284), .A4(new_n714), .ZN(new_n715));
  OR2_X1    g529(.A1(new_n715), .A2(KEYINPUT99), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(KEYINPUT99), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n281), .A3(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT100), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n718), .A2(new_n719), .A3(new_n189), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n719), .B1(new_n718), .B2(new_n189), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n669), .A2(new_n287), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n723), .A2(new_n580), .A3(new_n678), .A4(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n718), .A2(new_n189), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n722), .B1(new_n727), .B2(KEYINPUT100), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n718), .A2(new_n719), .A3(new_n189), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(new_n580), .A3(new_n678), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n726), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(KEYINPUT102), .B(G131), .Z(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G33));
  NAND4_X1  g549(.A1(new_n728), .A2(new_n580), .A3(new_n648), .A4(new_n729), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT103), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT104), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n229), .ZN(G36));
  NAND2_X1  g554(.A1(new_n283), .A2(new_n284), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n713), .A2(new_n284), .A3(new_n714), .ZN(new_n744));
  OAI211_X1 g558(.A(G469), .B(new_n743), .C1(new_n744), .C2(new_n742), .ZN(new_n745));
  INV_X1    g559(.A(new_n193), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT46), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT105), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n747), .A2(KEYINPUT46), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT105), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n747), .A2(new_n751), .A3(KEYINPUT46), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n749), .A2(new_n750), .A3(new_n685), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n189), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n754), .A2(new_n659), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n596), .A2(new_n656), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT43), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n612), .A3(new_n639), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n722), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n755), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  INV_X1    g581(.A(KEYINPUT47), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n754), .B(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n678), .ZN(new_n770));
  NOR4_X1   g584(.A1(new_n770), .A2(new_n522), .A3(new_n565), .A4(new_n722), .ZN(new_n771));
  XOR2_X1   g585(.A(new_n771), .B(KEYINPUT106), .Z(new_n772));
  NAND2_X1  g586(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G140), .ZN(G42));
  NAND3_X1  g588(.A1(new_n562), .A2(new_n629), .A3(new_n642), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT110), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n775), .B(new_n776), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n606), .A2(new_n657), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n727), .A2(new_n668), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n654), .A2(new_n679), .A3(new_n710), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT52), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n687), .A2(new_n690), .A3(new_n694), .A4(new_n702), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n783), .B1(new_n726), .B2(new_n732), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n770), .B1(new_n705), .B2(new_n708), .ZN(new_n785));
  AOI22_X1  g599(.A1(new_n785), .A2(new_n693), .B1(new_n677), .B2(new_n678), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n786), .A2(new_n787), .A3(new_n654), .A4(new_n780), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n723), .A2(new_n785), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT109), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n723), .A2(new_n785), .A3(KEYINPUT109), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n782), .A2(new_n784), .A3(new_n788), .A4(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n383), .A2(KEYINPUT107), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT107), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n621), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n656), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT108), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n799), .B1(new_n798), .B2(new_n597), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n701), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n614), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n803), .A2(new_n583), .A3(new_n635), .ZN(new_n804));
  NOR4_X1   g618(.A1(new_n613), .A2(new_n795), .A3(new_n797), .A4(new_n643), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n671), .A2(new_n600), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n652), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n804), .A2(new_n738), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n794), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT112), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n782), .A2(new_n784), .A3(new_n810), .A4(new_n788), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT53), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(KEYINPUT53), .B(new_n811), .C1(new_n794), .C2(new_n808), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT54), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n809), .A2(KEYINPUT53), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT111), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n809), .A2(KEYINPUT53), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT111), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n809), .A2(new_n819), .A3(KEYINPUT53), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n817), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n815), .B1(new_n821), .B2(KEYINPUT54), .ZN(new_n822));
  INV_X1    g636(.A(new_n386), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n758), .B2(new_n760), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n693), .A3(new_n700), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n806), .A2(new_n686), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n580), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT48), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n824), .A2(new_n700), .A3(new_n806), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT113), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n684), .A2(new_n685), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n189), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n833), .B1(new_n769), .B2(new_n836), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n699), .A2(new_n568), .A3(new_n190), .A4(new_n835), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n287), .B1(new_n670), .B2(new_n673), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n824), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT50), .ZN(new_n841));
  OR3_X1    g655(.A1(new_n840), .A2(KEYINPUT117), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT117), .B1(new_n840), .B2(new_n841), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n840), .B2(KEYINPUT114), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n838), .A2(new_n824), .A3(new_n848), .A4(new_n839), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n847), .B1(new_n846), .B2(new_n849), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n844), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n829), .A2(new_n709), .ZN(new_n853));
  AND4_X1   g667(.A1(new_n386), .A2(new_n827), .A3(new_n565), .A4(new_n668), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n854), .A2(new_n656), .A3(new_n595), .A4(new_n594), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n837), .A2(new_n852), .A3(new_n853), .A4(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n385), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n852), .A2(new_n857), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(KEYINPUT51), .A3(new_n837), .A4(new_n853), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n854), .A2(new_n599), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n831), .A2(new_n860), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n822), .A2(new_n825), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n865), .B1(G952), .B2(G953), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n757), .B(new_n189), .C1(KEYINPUT49), .C2(new_n835), .ZN(new_n867));
  AOI211_X1 g681(.A(new_n568), .B(new_n867), .C1(KEYINPUT49), .C2(new_n835), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n868), .A2(new_n287), .A3(new_n668), .A4(new_n674), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n866), .A2(new_n869), .ZN(G75));
  NAND2_X1  g684(.A1(new_n813), .A2(new_n814), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n871), .A2(new_n192), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(G210), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT56), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n320), .B(new_n325), .Z(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT55), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n873), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n876), .B1(new_n873), .B2(new_n874), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n384), .A2(G952), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT119), .Z(new_n880));
  NOR3_X1   g694(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(G51));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n871), .A2(new_n192), .A3(new_n745), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n193), .B(KEYINPUT57), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n813), .A2(KEYINPUT54), .A3(new_n814), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n884), .B1(new_n885), .B2(new_n815), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n883), .B1(new_n886), .B2(new_n682), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n882), .B1(new_n887), .B2(new_n879), .ZN(new_n888));
  INV_X1    g702(.A(new_n879), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT54), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n871), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n813), .A2(KEYINPUT54), .A3(new_n814), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n683), .B1(new_n893), .B2(new_n884), .ZN(new_n894));
  OAI211_X1 g708(.A(KEYINPUT120), .B(new_n889), .C1(new_n894), .C2(new_n883), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n888), .A2(new_n895), .ZN(G54));
  NAND3_X1  g710(.A1(new_n872), .A2(KEYINPUT58), .A3(G475), .ZN(new_n897));
  INV_X1    g711(.A(new_n443), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n900), .A3(new_n879), .ZN(G60));
  NAND2_X1  g715(.A1(G478), .A2(G902), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT59), .Z(new_n903));
  OAI211_X1 g717(.A(new_n592), .B(new_n591), .C1(new_n822), .C2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n880), .ZN(new_n905));
  INV_X1    g719(.A(new_n903), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n893), .A2(new_n593), .A3(new_n906), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(G63));
  NAND2_X1  g722(.A1(new_n553), .A2(new_n554), .ZN(new_n909));
  NAND2_X1  g723(.A1(G217), .A2(G902), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT121), .Z(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT60), .Z(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n909), .B1(new_n871), .B2(new_n913), .ZN(new_n914));
  OR2_X1    g728(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n813), .A2(new_n628), .A3(new_n814), .A4(new_n912), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n914), .A2(new_n905), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(G66));
  OAI21_X1  g733(.A(G953), .B1(new_n388), .B2(new_n323), .ZN(new_n920));
  NOR4_X1   g734(.A1(new_n783), .A2(new_n803), .A3(new_n583), .A4(new_n635), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n920), .B1(new_n921), .B2(G953), .ZN(new_n922));
  INV_X1    g736(.A(new_n320), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n923), .B1(G898), .B2(new_n384), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n922), .B(new_n924), .ZN(G69));
  NAND2_X1  g739(.A1(new_n395), .A2(new_n398), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n515), .B(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n928), .A2(G900), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT124), .B1(new_n929), .B2(G953), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n270), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  AOI211_X1 g746(.A(new_n384), .B(new_n930), .C1(G900), .C2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n384), .B1(new_n932), .B2(G900), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n786), .A2(new_n654), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n935), .A2(new_n675), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT62), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n567), .A2(new_n582), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n800), .A2(new_n801), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n938), .A2(new_n939), .A3(new_n660), .A4(new_n806), .ZN(new_n940));
  AND4_X1   g754(.A1(new_n766), .A2(new_n937), .A3(new_n773), .A4(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(G953), .B1(new_n941), .B2(new_n927), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n766), .A2(new_n654), .A3(new_n786), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(KEYINPUT123), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT123), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n766), .A2(new_n945), .A3(new_n654), .A4(new_n786), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n755), .A2(new_n580), .A3(new_n778), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n773), .A2(new_n733), .A3(new_n738), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n928), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n934), .B1(new_n942), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n933), .B1(new_n952), .B2(new_n930), .ZN(G72));
  NAND2_X1  g767(.A1(new_n941), .A2(new_n921), .ZN(new_n954));
  NAND2_X1  g768(.A1(G472), .A2(G902), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT63), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT125), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n958), .A2(new_n469), .A3(new_n495), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n947), .A2(new_n921), .A3(new_n949), .A4(new_n948), .ZN(new_n960));
  AOI211_X1 g774(.A(new_n469), .B(new_n495), .C1(new_n960), .C2(new_n957), .ZN(new_n961));
  OAI21_X1  g775(.A(KEYINPUT126), .B1(new_n961), .B2(new_n879), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n957), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n963), .A2(new_n471), .A3(new_n516), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT126), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n964), .A2(new_n965), .A3(new_n889), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n508), .A2(KEYINPUT127), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n956), .B1(new_n967), .B2(new_n496), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n821), .B(new_n968), .C1(new_n496), .C2(new_n967), .ZN(new_n969));
  AND4_X1   g783(.A1(new_n959), .A2(new_n962), .A3(new_n966), .A4(new_n969), .ZN(G57));
endmodule


