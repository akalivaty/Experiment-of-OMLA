

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582;

  NOR2_X1 U323 ( .A1(n515), .A2(n412), .ZN(n567) );
  XNOR2_X1 U324 ( .A(n442), .B(n441), .ZN(n530) );
  INV_X1 U325 ( .A(KEYINPUT112), .ZN(n358) );
  XNOR2_X1 U326 ( .A(n358), .B(KEYINPUT46), .ZN(n359) );
  XNOR2_X1 U327 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U328 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n391) );
  XNOR2_X1 U329 ( .A(n392), .B(n391), .ZN(n528) );
  XNOR2_X1 U330 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U331 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U332 ( .A(KEYINPUT37), .B(KEYINPUT101), .ZN(n464) );
  XNOR2_X1 U333 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U334 ( .A(n356), .B(n355), .ZN(n572) );
  XNOR2_X1 U335 ( .A(n465), .B(n464), .ZN(n514) );
  XNOR2_X1 U336 ( .A(n467), .B(n466), .ZN(n497) );
  XNOR2_X1 U337 ( .A(G169GAT), .B(KEYINPUT124), .ZN(n445) );
  XNOR2_X1 U338 ( .A(n468), .B(G43GAT), .ZN(n469) );
  XNOR2_X1 U339 ( .A(n446), .B(n445), .ZN(G1348GAT) );
  XNOR2_X1 U340 ( .A(n470), .B(n469), .ZN(G1330GAT) );
  XNOR2_X1 U341 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n291) );
  XNOR2_X1 U342 ( .A(n291), .B(KEYINPUT7), .ZN(n377) );
  XOR2_X1 U343 ( .A(G50GAT), .B(G22GAT), .Z(n292) );
  XOR2_X1 U344 ( .A(G141GAT), .B(n292), .Z(n414) );
  XOR2_X1 U345 ( .A(n377), .B(n414), .Z(n305) );
  XOR2_X1 U346 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n294) );
  XNOR2_X1 U347 ( .A(KEYINPUT69), .B(KEYINPUT67), .ZN(n293) );
  XNOR2_X1 U348 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U349 ( .A(G15GAT), .B(KEYINPUT30), .Z(n296) );
  NAND2_X1 U350 ( .A1(G229GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U351 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U352 ( .A(n298), .B(n297), .Z(n303) );
  XNOR2_X1 U353 ( .A(G29GAT), .B(G113GAT), .ZN(n299) );
  XNOR2_X1 U354 ( .A(n299), .B(G1GAT), .ZN(n319) );
  XOR2_X1 U355 ( .A(G8GAT), .B(G197GAT), .Z(n301) );
  XNOR2_X1 U356 ( .A(G169GAT), .B(G36GAT), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n405) );
  XNOR2_X1 U358 ( .A(n319), .B(n405), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U360 ( .A(n305), .B(n304), .ZN(n568) );
  XNOR2_X1 U361 ( .A(KEYINPUT70), .B(n568), .ZN(n535) );
  XOR2_X1 U362 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n307) );
  XNOR2_X1 U363 ( .A(KEYINPUT4), .B(KEYINPUT88), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n323) );
  XOR2_X1 U365 ( .A(G120GAT), .B(G57GAT), .Z(n340) );
  XOR2_X1 U366 ( .A(KEYINPUT1), .B(KEYINPUT87), .Z(n309) );
  XNOR2_X1 U367 ( .A(G141GAT), .B(G85GAT), .ZN(n308) );
  XNOR2_X1 U368 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U369 ( .A(n340), .B(n310), .Z(n312) );
  NAND2_X1 U370 ( .A1(G225GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U371 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U372 ( .A(KEYINPUT2), .B(G162GAT), .Z(n314) );
  XNOR2_X1 U373 ( .A(G155GAT), .B(G148GAT), .ZN(n313) );
  XNOR2_X1 U374 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U375 ( .A(KEYINPUT3), .B(n315), .Z(n421) );
  XOR2_X1 U376 ( .A(n316), .B(n421), .Z(n321) );
  XOR2_X1 U377 ( .A(G127GAT), .B(KEYINPUT81), .Z(n318) );
  XNOR2_X1 U378 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n317) );
  XNOR2_X1 U379 ( .A(n318), .B(n317), .ZN(n430) );
  XNOR2_X1 U380 ( .A(n319), .B(n430), .ZN(n320) );
  XNOR2_X1 U381 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U382 ( .A(n323), .B(n322), .Z(n454) );
  XNOR2_X1 U383 ( .A(KEYINPUT89), .B(n454), .ZN(n515) );
  XOR2_X1 U384 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n325) );
  XNOR2_X1 U385 ( .A(G8GAT), .B(KEYINPUT80), .ZN(n324) );
  XNOR2_X1 U386 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U387 ( .A(G71GAT), .B(KEYINPUT13), .Z(n341) );
  XOR2_X1 U388 ( .A(KEYINPUT15), .B(n341), .Z(n327) );
  XNOR2_X1 U389 ( .A(G211GAT), .B(G155GAT), .ZN(n326) );
  XNOR2_X1 U390 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U391 ( .A(n329), .B(n328), .Z(n331) );
  NAND2_X1 U392 ( .A1(G231GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U393 ( .A(n331), .B(n330), .ZN(n339) );
  XOR2_X1 U394 ( .A(G78GAT), .B(G127GAT), .Z(n333) );
  XNOR2_X1 U395 ( .A(G22GAT), .B(G183GAT), .ZN(n332) );
  XNOR2_X1 U396 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U397 ( .A(G64GAT), .B(G57GAT), .Z(n335) );
  XNOR2_X1 U398 ( .A(G1GAT), .B(G15GAT), .ZN(n334) );
  XNOR2_X1 U399 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U400 ( .A(n337), .B(n336), .Z(n338) );
  XNOR2_X1 U401 ( .A(n339), .B(n338), .ZN(n577) );
  XNOR2_X1 U402 ( .A(n341), .B(n340), .ZN(n343) );
  AND2_X1 U403 ( .A1(G230GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U405 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n345) );
  XNOR2_X1 U406 ( .A(KEYINPUT74), .B(KEYINPUT32), .ZN(n344) );
  XOR2_X1 U407 ( .A(n345), .B(n344), .Z(n346) );
  XNOR2_X1 U408 ( .A(n347), .B(n346), .ZN(n356) );
  XNOR2_X1 U409 ( .A(G99GAT), .B(G85GAT), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n348), .B(KEYINPUT71), .ZN(n376) );
  XNOR2_X1 U411 ( .A(G176GAT), .B(G92GAT), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n349), .B(G64GAT), .ZN(n404) );
  XNOR2_X1 U413 ( .A(n376), .B(n404), .ZN(n354) );
  XOR2_X1 U414 ( .A(G106GAT), .B(G78GAT), .Z(n413) );
  XOR2_X1 U415 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n351) );
  XNOR2_X1 U416 ( .A(G204GAT), .B(G148GAT), .ZN(n350) );
  XNOR2_X1 U417 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U418 ( .A(n413), .B(n352), .ZN(n353) );
  INV_X1 U419 ( .A(KEYINPUT41), .ZN(n357) );
  XNOR2_X1 U420 ( .A(n572), .B(n357), .ZN(n499) );
  INV_X1 U421 ( .A(n499), .ZN(n559) );
  NAND2_X1 U422 ( .A1(n559), .A2(n568), .ZN(n360) );
  NOR2_X1 U423 ( .A1(n577), .A2(n361), .ZN(n384) );
  NAND2_X1 U424 ( .A1(G232GAT), .A2(G233GAT), .ZN(n367) );
  XOR2_X1 U425 ( .A(KEYINPUT65), .B(G106GAT), .Z(n363) );
  XNOR2_X1 U426 ( .A(G50GAT), .B(G29GAT), .ZN(n362) );
  XNOR2_X1 U427 ( .A(n363), .B(n362), .ZN(n365) );
  XOR2_X1 U428 ( .A(G36GAT), .B(G218GAT), .Z(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U430 ( .A(n367), .B(n366), .ZN(n383) );
  XOR2_X1 U431 ( .A(KEYINPUT11), .B(KEYINPUT77), .Z(n369) );
  XNOR2_X1 U432 ( .A(KEYINPUT79), .B(KEYINPUT66), .ZN(n368) );
  XNOR2_X1 U433 ( .A(n369), .B(n368), .ZN(n381) );
  XOR2_X1 U434 ( .A(KEYINPUT78), .B(KEYINPUT10), .Z(n371) );
  XNOR2_X1 U435 ( .A(G162GAT), .B(KEYINPUT9), .ZN(n370) );
  XNOR2_X1 U436 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U437 ( .A(G92GAT), .B(KEYINPUT76), .Z(n373) );
  XNOR2_X1 U438 ( .A(G190GAT), .B(G134GAT), .ZN(n372) );
  XNOR2_X1 U439 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U440 ( .A(n375), .B(n374), .Z(n379) );
  XNOR2_X1 U441 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U443 ( .A(n381), .B(n380), .Z(n382) );
  XNOR2_X1 U444 ( .A(n383), .B(n382), .ZN(n471) );
  NAND2_X1 U445 ( .A1(n384), .A2(n471), .ZN(n385) );
  XNOR2_X1 U446 ( .A(n385), .B(KEYINPUT47), .ZN(n390) );
  INV_X1 U447 ( .A(n577), .ZN(n476) );
  XNOR2_X1 U448 ( .A(KEYINPUT36), .B(n471), .ZN(n580) );
  NOR2_X1 U449 ( .A1(n476), .A2(n580), .ZN(n386) );
  XNOR2_X1 U450 ( .A(KEYINPUT45), .B(n386), .ZN(n387) );
  NAND2_X1 U451 ( .A1(n387), .A2(n572), .ZN(n388) );
  NOR2_X1 U452 ( .A1(n388), .A2(n535), .ZN(n389) );
  NOR2_X1 U453 ( .A1(n390), .A2(n389), .ZN(n392) );
  XNOR2_X1 U454 ( .A(KEYINPUT85), .B(KEYINPUT18), .ZN(n393) );
  XNOR2_X1 U455 ( .A(n393), .B(KEYINPUT17), .ZN(n394) );
  XOR2_X1 U456 ( .A(n394), .B(KEYINPUT19), .Z(n396) );
  XNOR2_X1 U457 ( .A(G183GAT), .B(G190GAT), .ZN(n395) );
  XNOR2_X1 U458 ( .A(n396), .B(n395), .ZN(n432) );
  XOR2_X1 U459 ( .A(KEYINPUT86), .B(G218GAT), .Z(n398) );
  XNOR2_X1 U460 ( .A(G211GAT), .B(G204GAT), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U462 ( .A(KEYINPUT21), .B(n399), .ZN(n424) );
  INV_X1 U463 ( .A(n424), .ZN(n400) );
  XNOR2_X1 U464 ( .A(n432), .B(n400), .ZN(n409) );
  XOR2_X1 U465 ( .A(KEYINPUT90), .B(KEYINPUT92), .Z(n402) );
  NAND2_X1 U466 ( .A1(G226GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U467 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U468 ( .A(n403), .B(KEYINPUT91), .Z(n407) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U470 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n409), .B(n408), .ZN(n517) );
  XOR2_X1 U472 ( .A(KEYINPUT122), .B(n517), .Z(n410) );
  NOR2_X1 U473 ( .A1(n528), .A2(n410), .ZN(n411) );
  XOR2_X1 U474 ( .A(KEYINPUT54), .B(n411), .Z(n412) );
  XOR2_X1 U475 ( .A(n413), .B(KEYINPUT23), .Z(n416) );
  XNOR2_X1 U476 ( .A(n414), .B(KEYINPUT76), .ZN(n415) );
  XNOR2_X1 U477 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U478 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n418) );
  NAND2_X1 U479 ( .A1(G228GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U481 ( .A(n420), .B(n419), .Z(n423) );
  XNOR2_X1 U482 ( .A(G197GAT), .B(n421), .ZN(n422) );
  XNOR2_X1 U483 ( .A(n423), .B(n422), .ZN(n425) );
  XNOR2_X1 U484 ( .A(n425), .B(n424), .ZN(n456) );
  NAND2_X1 U485 ( .A1(n567), .A2(n456), .ZN(n426) );
  XNOR2_X1 U486 ( .A(n426), .B(KEYINPUT55), .ZN(n443) );
  XOR2_X1 U487 ( .A(KEYINPUT83), .B(G120GAT), .Z(n428) );
  XNOR2_X1 U488 ( .A(G113GAT), .B(G15GAT), .ZN(n427) );
  XNOR2_X1 U489 ( .A(n428), .B(n427), .ZN(n434) );
  XOR2_X1 U490 ( .A(G71GAT), .B(KEYINPUT82), .Z(n429) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n442) );
  NAND2_X1 U492 ( .A1(G227GAT), .A2(G233GAT), .ZN(n440) );
  XOR2_X1 U493 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n436) );
  XNOR2_X1 U494 ( .A(G169GAT), .B(G176GAT), .ZN(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n438) );
  XOR2_X1 U496 ( .A(G43GAT), .B(G99GAT), .Z(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U498 ( .A(n440), .B(n439), .ZN(n441) );
  NAND2_X1 U499 ( .A1(n443), .A2(n530), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n444), .B(KEYINPUT123), .ZN(n564) );
  NAND2_X1 U501 ( .A1(n535), .A2(n564), .ZN(n446) );
  XOR2_X1 U502 ( .A(KEYINPUT38), .B(KEYINPUT102), .Z(n467) );
  NAND2_X1 U503 ( .A1(n572), .A2(n535), .ZN(n447) );
  XNOR2_X1 U504 ( .A(n447), .B(KEYINPUT75), .ZN(n481) );
  INV_X1 U505 ( .A(KEYINPUT100), .ZN(n462) );
  NAND2_X1 U506 ( .A1(n517), .A2(n530), .ZN(n448) );
  NAND2_X1 U507 ( .A1(n456), .A2(n448), .ZN(n449) );
  XOR2_X1 U508 ( .A(KEYINPUT25), .B(n449), .Z(n452) );
  XNOR2_X1 U509 ( .A(n517), .B(KEYINPUT27), .ZN(n455) );
  NOR2_X1 U510 ( .A1(n530), .A2(n456), .ZN(n450) );
  XNOR2_X1 U511 ( .A(n450), .B(KEYINPUT26), .ZN(n566) );
  NAND2_X1 U512 ( .A1(n455), .A2(n566), .ZN(n451) );
  NAND2_X1 U513 ( .A1(n452), .A2(n451), .ZN(n453) );
  NAND2_X1 U514 ( .A1(n454), .A2(n453), .ZN(n459) );
  NAND2_X1 U515 ( .A1(n515), .A2(n455), .ZN(n527) );
  NOR2_X1 U516 ( .A1(n530), .A2(n527), .ZN(n457) );
  XNOR2_X1 U517 ( .A(n456), .B(KEYINPUT28), .ZN(n533) );
  NAND2_X1 U518 ( .A1(n457), .A2(n533), .ZN(n458) );
  NAND2_X1 U519 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U520 ( .A(KEYINPUT93), .B(n460), .ZN(n479) );
  NOR2_X1 U521 ( .A1(n479), .A2(n577), .ZN(n461) );
  XNOR2_X1 U522 ( .A(n462), .B(n461), .ZN(n463) );
  NOR2_X1 U523 ( .A1(n580), .A2(n463), .ZN(n465) );
  NAND2_X1 U524 ( .A1(n481), .A2(n514), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n497), .A2(n530), .ZN(n470) );
  XOR2_X1 U526 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n468) );
  INV_X1 U527 ( .A(G190GAT), .ZN(n475) );
  XOR2_X1 U528 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n473) );
  INV_X1 U529 ( .A(n471), .ZN(n555) );
  NAND2_X1 U530 ( .A1(n564), .A2(n555), .ZN(n472) );
  XNOR2_X1 U531 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n475), .B(n474), .ZN(G1351GAT) );
  XOR2_X1 U533 ( .A(KEYINPUT96), .B(KEYINPUT34), .Z(n484) );
  NOR2_X1 U534 ( .A1(n476), .A2(n555), .ZN(n477) );
  XOR2_X1 U535 ( .A(KEYINPUT16), .B(n477), .Z(n478) );
  NOR2_X1 U536 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U537 ( .A(KEYINPUT94), .B(n480), .ZN(n500) );
  NAND2_X1 U538 ( .A1(n500), .A2(n481), .ZN(n482) );
  XNOR2_X1 U539 ( .A(n482), .B(KEYINPUT95), .ZN(n491) );
  NAND2_X1 U540 ( .A1(n491), .A2(n515), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U542 ( .A(G1GAT), .B(n485), .Z(G1324GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n487) );
  NAND2_X1 U544 ( .A1(n491), .A2(n517), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U546 ( .A(G8GAT), .B(n488), .ZN(G1325GAT) );
  XOR2_X1 U547 ( .A(G15GAT), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U548 ( .A1(n491), .A2(n530), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  XOR2_X1 U550 ( .A(G22GAT), .B(KEYINPUT99), .Z(n493) );
  INV_X1 U551 ( .A(n533), .ZN(n521) );
  NAND2_X1 U552 ( .A1(n491), .A2(n521), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(G1327GAT) );
  XOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT39), .Z(n495) );
  NAND2_X1 U555 ( .A1(n497), .A2(n515), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(G1328GAT) );
  NAND2_X1 U557 ( .A1(n497), .A2(n517), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n496), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U559 ( .A1(n521), .A2(n497), .ZN(n498) );
  XNOR2_X1 U560 ( .A(G50GAT), .B(n498), .ZN(G1331GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n503) );
  NOR2_X1 U562 ( .A1(n499), .A2(n568), .ZN(n513) );
  NAND2_X1 U563 ( .A1(n500), .A2(n513), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n501), .B(KEYINPUT105), .ZN(n508) );
  NAND2_X1 U565 ( .A1(n508), .A2(n515), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U567 ( .A(G57GAT), .B(n504), .Z(G1332GAT) );
  NAND2_X1 U568 ( .A1(n508), .A2(n517), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n505), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U570 ( .A1(n530), .A2(n508), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n506), .B(KEYINPUT106), .ZN(n507) );
  XNOR2_X1 U572 ( .A(G71GAT), .B(n507), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U574 ( .A1(n508), .A2(n521), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(n512) );
  XOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT108), .Z(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  AND2_X1 U578 ( .A1(n514), .A2(n513), .ZN(n522) );
  NAND2_X1 U579 ( .A1(n522), .A2(n515), .ZN(n516) );
  XNOR2_X1 U580 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  NAND2_X1 U581 ( .A1(n522), .A2(n517), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n518), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U583 ( .A(G99GAT), .B(KEYINPUT109), .Z(n520) );
  NAND2_X1 U584 ( .A1(n522), .A2(n530), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(G1338GAT) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(KEYINPUT110), .ZN(n526) );
  XOR2_X1 U587 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n524) );
  NAND2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(G1339GAT) );
  NOR2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U592 ( .A(KEYINPUT113), .B(n529), .Z(n547) );
  NAND2_X1 U593 ( .A1(n547), .A2(n530), .ZN(n531) );
  XOR2_X1 U594 ( .A(KEYINPUT114), .B(n531), .Z(n532) );
  NAND2_X1 U595 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U596 ( .A(n534), .B(KEYINPUT115), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n543), .A2(n535), .ZN(n536) );
  XNOR2_X1 U598 ( .A(n536), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n538) );
  NAND2_X1 U600 ( .A1(n543), .A2(n559), .ZN(n537) );
  XNOR2_X1 U601 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U602 ( .A(G120GAT), .B(n539), .ZN(G1341GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n541) );
  NAND2_X1 U604 ( .A1(n543), .A2(n577), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U608 ( .A1(n543), .A2(n555), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(n546), .ZN(G1343GAT) );
  XOR2_X1 U611 ( .A(G141GAT), .B(KEYINPUT119), .Z(n549) );
  AND2_X1 U612 ( .A1(n547), .A2(n566), .ZN(n556) );
  NAND2_X1 U613 ( .A1(n556), .A2(n568), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(G1344GAT) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n553) );
  XOR2_X1 U616 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n551) );
  NAND2_X1 U617 ( .A1(n556), .A2(n559), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  NAND2_X1 U620 ( .A1(n577), .A2(n556), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U622 ( .A(G162GAT), .B(KEYINPUT121), .Z(n558) );
  NAND2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1347GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n561) );
  NAND2_X1 U626 ( .A1(n564), .A2(n559), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n563) );
  XOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT56), .Z(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  NAND2_X1 U630 ( .A1(n577), .A2(n564), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n570) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n579) );
  INV_X1 U634 ( .A(n579), .ZN(n576) );
  NAND2_X1 U635 ( .A1(n576), .A2(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n574) );
  OR2_X1 U639 ( .A1(n579), .A2(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U641 ( .A(G204GAT), .B(n575), .Z(G1353GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(KEYINPUT62), .B(n581), .Z(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

