//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n624, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1157;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT66), .Z(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  XNOR2_X1  g029(.A(G325), .B(KEYINPUT67), .ZN(G261));
  NAND2_X1  g030(.A1(new_n453), .A2(G567), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n456), .A2(KEYINPUT68), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(KEYINPUT68), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n451), .A2(G2106), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n469), .B1(new_n462), .B2(new_n463), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n469), .A2(G2104), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n471), .A2(G137), .B1(G101), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(G160));
  NOR2_X1   g049(.A1(new_n464), .A2(new_n469), .ZN(new_n475));
  AOI22_X1  g050(.A1(G124), .A2(new_n475), .B1(new_n471), .B2(G136), .ZN(new_n476));
  NOR2_X1   g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT69), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n476), .A2(new_n479), .ZN(G162));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(G138), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(KEYINPUT70), .B2(KEYINPUT4), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n471), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n475), .A2(G126), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n481), .B(new_n482), .C1(new_n470), .C2(new_n484), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G114), .C2(new_n469), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n486), .A2(new_n487), .A3(new_n488), .A4(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G164));
  NOR2_X1   g067(.A1(KEYINPUT6), .A2(G651), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  XNOR2_X1  g069(.A(KEYINPUT71), .B(G651), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT6), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT73), .B1(new_n498), .B2(KEYINPUT5), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT73), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(new_n501), .A3(G543), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n503), .B1(new_n501), .B2(G543), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n498), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n499), .A2(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n497), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n497), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n506), .A2(G62), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n495), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT74), .ZN(new_n515));
  OR3_X1    g090(.A1(new_n511), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n511), .B2(new_n514), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(G166));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT71), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n493), .B1(new_n523), .B2(KEYINPUT6), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n524), .A2(new_n498), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XOR2_X1   g102(.A(new_n527), .B(KEYINPUT7), .Z(new_n528));
  AND2_X1   g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n528), .B1(new_n506), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n497), .A2(new_n506), .A3(G89), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n526), .A2(new_n530), .A3(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  XOR2_X1   g108(.A(KEYINPUT75), .B(G90), .Z(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n507), .A2(new_n534), .B1(new_n509), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n495), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n536), .A2(new_n538), .ZN(G171));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n499), .A2(new_n502), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n504), .A2(new_n505), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n540), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(new_n523), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n525), .A2(G43), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n497), .A2(new_n506), .A3(G81), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  OAI21_X1  g130(.A(KEYINPUT76), .B1(new_n543), .B2(new_n524), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT76), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n497), .A2(new_n506), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n556), .A2(G91), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n496), .B1(new_n520), .B2(new_n522), .ZN(new_n560));
  OAI211_X1 g135(.A(G53), .B(G543), .C1(new_n560), .C2(new_n493), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n497), .A2(new_n563), .A3(G53), .A4(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n541), .A2(new_n542), .A3(G65), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g143(.A(KEYINPUT77), .B1(new_n568), .B2(G651), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n570));
  AOI211_X1 g145(.A(new_n570), .B(new_n519), .C1(new_n566), .C2(new_n567), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n559), .B(new_n565), .C1(new_n569), .C2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT78), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n570), .B1(new_n575), .B2(new_n519), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n568), .A2(KEYINPUT77), .A3(G651), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n578), .A2(KEYINPUT78), .A3(new_n559), .A4(new_n565), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G299));
  INV_X1    g156(.A(G171), .ZN(G301));
  AND2_X1   g157(.A1(new_n516), .A2(new_n517), .ZN(G303));
  NAND2_X1  g158(.A1(new_n556), .A2(new_n558), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n585), .A2(KEYINPUT79), .A3(G87), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n587));
  INV_X1    g162(.A(G87), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n506), .A2(G74), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(new_n525), .B2(G49), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n590), .A2(new_n592), .ZN(G288));
  NAND2_X1  g168(.A1(new_n585), .A2(G86), .ZN(new_n594));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G61), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n543), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(new_n523), .B1(new_n525), .B2(G48), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n594), .A2(new_n598), .ZN(G305));
  INV_X1    g174(.A(G85), .ZN(new_n600));
  INV_X1    g175(.A(G47), .ZN(new_n601));
  OAI22_X1  g176(.A1(new_n507), .A2(new_n600), .B1(new_n509), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(new_n495), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G290));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NOR2_X1   g182(.A1(G171), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT80), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n543), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G651), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n525), .A2(G54), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n556), .A2(G92), .A3(new_n558), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g193(.A1(new_n556), .A2(KEYINPUT10), .A3(G92), .A4(new_n558), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n615), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n609), .B1(G868), .B2(new_n620), .ZN(G284));
  XNOR2_X1  g196(.A(G284), .B(KEYINPUT81), .ZN(G321));
  NOR2_X1   g197(.A1(G286), .A2(new_n607), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n580), .B(KEYINPUT82), .Z(new_n624));
  AOI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(new_n607), .ZN(G297));
  AOI21_X1  g200(.A(new_n623), .B1(new_n624), .B2(new_n607), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n620), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n549), .A2(new_n607), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n618), .A2(new_n619), .ZN(new_n630));
  INV_X1    g205(.A(new_n615), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n632), .A2(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n629), .B1(new_n633), .B2(new_n607), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g210(.A1(new_n469), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT83), .B(KEYINPUT13), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G2100), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT84), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n475), .A2(G123), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n471), .A2(G135), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n469), .A2(G111), .ZN(new_n644));
  OAI21_X1  g219(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n642), .B(new_n643), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2096), .Z(new_n647));
  OAI211_X1 g222(.A(new_n641), .B(new_n647), .C1(G2100), .C2(new_n639), .ZN(G156));
  INV_X1    g223(.A(KEYINPUT14), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2430), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n652), .B2(new_n651), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n654), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(G14), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT85), .Z(G401));
  INV_X1    g239(.A(KEYINPUT18), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n666), .A2(new_n667), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2100), .ZN(new_n672));
  XOR2_X1   g247(.A(G2072), .B(G2078), .Z(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n668), .B2(KEYINPUT18), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2096), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n672), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1956), .B(G2474), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1961), .B(G1966), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n678), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n678), .A2(new_n681), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT20), .Z(new_n685));
  AOI211_X1 g260(.A(new_n683), .B(new_n685), .C1(new_n678), .C2(new_n682), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT86), .ZN(new_n687));
  XOR2_X1   g262(.A(G1981), .B(G1986), .Z(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n687), .B(new_n692), .ZN(G229));
  NOR2_X1   g268(.A1(G16), .A2(G24), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n605), .B2(G16), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT89), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT90), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n698), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n475), .A2(G119), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n471), .A2(G131), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n469), .A2(G107), .ZN(new_n703));
  OAI21_X1  g278(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n701), .B(new_n702), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  MUX2_X1   g280(.A(G25), .B(new_n705), .S(G29), .Z(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT35), .B(G1991), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT87), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT88), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n706), .B(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n710), .A2(KEYINPUT91), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n699), .A2(new_n700), .A3(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G23), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n590), .A2(new_n592), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n713), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT33), .B(G1976), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(G16), .A2(G22), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G166), .B2(G16), .ZN(new_n720));
  INV_X1    g295(.A(G1971), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n713), .A2(G6), .ZN(new_n723));
  INV_X1    g298(.A(G305), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(new_n713), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT32), .B(G1981), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n718), .A2(new_n722), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n712), .B1(new_n728), .B2(KEYINPUT34), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT34), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n718), .A2(new_n722), .A3(new_n730), .A4(new_n727), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT36), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT93), .B(KEYINPUT25), .Z(new_n735));
  NAND3_X1  g310(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G127), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n464), .A2(new_n738), .ZN(new_n739));
  AND2_X1   g314(.A1(G115), .A2(G2104), .ZN(new_n740));
  OAI21_X1  g315(.A(G2105), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n471), .A2(G139), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n737), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT94), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G29), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT95), .ZN(new_n746));
  NOR2_X1   g321(.A1(G29), .A2(G33), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT92), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n746), .B1(new_n745), .B2(new_n748), .ZN(new_n751));
  OAI21_X1  g326(.A(G2072), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(new_n751), .ZN(new_n753));
  INV_X1    g328(.A(G2072), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n753), .A2(new_n754), .A3(new_n749), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G29), .ZN(new_n757));
  NOR2_X1   g332(.A1(G164), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G27), .B2(new_n757), .ZN(new_n759));
  INV_X1    g334(.A(G2078), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G34), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n762), .A2(KEYINPUT24), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(KEYINPUT24), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n757), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G160), .B2(new_n757), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G2084), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n761), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(G5), .A2(G16), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT97), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G301), .B2(new_n713), .ZN(new_n771));
  INV_X1    g346(.A(G1961), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n768), .A2(new_n773), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n757), .A2(G32), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n471), .A2(G141), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT96), .Z(new_n777));
  AND2_X1   g352(.A1(new_n472), .A2(G105), .ZN(new_n778));
  NAND3_X1  g353(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT26), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n778), .B(new_n780), .C1(G129), .C2(new_n475), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n775), .B1(new_n782), .B2(G29), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT27), .B(G1996), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n759), .A2(new_n760), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n783), .A2(new_n784), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n774), .A2(new_n788), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n756), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT100), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n771), .A2(new_n772), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT98), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT31), .B(G11), .Z(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT30), .B(G28), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n795), .B1(new_n757), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n713), .A2(G21), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G286), .B2(G16), .ZN(new_n799));
  INV_X1    g374(.A(G1966), .ZN(new_n800));
  OAI221_X1 g375(.A(new_n797), .B1(new_n757), .B2(new_n646), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n800), .B2(new_n799), .ZN(new_n802));
  AOI21_X1  g377(.A(KEYINPUT99), .B1(new_n794), .B2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n794), .A2(KEYINPUT99), .A3(new_n802), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n790), .A2(new_n791), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n756), .A2(new_n805), .A3(new_n789), .ZN(new_n807));
  OAI21_X1  g382(.A(KEYINPUT100), .B1(new_n807), .B2(new_n803), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n713), .A2(G20), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT23), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n580), .B2(new_n713), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G1956), .ZN(new_n812));
  NOR2_X1   g387(.A1(G16), .A2(G19), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n550), .B2(G16), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(G1341), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n757), .A2(G35), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT101), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G162), .B2(new_n757), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT29), .B(G2090), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n757), .A2(G26), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT28), .Z(new_n822));
  NAND2_X1  g397(.A1(new_n475), .A2(G128), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n471), .A2(G140), .ZN(new_n824));
  OR2_X1    g399(.A1(G104), .A2(G2105), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n825), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n823), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n822), .B1(new_n827), .B2(G29), .ZN(new_n828));
  INV_X1    g403(.A(G2067), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n820), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(G4), .A2(G16), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n620), .B2(G16), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n815), .B(new_n831), .C1(G1348), .C2(new_n833), .ZN(new_n834));
  AOI211_X1 g409(.A(new_n812), .B(new_n834), .C1(G1348), .C2(new_n833), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n806), .A2(new_n808), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(KEYINPUT36), .B1(new_n729), .B2(new_n731), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT102), .ZN(new_n838));
  NOR4_X1   g413(.A1(new_n734), .A2(new_n836), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n836), .A2(new_n837), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n729), .A2(KEYINPUT36), .A3(new_n731), .ZN(new_n841));
  AOI21_X1  g416(.A(KEYINPUT102), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n839), .A2(new_n842), .ZN(G311));
  NAND2_X1  g418(.A1(new_n840), .A2(new_n841), .ZN(G150));
  INV_X1    g419(.A(G93), .ZN(new_n845));
  INV_X1    g420(.A(G55), .ZN(new_n846));
  OAI22_X1  g421(.A1(new_n507), .A2(new_n845), .B1(new_n509), .B2(new_n846), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n848), .A2(new_n495), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(G860), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT37), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n620), .A2(G559), .ZN(new_n854));
  XOR2_X1   g429(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n847), .A2(new_n849), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(new_n549), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n550), .A2(new_n850), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n856), .B(new_n860), .Z(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n862), .A2(KEYINPUT39), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n851), .B1(new_n862), .B2(KEYINPUT39), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n853), .B1(new_n863), .B2(new_n864), .ZN(G145));
  XNOR2_X1  g440(.A(G160), .B(new_n646), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G162), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n782), .B(new_n827), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n869), .A2(new_n491), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n491), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n744), .A2(KEYINPUT104), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n744), .A2(KEYINPUT104), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n705), .B(new_n637), .Z(new_n876));
  AOI22_X1  g451(.A1(G130), .A2(new_n475), .B1(new_n471), .B2(G142), .ZN(new_n877));
  OAI21_X1  g452(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n878));
  INV_X1    g453(.A(G118), .ZN(new_n879));
  AOI22_X1  g454(.A1(new_n878), .A2(KEYINPUT105), .B1(new_n879), .B2(G2105), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(KEYINPUT105), .B2(new_n878), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n876), .B(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n875), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n875), .A2(new_n883), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n868), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n875), .A2(new_n883), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n889), .A2(new_n867), .A3(new_n884), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT40), .ZN(G395));
  AOI21_X1  g467(.A(KEYINPUT109), .B1(new_n857), .B2(new_n607), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n633), .B(new_n860), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n574), .A2(new_n579), .A3(new_n620), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n620), .B1(new_n574), .B2(new_n579), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n559), .A2(new_n565), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT78), .B1(new_n900), .B2(new_n578), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n572), .A2(new_n573), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n632), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n574), .A2(new_n579), .A3(new_n620), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(KEYINPUT41), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n895), .B1(new_n899), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n903), .A2(new_n904), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT106), .B1(new_n907), .B2(new_n896), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n894), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT107), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n715), .A2(G305), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n516), .A2(G290), .A3(new_n517), .ZN(new_n912));
  AOI21_X1  g487(.A(G305), .B1(new_n590), .B2(new_n592), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(G166), .A2(new_n605), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n911), .A2(new_n912), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n912), .ZN(new_n917));
  NOR2_X1   g492(.A1(G288), .A2(new_n724), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n917), .B1(new_n918), .B2(new_n913), .ZN(new_n919));
  XOR2_X1   g494(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n920));
  AND3_X1   g495(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n916), .A2(new_n919), .B1(new_n922), .B2(KEYINPUT42), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n897), .A2(new_n898), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n894), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n928), .B(new_n894), .C1(new_n906), .C2(new_n908), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n910), .A2(new_n924), .A3(new_n927), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(G868), .ZN(new_n931));
  INV_X1    g506(.A(new_n894), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n897), .A2(new_n898), .A3(new_n896), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT41), .B1(new_n903), .B2(new_n904), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT106), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n895), .B1(new_n925), .B2(KEYINPUT41), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n926), .B1(new_n937), .B2(new_n928), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n924), .B1(new_n938), .B2(new_n910), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n893), .B1(new_n931), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n910), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n929), .A2(new_n927), .ZN(new_n942));
  OAI22_X1  g517(.A1(new_n941), .A2(new_n942), .B1(new_n921), .B2(new_n923), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n943), .A2(KEYINPUT109), .A3(G868), .A4(new_n930), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n940), .A2(new_n944), .ZN(G295));
  AND3_X1   g520(.A1(new_n940), .A2(KEYINPUT110), .A3(new_n944), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT110), .B1(new_n940), .B2(new_n944), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(G331));
  NAND2_X1  g523(.A1(new_n916), .A2(new_n919), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n858), .A2(G301), .A3(new_n859), .ZN(new_n950));
  AOI21_X1  g525(.A(G301), .B1(new_n858), .B2(new_n859), .ZN(new_n951));
  OAI21_X1  g526(.A(G286), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n857), .A2(new_n549), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n550), .A2(new_n850), .ZN(new_n954));
  OAI21_X1  g529(.A(G171), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n858), .A2(new_n859), .A3(G301), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(G168), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n952), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n907), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT112), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n961), .A3(new_n907), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n958), .B1(new_n899), .B2(new_n905), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n960), .B(new_n962), .C1(new_n963), .C2(KEYINPUT111), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n963), .A2(KEYINPUT111), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n949), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n957), .B(new_n952), .C1(new_n906), .C2(new_n908), .ZN(new_n968));
  INV_X1    g543(.A(new_n949), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(new_n969), .A3(new_n959), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n966), .A2(new_n967), .A3(new_n888), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n888), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n969), .B1(new_n968), .B2(new_n959), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT43), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n966), .A2(KEYINPUT43), .A3(new_n888), .A4(new_n970), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n967), .B1(new_n972), .B2(new_n973), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  MUX2_X1   g553(.A(new_n975), .B(new_n978), .S(KEYINPUT44), .Z(G397));
  NAND3_X1  g554(.A1(new_n468), .A2(new_n473), .A3(G40), .ZN(new_n980));
  INV_X1    g555(.A(G1384), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n491), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n980), .B1(new_n983), .B2(KEYINPUT45), .ZN(new_n984));
  XOR2_X1   g559(.A(KEYINPUT113), .B(KEYINPUT45), .Z(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  AOI211_X1 g561(.A(KEYINPUT114), .B(new_n986), .C1(new_n491), .C2(new_n981), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n982), .B2(new_n985), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n984), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT115), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n984), .B(new_n992), .C1(new_n987), .C2(new_n989), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(new_n721), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n982), .A2(KEYINPUT50), .ZN(new_n995));
  INV_X1    g570(.A(new_n980), .ZN(new_n996));
  XOR2_X1   g571(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n997));
  NAND3_X1  g572(.A1(new_n491), .A2(new_n981), .A3(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n995), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  OR2_X1    g574(.A1(new_n999), .A2(G2090), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n994), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT117), .ZN(new_n1002));
  NAND3_X1  g577(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1003));
  OR2_X1    g578(.A1(new_n1003), .A2(KEYINPUT118), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(KEYINPUT118), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n1006));
  INV_X1    g581(.A(G8), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1006), .B1(G166), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1004), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT117), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n994), .A2(new_n1010), .A3(new_n1000), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1002), .A2(new_n1009), .A3(G8), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n983), .A2(new_n996), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT119), .B(G8), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT120), .ZN(new_n1017));
  NOR2_X1   g592(.A1(G305), .A2(G1981), .ZN(new_n1018));
  INV_X1    g593(.A(G1981), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n497), .A2(new_n506), .A3(G86), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1019), .B1(new_n598), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1017), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1016), .B1(new_n1022), .B2(KEYINPUT49), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(KEYINPUT49), .B2(new_n1022), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1016), .B1(new_n715), .B2(G1976), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1025), .B(new_n1026), .C1(G1976), .C2(new_n715), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1024), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(G288), .A2(G1976), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1018), .B1(new_n1024), .B2(new_n1030), .ZN(new_n1031));
  OAI22_X1  g606(.A1(new_n1012), .A2(new_n1029), .B1(new_n1031), .B2(new_n1016), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n999), .A2(new_n772), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n983), .A2(new_n986), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n980), .B1(new_n982), .B2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1034), .A2(new_n1036), .A3(KEYINPUT53), .A4(new_n760), .ZN(new_n1037));
  AOI21_X1  g612(.A(G2078), .B1(new_n991), .B2(new_n993), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1033), .B(new_n1037), .C1(new_n1038), .C2(KEYINPUT53), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G171), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(G1966), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1042));
  INV_X1    g617(.A(G2084), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n995), .A2(new_n1043), .A3(new_n996), .A4(new_n998), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(G286), .B(new_n1015), .C1(new_n1042), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1042), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1007), .B1(new_n1047), .B2(new_n1044), .ZN(new_n1048));
  NOR2_X1   g623(.A1(G168), .A2(new_n1014), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1046), .B(KEYINPUT51), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1015), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1049), .A2(KEYINPUT51), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1050), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT62), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT127), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT127), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1050), .A2(new_n1057), .A3(KEYINPUT62), .A4(new_n1053), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1059));
  AND4_X1   g634(.A1(new_n1041), .A2(new_n1056), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1024), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n997), .B1(new_n491), .B2(new_n981), .ZN(new_n1062));
  OR3_X1    g637(.A1(new_n1062), .A2(KEYINPUT121), .A3(new_n980), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT121), .B1(new_n1062), .B2(new_n980), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1063), .B(new_n1064), .C1(KEYINPUT50), .C2(new_n982), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n994), .B1(G2090), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n1015), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1004), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1061), .A2(new_n1012), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1032), .B1(new_n1060), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT63), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1061), .A2(new_n1012), .A3(new_n1069), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n1051), .A2(G286), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1002), .A2(G8), .A3(new_n1011), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n1068), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1074), .A2(new_n1072), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1077), .A2(new_n1012), .A3(new_n1061), .A4(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1075), .A2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n983), .A2(new_n986), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1082), .A2(KEYINPUT53), .A3(new_n760), .A4(new_n984), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1033), .B(new_n1083), .C1(new_n1038), .C2(KEYINPUT53), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1040), .B1(G171), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1054), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT56), .B(G2072), .Z(new_n1088));
  OR2_X1    g663(.A1(new_n990), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n1090));
  INV_X1    g665(.A(G1956), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1065), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1090), .B1(new_n1065), .B2(new_n1091), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1089), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT123), .B(KEYINPUT57), .ZN(new_n1095));
  XOR2_X1   g670(.A(new_n572), .B(new_n1095), .Z(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1096), .B(new_n1089), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1099));
  INV_X1    g674(.A(G1348), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n999), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(G2067), .B2(new_n1013), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1099), .A2(new_n620), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n550), .B1(KEYINPUT125), .B2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT124), .B(G1996), .Z(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n984), .B(new_n1107), .C1(new_n987), .C2(new_n989), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT58), .B(G1341), .Z(new_n1109));
  NAND2_X1  g684(.A1(new_n1013), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1105), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1104), .A2(KEYINPUT125), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1111), .B(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1013), .A2(G2067), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(new_n1100), .B2(new_n999), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n632), .A2(KEYINPUT126), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n632), .A2(KEYINPUT126), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1115), .A2(new_n1116), .A3(KEYINPUT60), .A4(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT60), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1102), .A2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1102), .A2(new_n1119), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1118), .B(new_n1120), .C1(new_n1121), .C2(new_n1117), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1113), .B(new_n1122), .C1(new_n1099), .C2(KEYINPUT61), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1099), .A2(KEYINPUT61), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1098), .B(new_n1103), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1084), .A2(G171), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1126), .B(KEYINPUT54), .C1(G171), .C2(new_n1039), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1087), .A2(new_n1125), .A3(new_n1070), .A4(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1071), .A2(new_n1080), .A3(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1082), .A2(new_n980), .ZN(new_n1130));
  INV_X1    g705(.A(G1996), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n782), .B(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n827), .B(new_n829), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n705), .A2(new_n708), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n705), .A2(new_n708), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  XOR2_X1   g711(.A(new_n605), .B(G1986), .Z(new_n1137));
  OAI21_X1  g712(.A(new_n1130), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1129), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(KEYINPUT46), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1133), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1130), .B1(new_n782), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT47), .ZN(new_n1145));
  NOR2_X1   g720(.A1(G290), .A2(G1986), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1130), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1148), .A2(KEYINPUT48), .B1(new_n1136), .B2(new_n1130), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(KEYINPUT48), .B2(new_n1148), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1151));
  OAI22_X1  g726(.A1(new_n1151), .A2(new_n1135), .B1(G2067), .B2(new_n827), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n1130), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1145), .A2(new_n1150), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1139), .A2(new_n1154), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g730(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1157));
  NAND3_X1  g731(.A1(new_n975), .A2(new_n891), .A3(new_n1157), .ZN(G225));
  INV_X1    g732(.A(G225), .ZN(G308));
endmodule


