//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1268, new_n1269,
    new_n1270;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT0), .ZN(new_n206));
  NOR2_X1   g0006(.A1(G58), .A2(G68), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  OR2_X1    g0008(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n210));
  NAND3_X1  g0010(.A1(new_n209), .A2(G50), .A3(new_n210), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT65), .Z(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n212), .A2(G20), .A3(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G116), .ZN(new_n219));
  INV_X1    g0019(.A(G270), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT66), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AND2_X1   g0023(.A1(new_n221), .A2(new_n222), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n223), .B(new_n224), .C1(G107), .C2(G264), .ZN(new_n225));
  INV_X1    g0025(.A(G58), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  INV_X1    g0027(.A(G97), .ZN(new_n228));
  INV_X1    g0028(.A(G257), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n225), .B1(new_n226), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(G87), .ZN(new_n231));
  INV_X1    g0031(.A(G250), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n203), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n206), .B(new_n215), .C1(new_n234), .C2(KEYINPUT1), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n234), .ZN(G361));
  XNOR2_X1  g0036(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT68), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G264), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n220), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT69), .ZN(new_n248));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n250), .B(new_n253), .Z(G351));
  INV_X1    g0054(.A(G200), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G222), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G223), .A2(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(G77), .B2(new_n256), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT71), .ZN(new_n262));
  OR2_X1    g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(new_n262), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G41), .A2(G45), .ZN(new_n267));
  INV_X1    g0067(.A(G274), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n267), .A2(G1), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT70), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT70), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G1), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n267), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n264), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n269), .B1(new_n276), .B2(G226), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n255), .B1(new_n266), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n266), .A2(new_n277), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n278), .B1(G190), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G20), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n281), .B1(new_n271), .B2(new_n273), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n213), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n282), .A2(new_n217), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n281), .B1(new_n207), .B2(new_n217), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n286), .B1(G150), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT8), .B(G58), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT72), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OR3_X1    g0091(.A1(new_n290), .A2(new_n226), .A3(KEYINPUT8), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G33), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G20), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n288), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n285), .B1(new_n297), .B2(new_n284), .ZN(new_n298));
  INV_X1    g0098(.A(G13), .ZN(new_n299));
  AOI211_X1 g0099(.A(new_n299), .B(new_n281), .C1(new_n271), .C2(new_n273), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n217), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  OR2_X1    g0102(.A1(KEYINPUT77), .A2(KEYINPUT9), .ZN(new_n303));
  NAND2_X1  g0103(.A1(KEYINPUT77), .A2(KEYINPUT9), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n272), .A2(G1), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n270), .A2(KEYINPUT70), .ZN(new_n307));
  OAI211_X1 g0107(.A(G13), .B(G20), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n298), .B1(G50), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n309), .A2(KEYINPUT77), .A3(KEYINPUT9), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n280), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n280), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n218), .A2(new_n257), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n256), .B(new_n317), .C1(G232), .C2(new_n257), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT78), .B1(new_n294), .B2(new_n228), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT78), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(G33), .A3(G97), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n269), .B1(new_n323), .B2(new_n264), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT13), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n276), .A2(G238), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n325), .B1(new_n324), .B2(new_n326), .ZN(new_n328));
  OAI21_X1  g0128(.A(G200), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n324), .A2(new_n326), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT13), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(G190), .A3(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT76), .B1(new_n300), .B2(new_n284), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT76), .ZN(new_n335));
  INV_X1    g0135(.A(new_n284), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n308), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n282), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(G68), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT79), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT79), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n338), .A2(new_n342), .A3(G68), .A4(new_n339), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G68), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n300), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n346), .B(KEYINPUT12), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT11), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n295), .A2(G77), .B1(G20), .B2(new_n345), .ZN(new_n349));
  INV_X1    g0149(.A(new_n287), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(new_n217), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n348), .B1(new_n351), .B2(new_n284), .ZN(new_n352));
  AND3_X1   g0152(.A1(new_n351), .A2(new_n348), .A3(new_n284), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n347), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n329), .A2(new_n333), .A3(new_n344), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT80), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n354), .B1(new_n341), .B2(new_n343), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT80), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n358), .A2(new_n359), .A3(new_n329), .A4(new_n333), .ZN(new_n360));
  OAI21_X1  g0160(.A(G169), .B1(new_n327), .B2(new_n328), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT14), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n331), .A2(G179), .A3(new_n332), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT14), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n364), .B(G169), .C1(new_n327), .C2(new_n328), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n362), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n358), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n357), .A2(new_n360), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n309), .B1(new_n279), .B2(G169), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n369), .A2(KEYINPUT73), .ZN(new_n370));
  INV_X1    g0170(.A(G179), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n279), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(KEYINPUT73), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n370), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G238), .A2(G1698), .ZN(new_n375));
  AND2_X1   g0175(.A1(KEYINPUT3), .A2(G33), .ZN(new_n376));
  NOR2_X1   g0176(.A1(KEYINPUT3), .A2(G33), .ZN(new_n377));
  OAI221_X1 g0177(.A(new_n375), .B1(new_n227), .B2(G1698), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n378), .B(new_n264), .C1(G107), .C2(new_n256), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n276), .A2(G244), .ZN(new_n380));
  INV_X1    g0180(.A(new_n269), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G169), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n379), .A2(new_n380), .A3(new_n371), .A4(new_n381), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n338), .A2(G77), .A3(new_n339), .ZN(new_n387));
  INV_X1    g0187(.A(G77), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n300), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g0189(.A(new_n389), .B(KEYINPUT75), .ZN(new_n390));
  XOR2_X1   g0190(.A(KEYINPUT15), .B(G87), .Z(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n392), .A2(new_n296), .ZN(new_n393));
  OAI22_X1  g0193(.A1(new_n289), .A2(new_n350), .B1(new_n281), .B2(new_n388), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n284), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n387), .A2(new_n390), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n386), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n316), .A2(new_n368), .A3(new_n374), .A4(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n376), .A2(new_n377), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT7), .B1(new_n399), .B2(new_n281), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  NOR4_X1   g0201(.A1(new_n376), .A2(new_n377), .A3(new_n401), .A4(G20), .ZN(new_n402));
  OAI21_X1  g0202(.A(G68), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G58), .A2(G68), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(G20), .B1(new_n405), .B2(new_n207), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n287), .A2(G159), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT81), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n403), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n403), .A2(KEYINPUT16), .A3(new_n406), .A4(new_n408), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n284), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n293), .A2(new_n308), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n282), .A2(new_n284), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n414), .B1(new_n293), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT82), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n414), .B(KEYINPUT82), .C1(new_n293), .C2(new_n415), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n276), .A2(G232), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G41), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n214), .B1(new_n294), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n218), .A2(G1698), .ZN(new_n425));
  OAI221_X1 g0225(.A(new_n425), .B1(G223), .B2(G1698), .C1(new_n376), .C2(new_n377), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G87), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n424), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n422), .A2(new_n428), .A3(new_n269), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G190), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n428), .A2(new_n269), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n421), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G200), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n413), .A2(new_n420), .A3(new_n430), .A4(new_n433), .ZN(new_n434));
  XNOR2_X1  g0234(.A(KEYINPUT83), .B(KEYINPUT17), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g0236(.A1(KEYINPUT83), .A2(KEYINPUT17), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n413), .A2(new_n420), .ZN(new_n439));
  AOI21_X1  g0239(.A(G169), .B1(new_n431), .B2(new_n421), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n440), .B1(new_n371), .B2(new_n429), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n439), .A2(KEYINPUT18), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(KEYINPUT18), .B1(new_n439), .B2(new_n441), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n436), .A2(new_n438), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n382), .A2(G200), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n445), .A2(KEYINPUT74), .B1(new_n446), .B2(G190), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n446), .A2(KEYINPUT74), .A3(G190), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n447), .A2(new_n448), .A3(new_n396), .ZN(new_n449));
  OR2_X1    g0249(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n398), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT6), .ZN(new_n452));
  INV_X1    g0252(.A(G107), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n228), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(G97), .A2(G107), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n453), .A2(KEYINPUT6), .A3(G97), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n281), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(G107), .B1(new_n400), .B2(new_n402), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n350), .A2(new_n388), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n459), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n308), .A2(new_n336), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT84), .ZN(new_n465));
  XNOR2_X1  g0265(.A(KEYINPUT70), .B(G1), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n465), .B1(new_n466), .B2(new_n294), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n274), .A2(KEYINPUT84), .A3(G33), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n463), .A2(new_n284), .B1(new_n469), .B2(G97), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n300), .A2(new_n228), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT5), .B(G41), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n274), .A2(new_n472), .A3(G45), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n264), .A2(new_n268), .ZN(new_n475));
  INV_X1    g0275(.A(G45), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n476), .B1(new_n271), .B2(new_n273), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n264), .B1(new_n477), .B2(new_n472), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n474), .A2(new_n475), .B1(new_n478), .B2(G257), .ZN(new_n479));
  OAI211_X1 g0279(.A(G244), .B(new_n257), .C1(new_n376), .C2(new_n377), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT85), .ZN(new_n481));
  OR2_X1    g0281(.A1(new_n481), .A2(KEYINPUT4), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n256), .A2(G250), .A3(G1698), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n257), .A2(G244), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n256), .A2(new_n482), .A3(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n484), .A2(new_n485), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n264), .ZN(new_n490));
  INV_X1    g0290(.A(G190), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n479), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(G200), .B1(new_n479), .B2(new_n490), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n470), .B(new_n471), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n464), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n467), .A2(new_n468), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(G97), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n401), .B1(new_n256), .B2(G20), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n399), .A2(KEYINPUT7), .A3(new_n281), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n453), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n500), .A2(new_n458), .A3(new_n461), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n471), .B(new_n497), .C1(new_n501), .C2(new_n336), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n479), .A2(new_n490), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n383), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n479), .A2(new_n490), .A3(new_n371), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n494), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT86), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT21), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n283), .A2(new_n213), .B1(G20), .B2(new_n219), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n485), .B(new_n281), .C1(G33), .C2(new_n228), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n511), .A2(KEYINPUT20), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT20), .B1(new_n511), .B2(new_n512), .ZN(new_n514));
  OAI22_X1  g0314(.A1(new_n513), .A2(new_n514), .B1(G116), .B2(new_n308), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n219), .B1(new_n467), .B2(new_n468), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n515), .B1(new_n338), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n473), .A2(G270), .A3(new_n424), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n477), .A2(new_n424), .A3(G274), .A4(new_n472), .ZN(new_n519));
  OR2_X1    g0319(.A1(KEYINPUT3), .A2(G33), .ZN(new_n520));
  INV_X1    g0320(.A(G303), .ZN(new_n521));
  NAND2_X1  g0321(.A1(KEYINPUT3), .A2(G33), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G264), .A2(G1698), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n229), .B2(G1698), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n523), .B(new_n264), .C1(new_n399), .C2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n518), .A2(new_n519), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G169), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n510), .B1(new_n517), .B2(new_n528), .ZN(new_n529));
  AOI211_X1 g0329(.A(KEYINPUT76), .B(new_n284), .C1(new_n282), .C2(G13), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n335), .B1(new_n308), .B2(new_n336), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n516), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n514), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n511), .A2(KEYINPUT20), .A3(new_n512), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n533), .A2(new_n534), .B1(new_n219), .B2(new_n300), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n519), .A2(new_n526), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n383), .B1(new_n537), .B2(new_n518), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(KEYINPUT21), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(G179), .A3(new_n518), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n517), .A2(KEYINPUT89), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT89), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n527), .A2(new_n371), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(new_n536), .B2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n529), .B(new_n539), .C1(new_n541), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n229), .A2(G1698), .ZN(new_n546));
  OAI221_X1 g0346(.A(new_n546), .B1(G250), .B2(G1698), .C1(new_n376), .C2(new_n377), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G294), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n264), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n478), .A2(G264), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n550), .A2(new_n551), .A3(new_n519), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n383), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(G179), .B2(new_n552), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT24), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT23), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n281), .B2(G107), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n453), .A2(KEYINPUT23), .A3(G20), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n295), .A2(G116), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n281), .B(G87), .C1(new_n376), .C2(new_n377), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT22), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT22), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n256), .A2(new_n564), .A3(new_n281), .A4(G87), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n561), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n555), .B1(new_n566), .B2(KEYINPUT90), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n563), .A2(new_n565), .ZN(new_n568));
  INV_X1    g0368(.A(new_n561), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT90), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n570), .A2(new_n571), .A3(new_n555), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n284), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT25), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n308), .B2(G107), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n300), .A2(KEYINPUT25), .A3(new_n453), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n469), .A2(G107), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n554), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n527), .A2(new_n491), .ZN(new_n581));
  AOI211_X1 g0381(.A(new_n581), .B(new_n536), .C1(G200), .C2(new_n527), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n545), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n552), .A2(new_n255), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(G190), .B2(new_n552), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n575), .A2(new_n585), .A3(new_n579), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT88), .ZN(new_n587));
  OAI211_X1 g0387(.A(G238), .B(new_n257), .C1(new_n376), .C2(new_n377), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT87), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT87), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n256), .A2(new_n590), .A3(G238), .A4(new_n257), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G116), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n256), .A2(G244), .A3(G1698), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n589), .A2(new_n591), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n264), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n264), .B1(new_n477), .B2(new_n268), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n232), .B1(new_n466), .B2(new_n476), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n587), .B1(new_n599), .B2(G179), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n495), .A2(new_n391), .A3(new_n496), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n300), .A2(new_n392), .ZN(new_n602));
  NOR3_X1   g0402(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n319), .A2(new_n321), .A3(KEYINPUT19), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n603), .B1(new_n604), .B2(new_n281), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n256), .A2(new_n281), .A3(G68), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT19), .B1(new_n295), .B2(G97), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n605), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n601), .B(new_n602), .C1(new_n609), .C2(new_n336), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n599), .A2(new_n383), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n594), .A2(new_n264), .B1(new_n597), .B2(new_n596), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(KEYINPUT88), .A3(new_n371), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n600), .A2(new_n610), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n495), .A2(G87), .A3(new_n496), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n615), .B(new_n602), .C1(new_n609), .C2(new_n336), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n599), .A2(G200), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n595), .A2(G190), .A3(new_n598), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n586), .A2(new_n614), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n508), .B1(new_n494), .B2(new_n506), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n451), .A2(new_n509), .A3(new_n583), .A4(new_n623), .ZN(G372));
  NAND2_X1  g0424(.A1(new_n366), .A2(new_n367), .ZN(new_n625));
  INV_X1    g0425(.A(new_n356), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n625), .B1(new_n626), .B2(new_n397), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n434), .A2(new_n435), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(new_n437), .B2(new_n434), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n439), .A2(new_n441), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT18), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n439), .A2(KEYINPUT18), .A3(new_n441), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n316), .B1(new_n630), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n374), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n451), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n612), .A2(new_n371), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n611), .A2(new_n610), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n580), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n541), .A2(new_n544), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n529), .A2(new_n539), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT92), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n517), .A2(new_n510), .A3(new_n528), .ZN(new_n648));
  AOI21_X1  g0448(.A(KEYINPUT21), .B1(new_n536), .B2(new_n538), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT89), .B1(new_n517), .B2(new_n540), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n536), .A2(new_n542), .A3(new_n543), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT92), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n643), .B1(new_n647), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n642), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n616), .A2(KEYINPUT91), .ZN(new_n657));
  INV_X1    g0457(.A(new_n608), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n604), .A2(new_n281), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n606), .B(new_n658), .C1(new_n659), .C2(new_n603), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n284), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT91), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n661), .A2(new_n662), .A3(new_n602), .A4(new_n615), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n619), .B1(new_n255), .B2(new_n612), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  AND4_X1   g0467(.A1(new_n507), .A2(new_n586), .A3(new_n656), .A4(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n642), .B1(new_n655), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n665), .B1(new_n657), .B2(new_n663), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n670), .A2(new_n506), .A3(new_n642), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT93), .B1(new_n671), .B2(KEYINPUT26), .ZN(new_n672));
  INV_X1    g0472(.A(new_n506), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n673), .A2(new_n614), .A3(KEYINPUT26), .A4(new_n620), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n667), .A2(new_n656), .A3(new_n673), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT93), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n672), .A2(new_n674), .A3(new_n678), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n669), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n639), .B1(new_n640), .B2(new_n680), .ZN(G369));
  NOR2_X1   g0481(.A1(new_n545), .A2(new_n582), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n647), .A2(new_n654), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n281), .A2(G13), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n466), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT27), .ZN(new_n686));
  OR3_X1    g0486(.A1(new_n685), .A2(KEYINPUT94), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G213), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n685), .B2(new_n686), .ZN(new_n689));
  OAI21_X1  g0489(.A(KEYINPUT94), .B1(new_n685), .B2(new_n686), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n687), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g0492(.A(KEYINPUT95), .B(G343), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(new_n517), .ZN(new_n695));
  MUX2_X1   g0495(.A(new_n682), .B(new_n683), .S(new_n695), .Z(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n580), .A2(new_n694), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n575), .A2(new_n579), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n586), .B1(new_n701), .B2(new_n694), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n700), .B1(new_n702), .B2(new_n643), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n545), .ZN(new_n705));
  INV_X1    g0505(.A(new_n694), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(new_n700), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n704), .A2(new_n709), .ZN(G399));
  INV_X1    g0510(.A(new_n212), .ZN(new_n711));
  INV_X1    g0511(.A(new_n204), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G41), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n603), .A2(new_n219), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(G1), .ZN(new_n716));
  OAI22_X1  g0516(.A1(new_n711), .A2(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT28), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n705), .A2(new_n643), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n668), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n673), .A2(new_n614), .A3(new_n677), .A4(new_n620), .ZN(new_n722));
  OAI211_X1 g0522(.A(new_n656), .B(new_n722), .C1(new_n671), .C2(new_n677), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n694), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n706), .B1(new_n669), .B2(new_n679), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT96), .ZN(new_n726));
  OAI211_X1 g0526(.A(KEYINPUT29), .B(new_n724), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(G330), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n623), .A2(new_n583), .A3(new_n509), .A4(new_n694), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n543), .A2(new_n612), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n264), .A2(new_n549), .B1(new_n478), .B2(G264), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n479), .A2(new_n732), .A3(new_n490), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n730), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  AND3_X1   g0534(.A1(new_n479), .A2(new_n732), .A3(new_n490), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(KEYINPUT30), .A3(new_n543), .A4(new_n612), .ZN(new_n736));
  AOI21_X1  g0536(.A(G179), .B1(new_n479), .B2(new_n490), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n737), .A2(new_n552), .A3(new_n527), .A4(new_n599), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n734), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n706), .ZN(new_n740));
  AOI21_X1  g0540(.A(KEYINPUT31), .B1(new_n739), .B2(new_n706), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n728), .B1(new_n729), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT29), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(new_n725), .B2(KEYINPUT96), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n727), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n718), .B1(new_n748), .B2(G1), .ZN(new_n749));
  XOR2_X1   g0549(.A(new_n749), .B(KEYINPUT97), .Z(G364));
  OR2_X1    g0550(.A1(new_n696), .A2(G330), .ZN(new_n751));
  XOR2_X1   g0551(.A(new_n684), .B(KEYINPUT98), .Z(new_n752));
  AOI21_X1  g0552(.A(new_n716), .B1(G45), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n751), .A2(new_n697), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT99), .ZN(new_n756));
  OAI21_X1  g0556(.A(G20), .B1(KEYINPUT100), .B2(G169), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(KEYINPUT100), .A2(G169), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n213), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n281), .A2(G190), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n762), .A2(KEYINPUT101), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G179), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n762), .A2(KEYINPUT101), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G159), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n255), .A2(G179), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n763), .A2(new_n765), .A3(new_n770), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n769), .A2(KEYINPUT32), .B1(new_n453), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n281), .B1(new_n764), .B2(G190), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT102), .Z(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n772), .B1(G97), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n281), .A2(new_n491), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n770), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n231), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n371), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n491), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n256), .B1(new_n781), .B2(new_n226), .C1(new_n217), .C2(new_n784), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n779), .B(new_n785), .C1(new_n769), .C2(KEYINPUT32), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n776), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n782), .A2(G190), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n762), .A2(new_n780), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n787), .B1(new_n345), .B2(new_n789), .C1(new_n388), .C2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n778), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G303), .ZN(new_n793));
  INV_X1    g0593(.A(G329), .ZN(new_n794));
  INV_X1    g0594(.A(G311), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n766), .A2(new_n794), .B1(new_n795), .B2(new_n790), .ZN(new_n796));
  INV_X1    g0596(.A(new_n773), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n796), .B1(G294), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G317), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n789), .B1(KEYINPUT33), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(KEYINPUT33), .B2(new_n799), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n256), .B1(new_n783), .B2(G326), .ZN(new_n802));
  AND4_X1   g0602(.A1(new_n793), .A2(new_n798), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G283), .ZN(new_n804));
  INV_X1    g0604(.A(G322), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n803), .B1(new_n804), .B2(new_n771), .C1(new_n805), .C2(new_n781), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n761), .B1(new_n791), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n256), .A2(G355), .A3(new_n204), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n712), .A2(new_n256), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n711), .B2(G45), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n250), .A2(new_n476), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n808), .B1(G116), .B2(new_n204), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(G13), .A2(G33), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(G20), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n760), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n815), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n817), .B(new_n753), .C1(new_n696), .C2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n756), .B1(new_n807), .B2(new_n819), .ZN(G396));
  INV_X1    g0620(.A(KEYINPUT105), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n397), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n386), .A2(new_n396), .A3(KEYINPUT105), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n449), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n725), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n397), .A2(new_n694), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n706), .A2(new_n396), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n826), .B1(new_n824), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n825), .B1(new_n725), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(new_n743), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n754), .ZN(new_n832));
  INV_X1    g0632(.A(G294), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n774), .A2(new_n228), .B1(new_n833), .B2(new_n781), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT103), .ZN(new_n835));
  INV_X1    g0635(.A(new_n771), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n835), .B1(G87), .B2(new_n836), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n837), .B1(new_n219), .B2(new_n790), .C1(new_n795), .C2(new_n766), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n789), .A2(new_n804), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n784), .A2(new_n521), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n399), .B1(new_n778), .B2(new_n453), .ZN(new_n841));
  NOR4_X1   g0641(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n771), .A2(new_n345), .ZN(new_n843));
  INV_X1    g0643(.A(new_n766), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n399), .B1(new_n844), .B2(G132), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n781), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n847), .A2(G143), .B1(G150), .B2(new_n788), .ZN(new_n848));
  INV_X1    g0648(.A(G137), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n848), .B1(new_n849), .B2(new_n784), .C1(new_n767), .C2(new_n790), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT34), .ZN(new_n851));
  AOI22_X1  g0651(.A1(KEYINPUT104), .A2(new_n846), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT104), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n845), .A2(new_n853), .B1(G58), .B2(new_n797), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n852), .B(new_n854), .C1(new_n851), .C2(new_n850), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n843), .B(new_n855), .C1(G50), .C2(new_n792), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n760), .B1(new_n842), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n760), .A2(new_n813), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n388), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n828), .A2(new_n813), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n857), .A2(new_n753), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n832), .A2(new_n861), .ZN(G384));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n439), .A2(new_n692), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n863), .B1(new_n864), .B2(KEYINPUT107), .ZN(new_n865));
  AND4_X1   g0665(.A1(new_n413), .A2(new_n420), .A3(new_n430), .A4(new_n433), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n691), .B1(new_n413), .B2(new_n420), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n865), .A2(new_n868), .A3(new_n631), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n631), .A2(new_n864), .A3(new_n434), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT107), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT37), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n864), .B1(new_n635), .B2(new_n629), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n874), .A2(new_n876), .A3(KEYINPUT38), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n869), .A2(new_n873), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n878), .B1(new_n879), .B2(new_n875), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  AND4_X1   g0681(.A1(KEYINPUT37), .A2(new_n631), .A3(new_n864), .A4(new_n434), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n444), .B2(new_n867), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n870), .A2(new_n863), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT38), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NOR3_X1   g0685(.A1(new_n879), .A2(new_n875), .A3(new_n878), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT39), .ZN(new_n888));
  MUX2_X1   g0688(.A(new_n881), .B(new_n887), .S(new_n888), .Z(new_n889));
  NOR2_X1   g0689(.A1(new_n625), .A2(new_n706), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n822), .A2(new_n694), .A3(new_n823), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n825), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n358), .A2(new_n694), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n625), .A2(new_n356), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n368), .B2(new_n895), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n893), .A2(new_n897), .A3(new_n881), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n636), .A2(new_n691), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n891), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT109), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n727), .A2(new_n746), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n638), .B1(new_n902), .B2(new_n451), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n901), .B(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n828), .B1(new_n729), .B2(new_n742), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT108), .B1(new_n905), .B2(new_n897), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT40), .B1(new_n887), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT40), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n877), .A2(new_n908), .A3(new_n880), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n729), .A2(new_n742), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n897), .A2(new_n910), .A3(new_n829), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n908), .A2(KEYINPUT108), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n909), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n907), .A2(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n914), .A2(new_n910), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(G330), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n640), .A2(new_n744), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n915), .A2(new_n451), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n904), .B(new_n919), .Z(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n274), .B2(new_n752), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n212), .A2(G77), .A3(new_n404), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(G50), .B2(new_n345), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(new_n299), .A3(new_n466), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n456), .A2(new_n457), .ZN(new_n925));
  OAI211_X1 g0725(.A(G20), .B(new_n214), .C1(new_n925), .C2(KEYINPUT35), .ZN(new_n926));
  AOI211_X1 g0726(.A(new_n219), .B(new_n926), .C1(KEYINPUT35), .C2(new_n925), .ZN(new_n927));
  XNOR2_X1  g0727(.A(KEYINPUT106), .B(KEYINPUT36), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n927), .B(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n921), .A2(new_n924), .A3(new_n929), .ZN(G367));
  NAND3_X1  g0730(.A1(new_n792), .A2(KEYINPUT46), .A3(G116), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT46), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n778), .B2(new_n219), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n931), .B(new_n933), .C1(new_n833), .C2(new_n789), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n934), .A2(KEYINPUT111), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n766), .A2(new_n799), .B1(new_n521), .B2(new_n781), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n399), .B1(new_n773), .B2(new_n453), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n783), .A2(G311), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n771), .A2(new_n228), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n790), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n934), .A2(KEYINPUT111), .B1(G283), .B2(new_n942), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n938), .A2(new_n939), .A3(new_n941), .A4(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n774), .A2(new_n345), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n778), .A2(new_n226), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n783), .A2(G143), .ZN(new_n947));
  NOR4_X1   g0747(.A1(new_n945), .A2(new_n399), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n788), .A2(G159), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n771), .A2(new_n388), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(G150), .B2(new_n847), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n942), .A2(G50), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n948), .A2(new_n949), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n766), .A2(new_n849), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n944), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT47), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n760), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n706), .A2(new_n657), .A3(new_n663), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n656), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n667), .A2(new_n656), .A3(new_n958), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n959), .A2(new_n815), .A3(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n809), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n816), .B1(new_n204), .B2(new_n392), .C1(new_n245), .C2(new_n962), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n957), .A2(new_n961), .A3(new_n753), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n752), .A2(G45), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(G1), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n706), .A2(new_n502), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n507), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n506), .B2(new_n694), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n709), .A2(new_n969), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n970), .A2(KEYINPUT110), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n970), .A2(KEYINPUT110), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT45), .ZN(new_n973));
  OR3_X1    g0773(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n709), .A2(new_n969), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT44), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n973), .B1(new_n971), .B2(new_n972), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n974), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n704), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n978), .B(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n703), .B(new_n707), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n697), .B(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n748), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n713), .B(KEYINPUT41), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n966), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n708), .A2(new_n507), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT42), .Z(new_n987));
  OAI21_X1  g0787(.A(new_n506), .B1(new_n968), .B2(new_n643), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n694), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n959), .A2(new_n960), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n987), .A2(new_n989), .B1(KEYINPUT43), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n991), .B(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n979), .A2(new_n969), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n993), .B(new_n994), .Z(new_n995));
  OAI21_X1  g0795(.A(new_n964), .B1(new_n985), .B2(new_n995), .ZN(G387));
  OR2_X1    g0796(.A1(new_n747), .A2(new_n982), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n714), .B1(new_n747), .B2(new_n982), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n847), .A2(G317), .B1(G311), .B2(new_n788), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n521), .B2(new_n790), .C1(new_n805), .C2(new_n784), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT48), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n804), .B2(new_n773), .C1(new_n833), .C2(new_n778), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT49), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n256), .B1(new_n844), .B2(G326), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1004), .B(new_n1005), .C1(new_n219), .C2(new_n771), .ZN(new_n1006));
  INV_X1    g0806(.A(G150), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n766), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n774), .A2(new_n392), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1008), .B(new_n1009), .C1(G159), .C2(new_n783), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n293), .A2(new_n789), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n778), .A2(new_n388), .B1(new_n790), .B2(new_n345), .ZN(new_n1012));
  NOR3_X1   g0812(.A1(new_n940), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n847), .A2(G50), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1010), .A2(new_n256), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n761), .B1(new_n1006), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n809), .B1(new_n242), .B2(new_n476), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n715), .A2(new_n204), .A3(new_n256), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n289), .A2(G50), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT50), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1021), .B(new_n476), .C1(new_n345), .C2(new_n388), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1019), .B1(new_n715), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n712), .A2(new_n453), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n760), .B(new_n815), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n753), .B1(new_n703), .B2(new_n818), .ZN(new_n1026));
  OR3_X1    g0826(.A1(new_n1016), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n966), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n999), .B(new_n1027), .C1(new_n1028), .C2(new_n982), .ZN(G393));
  OAI21_X1  g0829(.A(new_n816), .B1(new_n228), .B2(new_n204), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n253), .B2(new_n809), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n847), .A2(G311), .B1(G317), .B2(new_n783), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT52), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n790), .A2(new_n833), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n771), .A2(new_n453), .B1(new_n804), .B2(new_n778), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n399), .B1(new_n789), .B2(new_n521), .ZN(new_n1036));
  NOR4_X1   g0836(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n219), .B2(new_n773), .C1(new_n805), .C2(new_n766), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT112), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n774), .A2(new_n388), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n778), .A2(new_n345), .B1(new_n790), .B2(new_n289), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n399), .B(new_n1041), .C1(new_n836), .C2(G87), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n784), .A2(new_n1007), .B1(new_n781), .B2(new_n767), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT51), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n844), .A2(G143), .B1(new_n788), .B2(G50), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1042), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1039), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n754), .B(new_n1031), .C1(new_n1047), .C2(new_n760), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n818), .B2(new_n969), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n980), .B2(new_n1028), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n980), .A2(new_n997), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n714), .B1(new_n980), .B2(new_n997), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1050), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(G390));
  XNOR2_X1  g0854(.A(new_n890), .B(KEYINPUT113), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n892), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n723), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n706), .B1(new_n1057), .B2(new_n720), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1056), .B1(new_n1058), .B2(new_n824), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n897), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1055), .B1(new_n886), .B2(new_n885), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n890), .B1(new_n893), .B2(new_n897), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1061), .B1(new_n1062), .B2(new_n889), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n911), .A2(G330), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1061), .B(new_n1064), .C1(new_n1062), .C2(new_n889), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT114), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n903), .B2(new_n918), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n640), .B1(new_n727), .B2(new_n746), .ZN(new_n1071));
  NOR4_X1   g0871(.A1(new_n1071), .A2(KEYINPUT114), .A3(new_n638), .A4(new_n917), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n905), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1060), .B1(new_n1073), .B2(new_n728), .ZN(new_n1074));
  AND3_X1   g0874(.A1(new_n1064), .A2(new_n1074), .A3(new_n1059), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1064), .A2(new_n1074), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1075), .B1(new_n893), .B2(new_n1076), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n1070), .A2(new_n1072), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT115), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1068), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n902), .A2(new_n451), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1081), .A2(new_n639), .A3(new_n918), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(KEYINPUT114), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1077), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n903), .A2(new_n1069), .A3(new_n918), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1086), .A2(KEYINPUT115), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1080), .A2(new_n713), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n858), .A2(new_n293), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n889), .A2(new_n814), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n843), .B(new_n1040), .C1(G97), .C2(new_n942), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n399), .B1(new_n781), .B2(new_n219), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n779), .B(new_n1093), .C1(G283), .C2(new_n783), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1095), .B1(new_n453), .B2(new_n789), .C1(new_n833), .C2(new_n766), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n847), .A2(G132), .ZN(new_n1097));
  INV_X1    g0897(.A(G128), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n256), .B1(new_n789), .B2(new_n849), .C1(new_n1098), .C2(new_n784), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1097), .B(new_n1099), .C1(G125), .C2(new_n844), .ZN(new_n1100));
  XOR2_X1   g0900(.A(KEYINPUT54), .B(G143), .Z(new_n1101));
  NAND2_X1  g0901(.A1(new_n942), .A2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n775), .A2(G159), .B1(G50), .B2(new_n836), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n778), .A2(new_n1007), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT53), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1100), .A2(new_n1102), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n761), .B1(new_n1096), .B2(new_n1106), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n1091), .A2(new_n754), .A3(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1068), .A2(new_n966), .B1(new_n1090), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1089), .A2(new_n1109), .ZN(G378));
  INV_X1    g0910(.A(new_n900), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n316), .A2(new_n374), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1112), .B(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n302), .A2(new_n691), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT119), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1114), .B(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n728), .B1(new_n907), .B2(new_n913), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1117), .B1(new_n1118), .B2(KEYINPUT120), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT120), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1120), .B(new_n728), .C1(new_n907), .C2(new_n913), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n916), .A2(new_n1117), .A3(new_n1120), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1111), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n916), .A2(new_n1120), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1118), .A2(KEYINPUT120), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1125), .A2(new_n1126), .A3(new_n1117), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1127), .A2(new_n1128), .A3(new_n900), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1124), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n966), .ZN(new_n1131));
  OR2_X1    g0931(.A1(new_n1117), .A2(new_n814), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n858), .A2(new_n217), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n945), .B1(G97), .B2(new_n788), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n423), .B(new_n399), .C1(new_n778), .C2(new_n388), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT116), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n766), .A2(new_n804), .B1(new_n219), .B2(new_n784), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(G58), .B2(new_n836), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1134), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(new_n453), .B2(new_n781), .C1(new_n392), .C2(new_n790), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT58), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n217), .B1(new_n376), .B2(G41), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(KEYINPUT117), .B(G124), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n766), .A2(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n775), .A2(G150), .B1(G137), .B2(new_n942), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n847), .A2(G128), .B1(G132), .B2(new_n788), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1101), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1145), .B(new_n1146), .C1(new_n778), .C2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(G125), .B2(new_n783), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT59), .ZN(new_n1150));
  AOI211_X1 g0950(.A(G41), .B(new_n1144), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1151), .B(new_n294), .C1(new_n767), .C2(new_n771), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1141), .B(new_n1142), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT118), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n760), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1132), .A2(new_n753), .A3(new_n1133), .A4(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1131), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1066), .A2(new_n1084), .A3(new_n1067), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n1122), .A2(new_n1111), .A3(new_n1123), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n900), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT57), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n714), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT121), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1124), .A2(new_n1129), .A3(new_n1167), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1127), .A2(new_n1128), .A3(KEYINPUT121), .A4(new_n900), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1168), .A2(KEYINPUT57), .A3(new_n1169), .A4(new_n1161), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1158), .B1(new_n1166), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(G375));
  NAND2_X1  g0972(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n1077), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1174), .A2(new_n984), .A3(new_n1086), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n771), .A2(new_n226), .B1(new_n789), .B2(new_n1147), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n399), .B(new_n1176), .C1(G132), .C2(new_n783), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n775), .A2(G50), .B1(G150), .B2(new_n942), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(new_n849), .C2(new_n781), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n766), .A2(new_n1098), .B1(new_n767), .B2(new_n778), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT122), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n766), .A2(new_n521), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n256), .B(new_n950), .C1(G294), .C2(new_n783), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1009), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n788), .A2(G116), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n778), .A2(new_n228), .B1(new_n790), .B2(new_n453), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G283), .B2(new_n847), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .A4(new_n1187), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n1179), .A2(new_n1181), .B1(new_n1182), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n760), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n753), .B(new_n1190), .C1(new_n897), .C2(new_n814), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n345), .B2(new_n858), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n1084), .B2(new_n966), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1175), .A2(new_n1193), .ZN(G381));
  NOR2_X1   g0994(.A1(G381), .A2(G384), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1053), .B(new_n964), .C1(new_n985), .C2(new_n995), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(G375), .A2(G378), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(G393), .A2(G396), .ZN(new_n1199));
  AND4_X1   g0999(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n1200), .A2(KEYINPUT123), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1200), .A2(KEYINPUT123), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1201), .A2(new_n1202), .ZN(G407));
  NOR2_X1   g1003(.A1(new_n693), .A2(new_n688), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT124), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1198), .A2(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(G213), .B(new_n1207), .C1(new_n1201), .C2(new_n1202), .ZN(G409));
  XNOR2_X1  g1008(.A(G393), .B(G396), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1209), .A2(KEYINPUT126), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(G387), .A2(G390), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1210), .B1(new_n1211), .B2(new_n1196), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1209), .B(KEYINPUT126), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1211), .A2(new_n1196), .A3(new_n1214), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1166), .A2(new_n1170), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1158), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1217), .A2(G378), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1157), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1124), .A2(new_n1129), .B1(new_n1160), .B2(new_n1159), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1220), .B1(new_n1221), .B2(new_n984), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1168), .A2(new_n966), .A3(new_n1169), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(G378), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1204), .B1(new_n1219), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT60), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1174), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1173), .A2(KEYINPUT60), .A3(new_n1077), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1229), .A2(new_n713), .A3(new_n1086), .A4(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1231), .A2(G384), .A3(new_n1193), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(G384), .B1(new_n1231), .B2(new_n1193), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT62), .B1(new_n1227), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(G378), .B1(new_n1223), .B2(new_n1222), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G378), .B2(new_n1171), .ZN(new_n1238));
  OAI21_X1  g1038(.A(KEYINPUT127), .B1(new_n1238), .B2(new_n1206), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1219), .A2(new_n1226), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT127), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1240), .A2(new_n1241), .A3(new_n1205), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1239), .A2(new_n1242), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1235), .A2(KEYINPUT62), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1236), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1231), .A2(new_n1193), .ZN(new_n1246));
  INV_X1    g1046(.A(G384), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1205), .B1(new_n1248), .B2(new_n1232), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1204), .A2(G2897), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(G2897), .A2(new_n1249), .B1(new_n1235), .B2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1239), .A2(new_n1242), .A3(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT61), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1216), .B1(new_n1245), .B2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1243), .A2(KEYINPUT63), .A3(new_n1235), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT61), .B1(new_n1213), .B2(new_n1215), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1227), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(KEYINPUT125), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT125), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1227), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n1251), .A3(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT63), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1235), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1263), .B1(new_n1258), .B2(new_n1264), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1256), .A2(new_n1257), .A3(new_n1262), .A4(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1255), .A2(new_n1266), .ZN(G405));
  NAND2_X1  g1067(.A1(G375), .A2(new_n1225), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1219), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1269), .B(new_n1235), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1270), .B(new_n1216), .ZN(G402));
endmodule


