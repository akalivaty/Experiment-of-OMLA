//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n574, new_n575,
    new_n576, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1126, new_n1127, new_n1128;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT66), .B(KEYINPUT67), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  OR4_X1    g029(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT68), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(new_n467), .A3(G137), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n468), .A2(KEYINPUT70), .A3(new_n469), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G113), .ZN(new_n476));
  INV_X1    g051(.A(G2104), .ZN(new_n477));
  OR3_X1    g052(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT69), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT69), .B1(new_n476), .B2(new_n477), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n477), .A2(KEYINPUT3), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n478), .B(new_n479), .C1(new_n480), .C2(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(KEYINPUT68), .B(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n475), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G160));
  NAND2_X1  g064(.A1(new_n467), .A2(new_n486), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n467), .A2(new_n462), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G136), .ZN(new_n495));
  OAI221_X1 g070(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n466), .C2(G112), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n492), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G162));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n466), .A2(new_n467), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n481), .A2(new_n483), .A3(G126), .ZN(new_n503));
  NAND2_X1  g078(.A1(G114), .A2(G2104), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G2105), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n462), .A2(G102), .A3(G2104), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n499), .A2(new_n501), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n466), .A2(new_n467), .A3(new_n508), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n502), .A2(new_n506), .A3(new_n507), .A4(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n512));
  AND3_X1   g087(.A1(new_n512), .A2(KEYINPUT6), .A3(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(KEYINPUT6), .B1(new_n512), .B2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(G50), .A2(new_n517), .B1(new_n522), .B2(G88), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n518), .A2(new_n520), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n524), .A2(KEYINPUT72), .A3(G62), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n527));
  INV_X1    g102(.A(G62), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n521), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n525), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n523), .A2(new_n531), .ZN(G303));
  INV_X1    g107(.A(G303), .ZN(G166));
  NAND2_X1  g108(.A1(new_n517), .A2(G51), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n513), .A2(new_n514), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n537), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n538));
  OAI211_X1 g113(.A(new_n534), .B(new_n536), .C1(new_n538), .C2(new_n521), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(G168));
  AOI22_X1  g115(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G651), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(G52), .B2(new_n517), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n522), .A2(G90), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  XNOR2_X1  g122(.A(KEYINPUT73), .B(G43), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n517), .A2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n537), .A2(new_n524), .ZN(new_n552));
  OAI221_X1 g127(.A(new_n549), .B1(new_n542), .B2(new_n550), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n537), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n517), .A2(KEYINPUT9), .A3(G53), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n521), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n522), .A2(G91), .B1(G651), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G299));
  NAND2_X1  g148(.A1(G168), .A2(KEYINPUT74), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n539), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(G286));
  NAND2_X1  g152(.A1(new_n517), .A2(G49), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n522), .A2(G87), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  AND2_X1   g156(.A1(new_n537), .A2(G48), .ZN(new_n582));
  AND2_X1   g157(.A1(G73), .A2(G651), .ZN(new_n583));
  OAI21_X1  g158(.A(G543), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n515), .A2(new_n585), .ZN(new_n586));
  AND2_X1   g161(.A1(G61), .A2(G651), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n524), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(G72), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G60), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n521), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n517), .A2(G47), .B1(G651), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n522), .A2(G85), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  INV_X1    g172(.A(G92), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n552), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n522), .A2(KEYINPUT10), .A3(G92), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n601), .A2(G66), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(G66), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n524), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G79), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n516), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n599), .A2(new_n600), .B1(G651), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n517), .A2(G54), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n596), .B1(new_n610), .B2(G868), .ZN(G284));
  OAI21_X1  g186(.A(new_n596), .B1(new_n610), .B2(G868), .ZN(G321));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(G299), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(G286), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n613), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(new_n613), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n610), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n553), .A2(new_n613), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n609), .A2(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n613), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g198(.A1(G123), .A2(new_n491), .B1(new_n494), .B2(G135), .ZN(new_n624));
  OAI221_X1 g199(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n466), .C2(G111), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT78), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2096), .ZN(new_n628));
  XOR2_X1   g203(.A(KEYINPUT76), .B(KEYINPUT12), .Z(new_n629));
  NOR3_X1   g204(.A1(new_n482), .A2(new_n477), .A3(G2105), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT77), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n631), .B(new_n634), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n628), .B(new_n635), .C1(KEYINPUT77), .C2(new_n632), .ZN(G156));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2430), .ZN(new_n638));
  XOR2_X1   g213(.A(KEYINPUT15), .B(G2435), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(KEYINPUT14), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2443), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n647), .B(new_n648), .Z(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(G14), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(G401));
  XOR2_X1   g226(.A(G2067), .B(G2678), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT18), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n653), .A2(new_n654), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n656), .B(KEYINPUT17), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(new_n661), .A3(new_n655), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n656), .B(KEYINPUT80), .Z(new_n663));
  OAI211_X1 g238(.A(new_n658), .B(new_n662), .C1(new_n660), .C2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2096), .B(G2100), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT81), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n664), .B(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n669), .A2(new_n670), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT82), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n675), .B1(new_n678), .B2(KEYINPUT20), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n672), .A2(new_n674), .A3(new_n676), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n679), .B(new_n680), .C1(KEYINPUT20), .C2(new_n678), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1986), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1981), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1991), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n683), .B(new_n686), .ZN(G229));
  INV_X1    g262(.A(G29), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G26), .ZN(new_n689));
  AOI22_X1  g264(.A1(G128), .A2(new_n491), .B1(new_n494), .B2(G140), .ZN(new_n690));
  OAI221_X1 g265(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n466), .C2(G116), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT84), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n689), .B1(new_n694), .B2(new_n688), .ZN(new_n695));
  MUX2_X1   g270(.A(new_n689), .B(new_n695), .S(KEYINPUT28), .Z(new_n696));
  XOR2_X1   g271(.A(KEYINPUT85), .B(G2067), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G4), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(new_n610), .B2(new_n699), .ZN(new_n701));
  INV_X1    g276(.A(G1348), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT87), .ZN(new_n704));
  NOR2_X1   g279(.A1(KEYINPUT24), .A2(G34), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(KEYINPUT24), .A2(G34), .ZN(new_n707));
  AOI21_X1  g282(.A(G29), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AOI22_X1  g283(.A1(G160), .A2(G29), .B1(new_n704), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(new_n704), .B2(new_n708), .ZN(new_n710));
  INV_X1    g285(.A(G2084), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n699), .A2(G19), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n554), .B2(new_n699), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G1341), .ZN(new_n715));
  AND4_X1   g290(.A1(new_n698), .A2(new_n703), .A3(new_n712), .A4(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n714), .A2(G1341), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n688), .A2(G35), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G162), .B2(new_n688), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT29), .Z(new_n721));
  INV_X1    g296(.A(G2090), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n699), .A2(G21), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G168), .B2(new_n699), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n721), .A2(new_n722), .B1(G1966), .B2(new_n725), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n725), .A2(G1966), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n710), .A2(new_n711), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n723), .A2(new_n726), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT31), .B(G11), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n688), .A2(G27), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G164), .B2(new_n688), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT90), .Z(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G2078), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n699), .A2(G5), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G171), .B2(new_n699), .ZN(new_n738));
  INV_X1    g313(.A(G1961), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT89), .B(G28), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT30), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(new_n688), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n626), .B2(new_n688), .ZN(new_n744));
  OR2_X1    g319(.A1(G29), .A2(G32), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT88), .B(KEYINPUT26), .Z(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n491), .A2(G129), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n494), .A2(G141), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n748), .A2(new_n749), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n745), .B1(new_n752), .B2(new_n688), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT27), .B(G1996), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n744), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n740), .B(new_n755), .C1(new_n753), .C2(new_n754), .ZN(new_n756));
  NOR4_X1   g331(.A1(new_n729), .A2(new_n730), .A3(new_n736), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n699), .A2(G20), .ZN(new_n758));
  OAI211_X1 g333(.A(KEYINPUT23), .B(new_n758), .C1(new_n572), .C2(new_n699), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(KEYINPUT23), .B2(new_n758), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT91), .B(G1956), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n735), .B2(new_n734), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n716), .A2(new_n718), .A3(new_n757), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n699), .A2(G23), .ZN(new_n765));
  INV_X1    g340(.A(G288), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n765), .B1(new_n766), .B2(new_n699), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT33), .ZN(new_n768));
  INV_X1    g343(.A(G1976), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n699), .A2(G6), .ZN(new_n771));
  INV_X1    g346(.A(G305), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(new_n699), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT32), .B(G1981), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n699), .A2(G22), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G166), .B2(new_n699), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(G1971), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n777), .A2(G1971), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n775), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n770), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT34), .ZN(new_n782));
  AOI22_X1  g357(.A1(G119), .A2(new_n491), .B1(new_n494), .B2(G131), .ZN(new_n783));
  OAI221_X1 g358(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n466), .C2(G107), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  MUX2_X1   g360(.A(G25), .B(new_n785), .S(G29), .Z(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT35), .B(G1991), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT83), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n786), .B(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G16), .A2(G24), .ZN(new_n790));
  INV_X1    g365(.A(G290), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(G16), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(G1986), .Z(new_n793));
  NAND3_X1  g368(.A1(new_n782), .A2(new_n789), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(KEYINPUT36), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT36), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n782), .A2(new_n796), .A3(new_n789), .A4(new_n793), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n764), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT25), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n494), .A2(G139), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n800), .B(new_n801), .C1(new_n466), .C2(new_n802), .ZN(new_n803));
  MUX2_X1   g378(.A(G33), .B(new_n803), .S(G29), .Z(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT86), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G2072), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n798), .A2(new_n807), .ZN(G311));
  NAND2_X1  g383(.A1(new_n798), .A2(new_n807), .ZN(G150));
  NAND2_X1  g384(.A1(new_n522), .A2(G93), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n517), .A2(G55), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n810), .B(new_n811), .C1(new_n542), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G860), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT37), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n553), .B(new_n813), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT92), .B(KEYINPUT38), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n609), .A2(new_n618), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT39), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n818), .B(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n815), .B1(new_n821), .B2(G860), .ZN(G145));
  NAND2_X1  g397(.A1(new_n491), .A2(G130), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT94), .ZN(new_n824));
  OAI221_X1 g399(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n466), .C2(G118), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n494), .A2(G142), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(new_n785), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(new_n631), .Z(new_n829));
  NOR2_X1   g404(.A1(new_n803), .A2(KEYINPUT93), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n752), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(G164), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(G164), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n694), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n834), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n836), .A2(new_n832), .A3(new_n693), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n829), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n488), .B(new_n626), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n497), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n693), .B1(new_n836), .B2(new_n832), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n833), .A2(new_n694), .A3(new_n834), .ZN(new_n842));
  INV_X1    g417(.A(new_n829), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n838), .A2(new_n840), .A3(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(G37), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n829), .A2(KEYINPUT95), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n837), .B2(new_n835), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n841), .B(new_n842), .C1(KEYINPUT95), .C2(new_n829), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n845), .B(new_n846), .C1(new_n850), .C2(new_n840), .ZN(new_n851));
  XOR2_X1   g426(.A(KEYINPUT96), .B(KEYINPUT40), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(G395));
  XNOR2_X1  g428(.A(new_n816), .B(new_n621), .ZN(new_n854));
  OAI21_X1  g429(.A(KEYINPUT97), .B1(new_n566), .B2(new_n571), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT97), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n564), .A2(new_n570), .A3(new_n856), .A4(new_n565), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n609), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n572), .A2(new_n856), .A3(new_n608), .A4(new_n607), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OR3_X1    g435(.A1(new_n854), .A2(KEYINPUT98), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(KEYINPUT41), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT41), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n858), .A2(new_n859), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n862), .A2(KEYINPUT99), .A3(new_n864), .ZN(new_n865));
  OR3_X1    g440(.A1(new_n860), .A2(KEYINPUT99), .A3(KEYINPUT41), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n866), .A3(new_n854), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT98), .B1(new_n854), .B2(new_n860), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n861), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT42), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT42), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n861), .A2(new_n867), .A3(new_n871), .A4(new_n868), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n791), .A2(G288), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n766), .A2(G290), .ZN(new_n875));
  OR3_X1    g450(.A1(new_n874), .A2(new_n875), .A3(KEYINPUT100), .ZN(new_n876));
  OAI21_X1  g451(.A(KEYINPUT100), .B1(new_n874), .B2(new_n875), .ZN(new_n877));
  XNOR2_X1  g452(.A(G166), .B(G305), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n878), .A2(new_n877), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n873), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n870), .A2(new_n881), .A3(new_n872), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(G868), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n813), .A2(new_n613), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(G295));
  INV_X1    g463(.A(KEYINPUT101), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n886), .A2(new_n889), .A3(new_n887), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n613), .B1(new_n883), .B2(new_n884), .ZN(new_n891));
  INV_X1    g466(.A(new_n887), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT101), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(new_n893), .ZN(G331));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n879), .A2(new_n880), .A3(KEYINPUT103), .ZN(new_n896));
  AOI21_X1  g471(.A(KEYINPUT103), .B1(new_n879), .B2(new_n880), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(G171), .A2(new_n539), .ZN(new_n899));
  AOI21_X1  g474(.A(G301), .B1(new_n574), .B2(new_n576), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n816), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n899), .A2(new_n900), .A3(new_n816), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n859), .B(new_n858), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n903), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n862), .A2(new_n864), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(new_n906), .A3(new_n901), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n898), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n865), .A2(new_n866), .A3(new_n901), .A4(new_n905), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(new_n881), .A3(new_n904), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n846), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n895), .B1(new_n912), .B2(KEYINPUT43), .ZN(new_n913));
  XOR2_X1   g488(.A(KEYINPUT102), .B(KEYINPUT43), .Z(new_n914));
  NAND2_X1  g489(.A1(new_n910), .A2(new_n904), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n898), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n916), .A2(new_n846), .A3(new_n911), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n913), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n914), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n912), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n916), .A2(new_n846), .A3(new_n914), .A4(new_n911), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(new_n921), .A3(new_n895), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n922), .A2(KEYINPUT104), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(KEYINPUT104), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n918), .B1(new_n923), .B2(new_n924), .ZN(G397));
  INV_X1    g500(.A(G1384), .ZN(new_n926));
  INV_X1    g501(.A(new_n504), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n927), .B1(new_n467), .B2(G126), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n507), .B(new_n509), .C1(new_n928), .C2(new_n462), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n484), .A2(new_n486), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT4), .B1(new_n930), .B2(G138), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n926), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n932), .A2(KEYINPUT105), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(KEYINPUT105), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(KEYINPUT106), .B(G40), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n472), .A2(new_n487), .A3(new_n473), .A4(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n693), .B(G2067), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n941), .A2(new_n942), .A3(new_n939), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n942), .B1(new_n941), .B2(new_n939), .ZN(new_n944));
  INV_X1    g519(.A(G1996), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n752), .B(new_n945), .ZN(new_n946));
  OAI22_X1  g521(.A1(new_n943), .A2(new_n944), .B1(new_n940), .B2(new_n946), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n947), .A2(KEYINPUT108), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(KEYINPUT108), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n785), .A2(new_n787), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G2067), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n694), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n940), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n785), .A2(new_n787), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n939), .B1(new_n950), .B2(new_n955), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n940), .A2(G1986), .A3(G290), .ZN(new_n957));
  XNOR2_X1  g532(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n957), .B(new_n958), .ZN(new_n959));
  AND4_X1   g534(.A1(new_n949), .A2(new_n948), .A3(new_n956), .A4(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n939), .B1(new_n941), .B2(new_n752), .ZN(new_n961));
  XNOR2_X1  g536(.A(KEYINPUT125), .B(KEYINPUT46), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(new_n940), .B2(G1996), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n939), .B(new_n945), .C1(KEYINPUT125), .C2(KEYINPUT46), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n961), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n965), .B(new_n966), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n954), .A2(new_n960), .A3(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n475), .A2(KEYINPUT123), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n472), .A2(KEYINPUT123), .A3(new_n473), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n487), .A2(KEYINPUT53), .A3(G40), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n510), .A2(KEYINPUT45), .A3(new_n926), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n972), .A2(new_n936), .A3(new_n735), .A4(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n932), .A2(KEYINPUT50), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n510), .A2(new_n976), .A3(new_n926), .ZN(new_n977));
  AND4_X1   g552(.A1(new_n472), .A2(new_n487), .A3(new_n473), .A4(new_n937), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n975), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n739), .ZN(new_n980));
  XNOR2_X1  g555(.A(KEYINPUT122), .B(KEYINPUT53), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n932), .A2(new_n934), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n982), .A2(new_n978), .A3(new_n973), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n981), .B1(new_n983), .B2(G2078), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n974), .A2(new_n980), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(G171), .ZN(new_n986));
  INV_X1    g561(.A(new_n983), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n987), .A2(KEYINPUT53), .A3(new_n735), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n988), .A2(G301), .A3(new_n980), .A4(new_n984), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n986), .A2(KEYINPUT54), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT124), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n988), .A2(new_n980), .A3(new_n984), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(G171), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(G171), .B2(new_n985), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT54), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n990), .A2(new_n991), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(new_n987), .B2(G1966), .ZN(new_n999));
  OR2_X1    g574(.A1(new_n979), .A2(G2084), .ZN(new_n1000));
  INV_X1    g575(.A(G1966), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n983), .A2(KEYINPUT114), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n1003), .A2(G8), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n539), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n999), .A2(new_n1000), .A3(G168), .A4(new_n1002), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT121), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(G8), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1007), .A2(KEYINPUT121), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1010), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1006), .A2(G8), .A3(new_n1008), .A4(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1005), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT109), .B(G1971), .Z(new_n1015));
  AND2_X1   g590(.A1(new_n983), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT110), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n983), .A2(new_n1015), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT110), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1017), .B(new_n1020), .C1(G2090), .C2(new_n979), .ZN(new_n1021));
  NAND2_X1  g596(.A1(G303), .A2(G8), .ZN(new_n1022));
  XOR2_X1   g597(.A(new_n1022), .B(KEYINPUT55), .Z(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(G8), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1023), .ZN(new_n1025));
  INV_X1    g600(.A(new_n977), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n976), .B1(new_n510), .B2(new_n926), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1027), .B1(new_n1028), .B2(new_n938), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n975), .A2(KEYINPUT113), .A3(new_n978), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1026), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1016), .B1(new_n722), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G8), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1025), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(G305), .B(G1981), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT49), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n938), .A2(new_n932), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1038), .A2(new_n1033), .ZN(new_n1039));
  OR2_X1    g614(.A1(G305), .A2(G1981), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G305), .A2(G1981), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(KEYINPUT49), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1037), .A2(new_n1039), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT111), .B1(G288), .B2(new_n769), .ZN(new_n1044));
  OR3_X1    g619(.A1(G288), .A2(KEYINPUT111), .A3(new_n769), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1039), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT52), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT52), .B1(G288), .B2(new_n769), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1039), .A2(new_n1044), .A3(new_n1045), .A4(new_n1048), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1043), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1024), .A2(new_n1034), .A3(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n992), .A2(new_n997), .A3(new_n1014), .A4(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT56), .B(G2072), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n987), .A2(new_n1053), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n1028), .A2(new_n1027), .A3(new_n938), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT113), .B1(new_n975), .B2(new_n978), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n977), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1956), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT115), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1031), .A2(new_n1060), .A3(G1956), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1054), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n570), .B1(KEYINPUT117), .B2(KEYINPUT57), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1063), .A2(new_n566), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n566), .A2(KEYINPUT116), .ZN(new_n1065));
  OR2_X1    g640(.A1(new_n570), .A2(KEYINPUT117), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n566), .A2(KEYINPUT116), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .A4(new_n1063), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1064), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1062), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1070), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1072), .B(new_n1054), .C1(new_n1059), .C2(new_n1061), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1071), .A2(KEYINPUT61), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT119), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT61), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n987), .A2(new_n945), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT58), .B(G1341), .Z(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n938), .B2(new_n932), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n553), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1082), .B(KEYINPUT59), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n979), .A2(new_n702), .B1(new_n952), .B2(new_n1038), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT60), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1085), .A2(KEYINPUT120), .A3(new_n609), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n609), .B1(new_n1085), .B2(KEYINPUT120), .ZN(new_n1087));
  OAI22_X1  g662(.A1(new_n1086), .A2(new_n1087), .B1(KEYINPUT120), .B2(new_n1085), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1084), .A2(KEYINPUT60), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1083), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1071), .A2(new_n1091), .A3(KEYINPUT61), .A4(new_n1073), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1075), .A2(new_n1078), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1057), .A2(KEYINPUT115), .A3(new_n1058), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1060), .B1(new_n1031), .B2(G1956), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1094), .A2(new_n1095), .B1(new_n987), .B2(new_n1053), .ZN(new_n1096));
  OAI22_X1  g671(.A1(new_n1096), .A2(new_n1072), .B1(new_n609), .B2(new_n1084), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1097), .A2(new_n1098), .A3(new_n1073), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1098), .B1(new_n1097), .B2(new_n1073), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1052), .B1(new_n1093), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1043), .A2(new_n769), .A3(new_n766), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n1040), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT112), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1104), .B(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n1039), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1050), .A2(G8), .A3(new_n1023), .A4(new_n1021), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT63), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1021), .A2(G8), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1109), .B1(new_n1110), .B2(new_n1025), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1004), .A2(new_n615), .ZN(new_n1112));
  AND4_X1   g687(.A1(new_n1024), .A2(new_n1111), .A3(new_n1112), .A4(new_n1050), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT63), .B1(new_n1051), .B2(new_n1112), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1107), .B(new_n1108), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n994), .B1(new_n1014), .B2(KEYINPUT62), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1005), .A2(new_n1011), .A3(new_n1117), .A4(new_n1013), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1116), .A2(new_n1051), .A3(new_n1118), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1102), .A2(new_n1115), .A3(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(G290), .B(G1986), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n939), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n948), .A2(new_n949), .A3(new_n956), .A4(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n968), .B1(new_n1120), .B2(new_n1123), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g699(.A1(new_n851), .A2(new_n650), .A3(new_n667), .ZN(new_n1126));
  NOR2_X1   g700(.A1(G229), .A2(new_n460), .ZN(new_n1127));
  NAND3_X1  g701(.A1(new_n920), .A2(new_n921), .A3(new_n1127), .ZN(new_n1128));
  NOR2_X1   g702(.A1(new_n1126), .A2(new_n1128), .ZN(G308));
  INV_X1    g703(.A(G308), .ZN(G225));
endmodule


