

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581;

  XOR2_X1 U322 ( .A(n325), .B(n324), .Z(n550) );
  AND2_X1 U323 ( .A1(G232GAT), .A2(G233GAT), .ZN(n290) );
  INV_X1 U324 ( .A(KEYINPUT96), .ZN(n452) );
  INV_X1 U325 ( .A(KEYINPUT97), .ZN(n456) );
  AND2_X1 U326 ( .A1(n385), .A2(n565), .ZN(n386) );
  XNOR2_X1 U327 ( .A(G92GAT), .B(KEYINPUT93), .ZN(n390) );
  XNOR2_X1 U328 ( .A(n314), .B(n290), .ZN(n315) );
  XNOR2_X1 U329 ( .A(n391), .B(n390), .ZN(n392) );
  NOR2_X1 U330 ( .A1(n426), .A2(n540), .ZN(n564) );
  XNOR2_X1 U331 ( .A(n400), .B(n399), .ZN(n401) );
  INV_X1 U332 ( .A(G190GAT), .ZN(n446) );
  XNOR2_X1 U333 ( .A(n402), .B(n401), .ZN(n489) );
  XNOR2_X1 U334 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U335 ( .A(n449), .B(n448), .ZN(G1351GAT) );
  XOR2_X1 U336 ( .A(G204GAT), .B(KEYINPUT86), .Z(n292) );
  XNOR2_X1 U337 ( .A(KEYINPUT88), .B(KEYINPUT24), .ZN(n291) );
  XNOR2_X1 U338 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U339 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n294) );
  XOR2_X1 U340 ( .A(G50GAT), .B(G162GAT), .Z(n314) );
  XOR2_X1 U341 ( .A(G22GAT), .B(G155GAT), .Z(n326) );
  XNOR2_X1 U342 ( .A(n314), .B(n326), .ZN(n293) );
  XNOR2_X1 U343 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U344 ( .A(n296), .B(n295), .Z(n298) );
  NAND2_X1 U345 ( .A1(G228GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n300) );
  XNOR2_X1 U347 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n299) );
  XNOR2_X1 U348 ( .A(n299), .B(KEYINPUT2), .ZN(n416) );
  XOR2_X1 U349 ( .A(n300), .B(n416), .Z(n306) );
  XOR2_X1 U350 ( .A(KEYINPUT87), .B(G218GAT), .Z(n302) );
  XNOR2_X1 U351 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n301) );
  XNOR2_X1 U352 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U353 ( .A(G197GAT), .B(n303), .Z(n398) );
  XNOR2_X1 U354 ( .A(G106GAT), .B(G78GAT), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n304), .B(G148GAT), .ZN(n371) );
  XNOR2_X1 U356 ( .A(n398), .B(n371), .ZN(n305) );
  XNOR2_X1 U357 ( .A(n306), .B(n305), .ZN(n463) );
  XNOR2_X1 U358 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n404) );
  XNOR2_X1 U359 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n389) );
  XOR2_X1 U360 ( .A(KEYINPUT78), .B(KEYINPUT9), .Z(n308) );
  XNOR2_X1 U361 ( .A(G106GAT), .B(KEYINPUT76), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U363 ( .A(G36GAT), .B(G190GAT), .Z(n393) );
  XOR2_X1 U364 ( .A(n309), .B(n393), .Z(n311) );
  XNOR2_X1 U365 ( .A(G134GAT), .B(G218GAT), .ZN(n310) );
  XNOR2_X1 U366 ( .A(n311), .B(n310), .ZN(n317) );
  XOR2_X1 U367 ( .A(G85GAT), .B(G92GAT), .Z(n313) );
  XNOR2_X1 U368 ( .A(G99GAT), .B(KEYINPUT74), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n313), .B(n312), .ZN(n363) );
  XNOR2_X1 U370 ( .A(n363), .B(n315), .ZN(n316) );
  XOR2_X1 U371 ( .A(n317), .B(n316), .Z(n325) );
  XOR2_X1 U372 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n319) );
  XNOR2_X1 U373 ( .A(G43GAT), .B(G29GAT), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U375 ( .A(KEYINPUT70), .B(n320), .Z(n359) );
  XOR2_X1 U376 ( .A(KEYINPUT77), .B(KEYINPUT11), .Z(n322) );
  XNOR2_X1 U377 ( .A(KEYINPUT79), .B(KEYINPUT10), .ZN(n321) );
  XNOR2_X1 U378 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U379 ( .A(n359), .B(n323), .ZN(n324) );
  INV_X1 U380 ( .A(n550), .ZN(n468) );
  XOR2_X1 U381 ( .A(G8GAT), .B(G183GAT), .Z(n391) );
  XOR2_X1 U382 ( .A(n391), .B(n326), .Z(n328) );
  XOR2_X1 U383 ( .A(KEYINPUT71), .B(G1GAT), .Z(n345) );
  XOR2_X1 U384 ( .A(G15GAT), .B(G127GAT), .Z(n435) );
  XNOR2_X1 U385 ( .A(n345), .B(n435), .ZN(n327) );
  XNOR2_X1 U386 ( .A(n328), .B(n327), .ZN(n334) );
  XOR2_X1 U387 ( .A(G57GAT), .B(KEYINPUT72), .Z(n330) );
  XNOR2_X1 U388 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n329) );
  XNOR2_X1 U389 ( .A(n330), .B(n329), .ZN(n370) );
  XOR2_X1 U390 ( .A(n370), .B(KEYINPUT80), .Z(n332) );
  NAND2_X1 U391 ( .A1(G231GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U392 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U393 ( .A(n334), .B(n333), .Z(n342) );
  XOR2_X1 U394 ( .A(KEYINPUT12), .B(G64GAT), .Z(n336) );
  XNOR2_X1 U395 ( .A(G211GAT), .B(G78GAT), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U397 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n338) );
  XNOR2_X1 U398 ( .A(KEYINPUT81), .B(KEYINPUT82), .ZN(n337) );
  XNOR2_X1 U399 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U400 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n342), .B(n341), .ZN(n575) );
  XNOR2_X1 U402 ( .A(KEYINPUT110), .B(KEYINPUT46), .ZN(n376) );
  XOR2_X1 U403 ( .A(KEYINPUT69), .B(KEYINPUT67), .Z(n344) );
  XNOR2_X1 U404 ( .A(KEYINPUT30), .B(KEYINPUT68), .ZN(n343) );
  XNOR2_X1 U405 ( .A(n344), .B(n343), .ZN(n349) );
  XOR2_X1 U406 ( .A(G36GAT), .B(G50GAT), .Z(n347) );
  XNOR2_X1 U407 ( .A(n345), .B(KEYINPUT29), .ZN(n346) );
  XNOR2_X1 U408 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U409 ( .A(n349), .B(n348), .Z(n351) );
  NAND2_X1 U410 ( .A1(G229GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U411 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U412 ( .A(G197GAT), .B(G113GAT), .Z(n353) );
  XNOR2_X1 U413 ( .A(G169GAT), .B(G15GAT), .ZN(n352) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U415 ( .A(n355), .B(n354), .Z(n361) );
  XOR2_X1 U416 ( .A(KEYINPUT66), .B(G8GAT), .Z(n357) );
  XNOR2_X1 U417 ( .A(G141GAT), .B(G22GAT), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U419 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U420 ( .A(n361), .B(n360), .Z(n497) );
  INV_X1 U421 ( .A(n497), .ZN(n565) );
  XNOR2_X1 U422 ( .A(G176GAT), .B(G204GAT), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n362), .B(G64GAT), .ZN(n399) );
  XOR2_X1 U424 ( .A(KEYINPUT31), .B(n363), .Z(n365) );
  NAND2_X1 U425 ( .A1(G230GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n365), .B(n364), .ZN(n369) );
  XOR2_X1 U427 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n367) );
  XNOR2_X1 U428 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U430 ( .A(n369), .B(n368), .Z(n373) );
  XNOR2_X1 U431 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U432 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U433 ( .A(n399), .B(n374), .ZN(n571) );
  XNOR2_X1 U434 ( .A(KEYINPUT41), .B(n571), .ZN(n544) );
  NOR2_X1 U435 ( .A1(n565), .A2(n544), .ZN(n375) );
  XOR2_X1 U436 ( .A(n376), .B(n375), .Z(n377) );
  NAND2_X1 U437 ( .A1(n575), .A2(n377), .ZN(n378) );
  NOR2_X1 U438 ( .A1(n468), .A2(n378), .ZN(n380) );
  XNOR2_X1 U439 ( .A(KEYINPUT111), .B(KEYINPUT47), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n380), .B(n379), .ZN(n387) );
  XNOR2_X1 U441 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n382) );
  XNOR2_X1 U442 ( .A(n550), .B(KEYINPUT36), .ZN(n578) );
  NOR2_X1 U443 ( .A1(n575), .A2(n578), .ZN(n381) );
  XNOR2_X1 U444 ( .A(n382), .B(n381), .ZN(n383) );
  NOR2_X1 U445 ( .A1(n571), .A2(n383), .ZN(n384) );
  XNOR2_X1 U446 ( .A(n384), .B(KEYINPUT112), .ZN(n385) );
  NOR2_X1 U447 ( .A1(n387), .A2(n386), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n538) );
  XOR2_X1 U449 ( .A(n393), .B(n392), .Z(n395) );
  NAND2_X1 U450 ( .A1(G226GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n395), .B(n394), .ZN(n402) );
  XOR2_X1 U452 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n397) );
  XNOR2_X1 U453 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n438) );
  XNOR2_X1 U455 ( .A(n438), .B(n398), .ZN(n400) );
  INV_X1 U456 ( .A(n489), .ZN(n513) );
  NOR2_X1 U457 ( .A1(n538), .A2(n513), .ZN(n403) );
  XNOR2_X1 U458 ( .A(n404), .B(n403), .ZN(n426) );
  XOR2_X1 U459 ( .A(KEYINPUT91), .B(KEYINPUT1), .Z(n406) );
  XNOR2_X1 U460 ( .A(KEYINPUT92), .B(KEYINPUT89), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n425) );
  XOR2_X1 U462 ( .A(G155GAT), .B(G148GAT), .Z(n408) );
  XNOR2_X1 U463 ( .A(G29GAT), .B(G127GAT), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U465 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n410) );
  XNOR2_X1 U466 ( .A(G1GAT), .B(G57GAT), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U468 ( .A(n412), .B(n411), .Z(n418) );
  XOR2_X1 U469 ( .A(G85GAT), .B(G162GAT), .Z(n414) );
  NAND2_X1 U470 ( .A1(G225GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U474 ( .A(n419), .B(KEYINPUT6), .Z(n423) );
  XOR2_X1 U475 ( .A(G120GAT), .B(KEYINPUT0), .Z(n421) );
  XNOR2_X1 U476 ( .A(G113GAT), .B(G134GAT), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n434) );
  XNOR2_X1 U478 ( .A(n434), .B(KEYINPUT90), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n425), .B(n424), .ZN(n510) );
  INV_X1 U481 ( .A(n510), .ZN(n540) );
  NAND2_X1 U482 ( .A1(n463), .A2(n564), .ZN(n427) );
  XNOR2_X1 U483 ( .A(KEYINPUT55), .B(n427), .ZN(n444) );
  XOR2_X1 U484 ( .A(KEYINPUT84), .B(G190GAT), .Z(n429) );
  XNOR2_X1 U485 ( .A(G43GAT), .B(G99GAT), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U487 ( .A(G183GAT), .B(KEYINPUT83), .Z(n431) );
  XNOR2_X1 U488 ( .A(KEYINPUT20), .B(KEYINPUT85), .ZN(n430) );
  XNOR2_X1 U489 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n443) );
  XOR2_X1 U491 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U492 ( .A1(G227GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n437), .B(n436), .ZN(n439) );
  XOR2_X1 U494 ( .A(n439), .B(n438), .Z(n441) );
  XNOR2_X1 U495 ( .A(G176GAT), .B(G71GAT), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U497 ( .A(n443), .B(n442), .Z(n516) );
  INV_X1 U498 ( .A(n516), .ZN(n525) );
  NAND2_X1 U499 ( .A1(n444), .A2(n525), .ZN(n445) );
  XNOR2_X2 U500 ( .A(KEYINPUT120), .B(n445), .ZN(n561) );
  NOR2_X1 U501 ( .A1(n561), .A2(n550), .ZN(n449) );
  XNOR2_X1 U502 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n447) );
  NOR2_X1 U503 ( .A1(n565), .A2(n571), .ZN(n450) );
  XOR2_X1 U504 ( .A(KEYINPUT75), .B(n450), .Z(n485) );
  XNOR2_X1 U505 ( .A(n489), .B(KEYINPUT27), .ZN(n462) );
  NOR2_X1 U506 ( .A1(n463), .A2(n525), .ZN(n451) );
  XNOR2_X1 U507 ( .A(n451), .B(KEYINPUT26), .ZN(n563) );
  NAND2_X1 U508 ( .A1(n462), .A2(n563), .ZN(n537) );
  XNOR2_X1 U509 ( .A(n537), .B(KEYINPUT95), .ZN(n459) );
  NOR2_X1 U510 ( .A1(n513), .A2(n516), .ZN(n453) );
  XNOR2_X1 U511 ( .A(n453), .B(n452), .ZN(n454) );
  NAND2_X1 U512 ( .A1(n454), .A2(n463), .ZN(n455) );
  XNOR2_X1 U513 ( .A(n455), .B(KEYINPUT25), .ZN(n457) );
  XNOR2_X1 U514 ( .A(n457), .B(n456), .ZN(n458) );
  NOR2_X1 U515 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U516 ( .A(n460), .B(KEYINPUT98), .ZN(n461) );
  NOR2_X1 U517 ( .A1(n540), .A2(n461), .ZN(n467) );
  AND2_X1 U518 ( .A1(n540), .A2(n462), .ZN(n464) );
  XOR2_X1 U519 ( .A(n463), .B(KEYINPUT28), .Z(n495) );
  INV_X1 U520 ( .A(n495), .ZN(n519) );
  NAND2_X1 U521 ( .A1(n464), .A2(n519), .ZN(n523) );
  NOR2_X1 U522 ( .A1(n525), .A2(n523), .ZN(n465) );
  XNOR2_X1 U523 ( .A(n465), .B(KEYINPUT94), .ZN(n466) );
  NOR2_X1 U524 ( .A1(n467), .A2(n466), .ZN(n482) );
  NOR2_X1 U525 ( .A1(n468), .A2(n575), .ZN(n469) );
  XOR2_X1 U526 ( .A(KEYINPUT16), .B(n469), .Z(n470) );
  NOR2_X1 U527 ( .A1(n482), .A2(n470), .ZN(n498) );
  NAND2_X1 U528 ( .A1(n485), .A2(n498), .ZN(n478) );
  NOR2_X1 U529 ( .A1(n510), .A2(n478), .ZN(n472) );
  XNOR2_X1 U530 ( .A(KEYINPUT99), .B(KEYINPUT34), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U532 ( .A(G1GAT), .B(n473), .ZN(G1324GAT) );
  NOR2_X1 U533 ( .A1(n513), .A2(n478), .ZN(n474) );
  XOR2_X1 U534 ( .A(G8GAT), .B(n474), .Z(G1325GAT) );
  NOR2_X1 U535 ( .A1(n516), .A2(n478), .ZN(n476) );
  XNOR2_X1 U536 ( .A(KEYINPUT35), .B(KEYINPUT100), .ZN(n475) );
  XNOR2_X1 U537 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U538 ( .A(G15GAT), .B(n477), .ZN(G1326GAT) );
  NOR2_X1 U539 ( .A1(n519), .A2(n478), .ZN(n479) );
  XOR2_X1 U540 ( .A(G22GAT), .B(n479), .Z(G1327GAT) );
  XOR2_X1 U541 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n481) );
  XNOR2_X1 U542 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n480) );
  XNOR2_X1 U543 ( .A(n481), .B(n480), .ZN(n488) );
  NOR2_X1 U544 ( .A1(n578), .A2(n482), .ZN(n483) );
  NAND2_X1 U545 ( .A1(n575), .A2(n483), .ZN(n484) );
  XNOR2_X1 U546 ( .A(KEYINPUT37), .B(n484), .ZN(n509) );
  NAND2_X1 U547 ( .A1(n509), .A2(n485), .ZN(n486) );
  XOR2_X1 U548 ( .A(KEYINPUT38), .B(n486), .Z(n494) );
  NAND2_X1 U549 ( .A1(n494), .A2(n540), .ZN(n487) );
  XOR2_X1 U550 ( .A(n488), .B(n487), .Z(G1328GAT) );
  NAND2_X1 U551 ( .A1(n489), .A2(n494), .ZN(n490) );
  XNOR2_X1 U552 ( .A(G36GAT), .B(n490), .ZN(G1329GAT) );
  NAND2_X1 U553 ( .A1(n494), .A2(n525), .ZN(n492) );
  XOR2_X1 U554 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n493), .ZN(G1330GAT) );
  NAND2_X1 U557 ( .A1(n495), .A2(n494), .ZN(n496) );
  XNOR2_X1 U558 ( .A(G50GAT), .B(n496), .ZN(G1331GAT) );
  XNOR2_X1 U559 ( .A(n544), .B(KEYINPUT104), .ZN(n555) );
  NOR2_X1 U560 ( .A1(n497), .A2(n555), .ZN(n508) );
  NAND2_X1 U561 ( .A1(n508), .A2(n498), .ZN(n504) );
  NOR2_X1 U562 ( .A1(n510), .A2(n504), .ZN(n499) );
  XOR2_X1 U563 ( .A(G57GAT), .B(n499), .Z(n500) );
  XNOR2_X1 U564 ( .A(KEYINPUT42), .B(n500), .ZN(G1332GAT) );
  NOR2_X1 U565 ( .A1(n513), .A2(n504), .ZN(n502) );
  XNOR2_X1 U566 ( .A(G64GAT), .B(KEYINPUT105), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n502), .B(n501), .ZN(G1333GAT) );
  NOR2_X1 U568 ( .A1(n516), .A2(n504), .ZN(n503) );
  XOR2_X1 U569 ( .A(G71GAT), .B(n503), .Z(G1334GAT) );
  NOR2_X1 U570 ( .A1(n519), .A2(n504), .ZN(n506) );
  XNOR2_X1 U571 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U573 ( .A(G78GAT), .B(n507), .ZN(G1335GAT) );
  NAND2_X1 U574 ( .A1(n509), .A2(n508), .ZN(n518) );
  NOR2_X1 U575 ( .A1(n510), .A2(n518), .ZN(n512) );
  XNOR2_X1 U576 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(G1336GAT) );
  NOR2_X1 U578 ( .A1(n513), .A2(n518), .ZN(n514) );
  XOR2_X1 U579 ( .A(KEYINPUT108), .B(n514), .Z(n515) );
  XNOR2_X1 U580 ( .A(G92GAT), .B(n515), .ZN(G1337GAT) );
  NOR2_X1 U581 ( .A1(n516), .A2(n518), .ZN(n517) );
  XOR2_X1 U582 ( .A(G99GAT), .B(n517), .Z(G1338GAT) );
  NOR2_X1 U583 ( .A1(n519), .A2(n518), .ZN(n521) );
  XNOR2_X1 U584 ( .A(KEYINPUT44), .B(KEYINPUT109), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n522), .ZN(G1339GAT) );
  NOR2_X1 U587 ( .A1(n538), .A2(n523), .ZN(n524) );
  NAND2_X1 U588 ( .A1(n525), .A2(n524), .ZN(n533) );
  NOR2_X1 U589 ( .A1(n565), .A2(n533), .ZN(n527) );
  XNOR2_X1 U590 ( .A(G113GAT), .B(KEYINPUT113), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n527), .B(n526), .ZN(G1340GAT) );
  NOR2_X1 U592 ( .A1(n555), .A2(n533), .ZN(n529) );
  XNOR2_X1 U593 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U595 ( .A(G120GAT), .B(n530), .ZN(G1341GAT) );
  NOR2_X1 U596 ( .A1(n575), .A2(n533), .ZN(n531) );
  XOR2_X1 U597 ( .A(KEYINPUT50), .B(n531), .Z(n532) );
  XNOR2_X1 U598 ( .A(G127GAT), .B(n532), .ZN(G1342GAT) );
  NOR2_X1 U599 ( .A1(n550), .A2(n533), .ZN(n535) );
  XNOR2_X1 U600 ( .A(KEYINPUT51), .B(KEYINPUT115), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U602 ( .A(G134GAT), .B(n536), .Z(G1343GAT) );
  NOR2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U604 ( .A1(n540), .A2(n539), .ZN(n549) );
  NOR2_X1 U605 ( .A1(n565), .A2(n549), .ZN(n542) );
  XNOR2_X1 U606 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(n543), .ZN(G1344GAT) );
  NOR2_X1 U609 ( .A1(n544), .A2(n549), .ZN(n546) );
  XNOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(n547), .ZN(G1345GAT) );
  NOR2_X1 U613 ( .A1(n575), .A2(n549), .ZN(n548) );
  XOR2_X1 U614 ( .A(G155GAT), .B(n548), .Z(G1346GAT) );
  NOR2_X1 U615 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U616 ( .A(KEYINPUT118), .B(n551), .Z(n552) );
  XNOR2_X1 U617 ( .A(G162GAT), .B(n552), .ZN(G1347GAT) );
  XNOR2_X1 U618 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n554) );
  NOR2_X1 U619 ( .A1(n565), .A2(n561), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(G1348GAT) );
  NOR2_X1 U621 ( .A1(n561), .A2(n555), .ZN(n560) );
  XOR2_X1 U622 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n557) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(KEYINPUT56), .B(n558), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  NOR2_X1 U627 ( .A1(n575), .A2(n561), .ZN(n562) );
  XOR2_X1 U628 ( .A(G183GAT), .B(n562), .Z(G1350GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n577) );
  NOR2_X1 U630 ( .A1(n565), .A2(n577), .ZN(n570) );
  XOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n567) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(KEYINPUT59), .B(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(G204GAT), .B(KEYINPUT61), .Z(n574) );
  INV_X1 U637 ( .A(n577), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n577), .ZN(n576) );
  XOR2_X1 U641 ( .A(G211GAT), .B(n576), .Z(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

