//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n807,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005;
  INV_X1    g000(.A(G36gat), .ZN(new_n202));
  AND2_X1   g001(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n206), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G50gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G43gat), .ZN(new_n210));
  INV_X1    g009(.A(G43gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G50gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n212), .A3(KEYINPUT15), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n208), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n211), .A2(G50gat), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT15), .B1(new_n216), .B2(KEYINPUT90), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT90), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n210), .A2(new_n212), .A3(new_n218), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n217), .A2(new_n219), .B1(new_n205), .B2(new_n207), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n215), .B1(new_n220), .B2(new_n214), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT91), .B1(new_n221), .B2(KEYINPUT17), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n217), .A2(new_n219), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(new_n208), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(new_n213), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT91), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT17), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n215), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G15gat), .B(G22gat), .ZN(new_n230));
  INV_X1    g029(.A(G1gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT16), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(G1gat), .B2(new_n230), .ZN(new_n234));
  INV_X1    g033(.A(G8gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n234), .B(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT17), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n229), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(KEYINPUT92), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n234), .B(G8gat), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT92), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n213), .B1(new_n205), .B2(new_n207), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n243), .B1(new_n224), .B2(new_n213), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n239), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n238), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G229gat), .A2(G233gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(KEYINPUT18), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n239), .A2(new_n242), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n221), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n245), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n247), .B(KEYINPUT13), .Z(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n238), .A2(new_n247), .A3(new_n245), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT18), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n248), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT89), .ZN(new_n258));
  XNOR2_X1  g057(.A(G113gat), .B(G141gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(G197gat), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT11), .B(G169gat), .Z(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(new_n262), .B(KEYINPUT12), .Z(new_n263));
  NAND2_X1  g062(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n263), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n257), .A2(KEYINPUT89), .A3(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT88), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT30), .ZN(new_n270));
  XNOR2_X1  g069(.A(G8gat), .B(G36gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(G64gat), .B(G92gat), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n271), .B(new_n272), .Z(new_n273));
  INV_X1    g072(.A(G226gat), .ZN(new_n274));
  INV_X1    g073(.A(G233gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G183gat), .A2(G190gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT65), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n279), .A2(G169gat), .A3(G176gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT26), .ZN(new_n281));
  INV_X1    g080(.A(G169gat), .ZN(new_n282));
  INV_X1    g081(.A(G176gat), .ZN(new_n283));
  OAI22_X1  g082(.A1(new_n280), .A2(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n283), .ZN(new_n285));
  NOR3_X1   g084(.A1(new_n285), .A2(new_n279), .A3(KEYINPUT26), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n278), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT66), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT27), .B(G183gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n290), .A2(KEYINPUT64), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT27), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT64), .B1(new_n292), .B2(G183gat), .ZN(new_n293));
  INV_X1    g092(.A(G190gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n289), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n290), .A2(KEYINPUT28), .A3(new_n294), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT66), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n299), .B(new_n278), .C1(new_n284), .C2(new_n286), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n288), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n285), .B(KEYINPUT23), .ZN(new_n302));
  INV_X1    g101(.A(new_n278), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT24), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n303), .A2(new_n304), .B1(G169gat), .B2(G176gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306));
  OR3_X1    g105(.A1(new_n303), .A2(new_n306), .A3(new_n304), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n302), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT25), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n302), .A2(new_n305), .A3(KEYINPUT25), .A4(new_n307), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n301), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n301), .A2(KEYINPUT74), .A3(new_n312), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n277), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G211gat), .B(G218gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n321));
  INV_X1    g120(.A(G197gat), .ZN(new_n322));
  INV_X1    g121(.A(G204gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G197gat), .A2(G204gat), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n321), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n320), .B(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n276), .A2(KEYINPUT29), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NOR3_X1   g129(.A1(new_n317), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n320), .A2(new_n326), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n320), .A2(new_n326), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n315), .A2(new_n328), .A3(new_n316), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n313), .A2(new_n277), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n334), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n273), .B1(new_n331), .B2(new_n338), .ZN(new_n339));
  AND3_X1   g138(.A1(new_n301), .A2(KEYINPUT74), .A3(new_n312), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT74), .B1(new_n301), .B2(new_n312), .ZN(new_n341));
  INV_X1    g140(.A(new_n328), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n327), .B1(new_n343), .B2(new_n336), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n273), .B(KEYINPUT75), .Z(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n276), .B1(new_n340), .B2(new_n341), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(new_n334), .A3(new_n329), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n344), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n270), .B1(new_n339), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n273), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n351), .B1(new_n344), .B2(new_n348), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n352), .A2(KEYINPUT30), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  XOR2_X1   g154(.A(G78gat), .B(G106gat), .Z(new_n356));
  XNOR2_X1  g155(.A(new_n356), .B(KEYINPUT84), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT31), .B(G50gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT2), .ZN(new_n361));
  INV_X1    g160(.A(G155gat), .ZN(new_n362));
  INV_X1    g161(.A(G162gat), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n364), .B1(new_n362), .B2(new_n363), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n366));
  INV_X1    g165(.A(G148gat), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n366), .B1(new_n367), .B2(G141gat), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n369));
  INV_X1    g168(.A(G141gat), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n369), .B1(new_n370), .B2(G148gat), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n367), .A2(KEYINPUT77), .A3(G141gat), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n368), .A2(new_n371), .A3(new_n372), .A4(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n367), .A2(G141gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n370), .A2(G148gat), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n361), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  XOR2_X1   g176(.A(G155gat), .B(G162gat), .Z(new_n378));
  AOI22_X1  g177(.A1(new_n365), .A2(new_n374), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT29), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n334), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT3), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n379), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n379), .A2(new_n382), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n380), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n327), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(G22gat), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(G228gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n389), .A2(new_n275), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT85), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n390), .B1(new_n383), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n382), .B1(new_n327), .B2(KEYINPUT29), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n374), .A2(new_n365), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n378), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(G22gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n398), .A3(new_n386), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n388), .A2(new_n392), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n392), .B1(new_n388), .B2(new_n399), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n360), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n399), .ZN(new_n404));
  INV_X1    g203(.A(new_n392), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n406), .A2(new_n359), .A3(new_n400), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G127gat), .B(G134gat), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT1), .ZN(new_n410));
  INV_X1    g209(.A(G113gat), .ZN(new_n411));
  INV_X1    g210(.A(G120gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G113gat), .A2(G120gat), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n409), .A2(new_n410), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  AND2_X1   g215(.A1(G113gat), .A2(G120gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(G113gat), .A2(G120gat), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT67), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT67), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n413), .A2(new_n420), .A3(new_n414), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n421), .A3(new_n410), .ZN(new_n422));
  INV_X1    g221(.A(new_n409), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT68), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT68), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n422), .A2(new_n426), .A3(new_n423), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n416), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n313), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(G227gat), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n430), .A2(new_n275), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n422), .A2(new_n426), .A3(new_n423), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n426), .B1(new_n422), .B2(new_n423), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n415), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n301), .A2(new_n434), .A3(new_n312), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n429), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT32), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT33), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  XOR2_X1   g238(.A(G15gat), .B(G43gat), .Z(new_n440));
  XNOR2_X1  g239(.A(G71gat), .B(G99gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n437), .A2(new_n439), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n442), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n436), .B(KEYINPUT32), .C1(new_n438), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n431), .B1(new_n429), .B2(new_n435), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT69), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n449), .A2(KEYINPUT34), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(KEYINPUT34), .ZN(new_n452));
  XOR2_X1   g251(.A(new_n452), .B(KEYINPUT70), .Z(new_n453));
  NAND3_X1  g252(.A1(new_n448), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n453), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n455), .B1(new_n447), .B2(new_n450), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n446), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT71), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n443), .A2(new_n445), .B1(new_n454), .B2(new_n456), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT71), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n443), .A2(new_n445), .A3(new_n454), .A4(new_n456), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n408), .A2(new_n459), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT82), .ZN(new_n465));
  XNOR2_X1  g264(.A(G1gat), .B(G29gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(KEYINPUT0), .ZN(new_n467));
  XNOR2_X1  g266(.A(G57gat), .B(G85gat), .ZN(new_n468));
  XOR2_X1   g267(.A(new_n467), .B(new_n468), .Z(new_n469));
  AND3_X1   g268(.A1(new_n394), .A2(new_n415), .A3(new_n395), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n470), .B1(new_n432), .B2(new_n433), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT80), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n434), .A2(new_n396), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n425), .A2(new_n427), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n475), .A2(KEYINPUT80), .A3(new_n470), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(G225gat), .A2(G233gat), .ZN(new_n478));
  XOR2_X1   g277(.A(new_n478), .B(KEYINPUT79), .Z(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT5), .ZN(new_n481));
  INV_X1    g280(.A(new_n479), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n470), .B(KEYINPUT4), .C1(new_n433), .C2(new_n432), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT78), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n379), .B2(new_n382), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n396), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(new_n486), .A3(new_n384), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n482), .B(new_n483), .C1(new_n487), .C2(new_n428), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n394), .A2(new_n395), .A3(new_n415), .ZN(new_n489));
  AOI211_X1 g288(.A(new_n472), .B(new_n489), .C1(new_n425), .C2(new_n427), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT80), .B1(new_n475), .B2(new_n470), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT4), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n488), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n469), .B1(new_n481), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n434), .A2(new_n486), .A3(new_n485), .A4(new_n384), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT5), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n497), .A3(new_n482), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n493), .B1(new_n473), .B2(new_n476), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n471), .A2(new_n493), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT81), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT4), .B1(new_n490), .B2(new_n491), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT81), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(new_n504), .A3(new_n500), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n498), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n465), .B1(new_n495), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n498), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n504), .B1(new_n503), .B2(new_n500), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n499), .A2(KEYINPUT81), .A3(new_n501), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n469), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n497), .B1(new_n477), .B2(new_n479), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n473), .A2(new_n493), .A3(new_n476), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n514), .A2(new_n482), .A3(new_n496), .A4(new_n483), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n512), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n511), .A2(KEYINPUT82), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n507), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT83), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n513), .A2(new_n515), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n512), .B1(new_n506), .B2(new_n522), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n507), .A2(new_n517), .A3(KEYINPUT83), .A4(new_n518), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n523), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT6), .ZN(new_n527));
  AOI211_X1 g326(.A(new_n355), .B(new_n464), .C1(new_n525), .C2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT35), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n269), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n525), .A2(new_n527), .ZN(new_n531));
  INV_X1    g330(.A(new_n464), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(new_n354), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n533), .A2(KEYINPUT88), .A3(KEYINPUT35), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n446), .A2(new_n457), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n536), .A2(new_n460), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n355), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n507), .A2(new_n517), .A3(new_n523), .A4(new_n518), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n527), .ZN(new_n541));
  INV_X1    g340(.A(new_n408), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(KEYINPUT35), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n539), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n535), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT72), .B1(new_n537), .B2(KEYINPUT36), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n459), .A2(new_n462), .A3(KEYINPUT36), .A4(new_n463), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT72), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT36), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n548), .B(new_n549), .C1(new_n536), .C2(new_n460), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n546), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n345), .A2(KEYINPUT38), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n344), .A2(new_n348), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT86), .B(KEYINPUT37), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n552), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n327), .B1(new_n317), .B2(new_n330), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n335), .A2(new_n337), .A3(new_n334), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(KEYINPUT37), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n352), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n527), .A2(new_n540), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT87), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n527), .A2(new_n540), .A3(new_n560), .A4(KEYINPUT87), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT37), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n351), .B1(new_n553), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n554), .B1(new_n344), .B2(new_n348), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT38), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n563), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n492), .A2(new_n482), .A3(new_n474), .ZN(new_n570));
  INV_X1    g369(.A(new_n496), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n571), .B1(new_n502), .B2(new_n505), .ZN(new_n572));
  OAI211_X1 g371(.A(KEYINPUT39), .B(new_n570), .C1(new_n572), .C2(new_n482), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n496), .B1(new_n509), .B2(new_n510), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT39), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(new_n575), .A3(new_n479), .ZN(new_n576));
  AND4_X1   g375(.A1(KEYINPUT40), .A2(new_n573), .A3(new_n469), .A4(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n523), .B1(new_n350), .B2(new_n353), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n573), .A2(new_n576), .A3(new_n469), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT40), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n542), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n551), .B1(new_n569), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n526), .B1(new_n519), .B2(new_n520), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n585), .A2(new_n524), .B1(KEYINPUT6), .B2(new_n526), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n542), .B1(new_n586), .B2(new_n355), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n268), .B1(new_n545), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(KEYINPUT93), .A2(G64gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(KEYINPUT93), .A2(G64gat), .ZN(new_n591));
  OAI21_X1  g390(.A(G57gat), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT94), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT94), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n594), .B(G57gat), .C1(new_n590), .C2(new_n591), .ZN(new_n595));
  INV_X1    g394(.A(G64gat), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n593), .B(new_n595), .C1(G57gat), .C2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G71gat), .A2(G78gat), .ZN(new_n598));
  OR2_X1    g397(.A1(G71gat), .A2(G78gat), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT9), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G57gat), .B(G64gat), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n598), .B(new_n599), .C1(new_n603), .C2(new_n600), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n602), .A2(KEYINPUT21), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n249), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT97), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT97), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n249), .A2(new_n608), .A3(new_n605), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G127gat), .B(G155gat), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT96), .ZN(new_n612));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n613), .B(KEYINPUT95), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n612), .B(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n610), .B(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT21), .B1(new_n602), .B2(new_n604), .ZN(new_n618));
  XOR2_X1   g417(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G183gat), .B(G211gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n617), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G99gat), .B(G106gat), .ZN(new_n624));
  INV_X1    g423(.A(G99gat), .ZN(new_n625));
  INV_X1    g424(.A(G106gat), .ZN(new_n626));
  OAI21_X1  g425(.A(KEYINPUT99), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT99), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n628), .A2(G99gat), .A3(G106gat), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n627), .A2(KEYINPUT8), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(G92gat), .ZN(new_n633));
  INV_X1    g432(.A(G92gat), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n631), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n624), .B1(new_n630), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n637), .A2(KEYINPUT101), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n639));
  AOI211_X1 g438(.A(new_n639), .B(new_n624), .C1(new_n630), .C2(new_n636), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n630), .A2(new_n636), .ZN(new_n643));
  INV_X1    g442(.A(new_n624), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n630), .A2(new_n636), .A3(KEYINPUT100), .A4(new_n624), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI22_X1  g446(.A1(new_n641), .A2(new_n647), .B1(KEYINPUT17), .B2(new_n221), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n648), .A2(KEYINPUT102), .A3(new_n229), .ZN(new_n649));
  AOI21_X1  g448(.A(KEYINPUT102), .B1(new_n648), .B2(new_n229), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n641), .A2(new_n244), .A3(new_n647), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT103), .ZN(new_n652));
  NAND3_X1  g451(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n653));
  AND3_X1   g452(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n652), .B1(new_n651), .B2(new_n653), .ZN(new_n655));
  OAI22_X1  g454(.A1(new_n649), .A2(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G190gat), .B(G218gat), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n657), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n222), .A2(new_n228), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n637), .A2(KEYINPUT101), .ZN(new_n662));
  INV_X1    g461(.A(new_n640), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n647), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n237), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n660), .B1(new_n661), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n648), .A2(new_n229), .A3(KEYINPUT102), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n651), .A2(new_n653), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(KEYINPUT103), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n659), .B1(new_n668), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT98), .ZN(new_n675));
  XNOR2_X1  g474(.A(G134gat), .B(G162gat), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n675), .B(new_n676), .Z(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  OR3_X1    g477(.A1(new_n658), .A2(new_n673), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n668), .A2(new_n659), .A3(new_n672), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n681), .B1(new_n673), .B2(KEYINPUT104), .ZN(new_n682));
  OR3_X1    g481(.A1(new_n656), .A2(KEYINPUT104), .A3(new_n657), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n680), .B1(new_n684), .B2(new_n678), .ZN(new_n685));
  AOI211_X1 g484(.A(KEYINPUT105), .B(new_n677), .C1(new_n682), .C2(new_n683), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n623), .B(new_n679), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT104), .B1(new_n656), .B2(new_n657), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(new_n658), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n656), .A2(KEYINPUT104), .A3(new_n657), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n678), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(KEYINPUT105), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n684), .A2(new_n680), .A3(new_n678), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n696), .A2(KEYINPUT106), .A3(new_n623), .A4(new_n679), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n602), .A2(new_n604), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n664), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n643), .A2(new_n644), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n698), .A2(new_n700), .A3(new_n637), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n699), .A2(new_n701), .A3(KEYINPUT10), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT10), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n664), .A2(new_n698), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(G230gat), .ZN(new_n705));
  OAI22_X1  g504(.A1(new_n702), .A2(new_n704), .B1(new_n705), .B2(new_n275), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n275), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(new_n699), .B2(new_n701), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n708), .A2(KEYINPUT107), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(KEYINPUT107), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n706), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(G120gat), .B(G148gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(G176gat), .B(G204gat), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n712), .B(new_n713), .Z(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n711), .A2(new_n715), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n689), .A2(new_n697), .A3(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n689), .A2(new_n697), .A3(KEYINPUT108), .A4(new_n718), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n589), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n531), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(new_n231), .ZN(G1324gat));
  NOR2_X1   g525(.A1(new_n724), .A2(new_n354), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT109), .B(KEYINPUT16), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(new_n235), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n727), .B2(new_n235), .ZN(new_n731));
  MUX2_X1   g530(.A(new_n730), .B(new_n731), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g531(.A(new_n724), .ZN(new_n733));
  AOI21_X1  g532(.A(G15gat), .B1(new_n733), .B2(new_n537), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n551), .A2(G15gat), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT110), .Z(new_n736));
  AOI21_X1  g535(.A(new_n734), .B1(new_n733), .B2(new_n736), .ZN(G1326gat));
  NAND3_X1  g536(.A1(new_n733), .A2(KEYINPUT111), .A3(new_n542), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n724), .B2(new_n408), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(KEYINPUT43), .B(G22gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1327gat));
  NAND2_X1  g542(.A1(new_n696), .A2(new_n679), .ZN(new_n744));
  INV_X1    g543(.A(new_n544), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n745), .B1(new_n530), .B2(new_n534), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n355), .B1(new_n525), .B2(new_n527), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT112), .B1(new_n747), .B2(new_n408), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n749), .B(new_n542), .C1(new_n586), .C2(new_n355), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n584), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n744), .B1(new_n746), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n588), .ZN(new_n755));
  OAI211_X1 g554(.A(KEYINPUT44), .B(new_n744), .C1(new_n746), .C2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n623), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n718), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n758), .A2(new_n268), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n754), .A2(new_n756), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(G29gat), .B1(new_n760), .B2(new_n531), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n696), .A2(new_n679), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(new_n758), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n589), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n531), .A2(G29gat), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n762), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n589), .A2(KEYINPUT45), .A3(new_n764), .A4(new_n766), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n761), .A2(new_n768), .A3(new_n769), .ZN(G1328gat));
  NOR3_X1   g569(.A1(new_n765), .A2(G36gat), .A3(new_n354), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(KEYINPUT113), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(G36gat), .B1(new_n760), .B2(new_n354), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT113), .B(KEYINPUT46), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n773), .B(new_n774), .C1(new_n771), .C2(new_n775), .ZN(G1329gat));
  OAI21_X1  g575(.A(new_n211), .B1(new_n765), .B2(new_n538), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n551), .A2(G43gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n760), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g579(.A(new_n209), .B1(new_n765), .B2(new_n408), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n542), .A2(G50gat), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n760), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT48), .ZN(G1331gat));
  OR2_X1    g583(.A1(new_n746), .A2(new_n751), .ZN(new_n785));
  INV_X1    g584(.A(new_n718), .ZN(new_n786));
  AND4_X1   g585(.A1(new_n268), .A2(new_n689), .A3(new_n697), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n586), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g590(.A(new_n354), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT114), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n793), .A2(KEYINPUT114), .ZN(new_n796));
  OAI22_X1  g595(.A1(new_n795), .A2(new_n796), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n797));
  INV_X1    g596(.A(new_n796), .ZN(new_n798));
  NOR2_X1   g597(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(new_n794), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n797), .A2(new_n800), .ZN(G1333gat));
  INV_X1    g600(.A(new_n551), .ZN(new_n802));
  OAI21_X1  g601(.A(G71gat), .B1(new_n788), .B2(new_n802), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n538), .A2(G71gat), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n788), .B2(new_n804), .ZN(new_n805));
  XOR2_X1   g604(.A(new_n805), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g605(.A1(new_n788), .A2(new_n408), .ZN(new_n807));
  XOR2_X1   g606(.A(KEYINPUT115), .B(G78gat), .Z(new_n808));
  XNOR2_X1  g607(.A(new_n807), .B(new_n808), .ZN(G1335gat));
  NOR2_X1   g608(.A1(new_n267), .A2(new_n623), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n785), .A2(KEYINPUT51), .A3(new_n744), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT116), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n744), .B(new_n810), .C1(new_n746), .C2(new_n751), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT51), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OR3_X1    g614(.A1(new_n813), .A2(KEYINPUT116), .A3(new_n814), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n812), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n531), .A2(G85gat), .A3(new_n718), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n810), .A2(new_n786), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n754), .A2(new_n756), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(G85gat), .B1(new_n822), .B2(new_n531), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n819), .A2(new_n823), .ZN(G1336gat));
  NOR3_X1   g623(.A1(new_n718), .A2(new_n354), .A3(G92gat), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n817), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n754), .A2(new_n355), .A3(new_n756), .A4(new_n821), .ZN(new_n827));
  AOI21_X1  g626(.A(KEYINPUT52), .B1(new_n827), .B2(G92gat), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n827), .A2(new_n830), .A3(G92gat), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n830), .B1(new_n827), .B2(G92gat), .ZN(new_n832));
  INV_X1    g631(.A(new_n825), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n833), .B1(new_n811), .B2(new_n815), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n831), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n829), .B1(new_n835), .B2(new_n836), .ZN(G1337gat));
  NAND3_X1  g636(.A1(new_n786), .A2(new_n625), .A3(new_n537), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT118), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n817), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(G99gat), .B1(new_n822), .B2(new_n802), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1338gat));
  NOR3_X1   g641(.A1(new_n718), .A2(G106gat), .A3(new_n408), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n817), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n754), .A2(new_n542), .A3(new_n756), .A4(new_n821), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(G106gat), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n811), .A2(new_n815), .ZN(new_n849));
  AOI22_X1  g648(.A1(new_n849), .A2(new_n843), .B1(new_n845), .B2(G106gat), .ZN(new_n850));
  OAI22_X1  g649(.A1(new_n844), .A2(new_n848), .B1(new_n847), .B2(new_n850), .ZN(G1339gat));
  OR3_X1    g650(.A1(new_n699), .A2(KEYINPUT10), .A3(new_n701), .ZN(new_n852));
  INV_X1    g651(.A(new_n704), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n707), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n714), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n852), .A2(new_n707), .A3(new_n853), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n706), .A3(KEYINPUT54), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n856), .A2(KEYINPUT55), .A3(new_n858), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n859), .A2(new_n716), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n246), .A2(new_n247), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n251), .A2(new_n252), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n262), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(new_n257), .B2(new_n263), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n856), .A2(new_n858), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT55), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n864), .A2(new_n865), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n860), .A2(new_n866), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n763), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n864), .B1(new_n716), .B2(new_n717), .ZN(new_n873));
  AND4_X1   g672(.A1(new_n264), .A2(new_n859), .A3(new_n716), .A4(new_n266), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n874), .B2(new_n869), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n875), .A2(new_n744), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n757), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n689), .A2(new_n697), .A3(new_n268), .A4(new_n718), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(KEYINPUT120), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n877), .A2(new_n881), .A3(new_n878), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n883), .A2(new_n586), .A3(new_n408), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n539), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n885), .A2(new_n411), .A3(new_n268), .ZN(new_n886));
  AND4_X1   g685(.A1(new_n354), .A2(new_n459), .A3(new_n462), .A4(new_n463), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n884), .A2(new_n267), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n886), .B1(new_n411), .B2(new_n888), .ZN(G1340gat));
  NOR3_X1   g688(.A1(new_n885), .A2(new_n412), .A3(new_n718), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n884), .A2(new_n786), .A3(new_n887), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n890), .B1(new_n412), .B2(new_n891), .ZN(G1341gat));
  OAI21_X1  g691(.A(G127gat), .B1(new_n885), .B2(new_n757), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n884), .A2(new_n887), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n757), .A2(G127gat), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(G1342gat));
  OAI21_X1  g695(.A(G134gat), .B1(new_n885), .B2(new_n763), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n763), .A2(G134gat), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT56), .B1(new_n894), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n884), .A2(new_n901), .A3(new_n887), .A4(new_n898), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n897), .A2(new_n900), .A3(new_n902), .ZN(G1343gat));
  AOI21_X1  g702(.A(KEYINPUT123), .B1(new_n802), .B2(new_n542), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n551), .A2(new_n905), .A3(new_n408), .ZN(new_n906));
  NOR4_X1   g705(.A1(new_n904), .A2(new_n906), .A3(new_n531), .A4(new_n355), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n880), .A2(new_n907), .A3(new_n882), .ZN(new_n908));
  AOI21_X1  g707(.A(G141gat), .B1(new_n908), .B2(new_n267), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n802), .A2(new_n586), .A3(new_n354), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n880), .A2(new_n542), .A3(new_n882), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT57), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT121), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n914), .B1(new_n867), .B2(new_n868), .ZN(new_n915));
  AOI211_X1 g714(.A(KEYINPUT121), .B(KEYINPUT55), .C1(new_n856), .C2(new_n858), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n873), .B1(new_n917), .B2(new_n874), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n918), .A2(new_n744), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n919), .A2(KEYINPUT122), .B1(new_n763), .B2(new_n871), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n919), .A2(KEYINPUT122), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n757), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n878), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n408), .A2(new_n912), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n910), .B1(new_n913), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n268), .A2(new_n370), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n909), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n929));
  OAI21_X1  g728(.A(KEYINPUT58), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT58), .ZN(new_n931));
  INV_X1    g730(.A(new_n927), .ZN(new_n932));
  AOI211_X1 g731(.A(new_n910), .B(new_n932), .C1(new_n913), .C2(new_n925), .ZN(new_n933));
  OAI211_X1 g732(.A(KEYINPUT124), .B(new_n931), .C1(new_n933), .C2(new_n909), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n930), .A2(new_n934), .ZN(G1344gat));
  NAND3_X1  g734(.A1(new_n908), .A2(new_n367), .A3(new_n786), .ZN(new_n936));
  AOI211_X1 g735(.A(KEYINPUT59), .B(new_n367), .C1(new_n926), .C2(new_n786), .ZN(new_n937));
  XOR2_X1   g736(.A(KEYINPUT125), .B(KEYINPUT59), .Z(new_n938));
  NOR2_X1   g737(.A1(new_n910), .A2(new_n718), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n880), .A2(new_n882), .A3(new_n924), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n721), .A2(new_n268), .A3(new_n722), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n757), .B1(new_n872), .B2(new_n919), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT57), .B1(new_n943), .B2(new_n542), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n940), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI211_X1 g745(.A(KEYINPUT126), .B(KEYINPUT57), .C1(new_n943), .C2(new_n542), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n939), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n938), .B1(new_n948), .B2(G148gat), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n936), .B1(new_n937), .B2(new_n949), .ZN(G1345gat));
  INV_X1    g749(.A(new_n926), .ZN(new_n951));
  OAI21_X1  g750(.A(G155gat), .B1(new_n951), .B2(new_n757), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n908), .A2(new_n362), .A3(new_n623), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1346gat));
  OAI21_X1  g753(.A(G162gat), .B1(new_n951), .B2(new_n763), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n908), .A2(new_n363), .A3(new_n744), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1347gat));
  NOR3_X1   g756(.A1(new_n586), .A2(new_n354), .A3(new_n464), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n883), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(G169gat), .B1(new_n959), .B2(new_n267), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n586), .A2(new_n354), .A3(new_n538), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n883), .A2(new_n408), .A3(new_n961), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n962), .A2(new_n282), .A3(new_n268), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n960), .A2(new_n963), .ZN(G1348gat));
  NAND3_X1  g763(.A1(new_n959), .A2(new_n283), .A3(new_n786), .ZN(new_n965));
  OAI21_X1  g764(.A(G176gat), .B1(new_n962), .B2(new_n718), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(G1349gat));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n623), .A2(new_n290), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n959), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(G183gat), .B1(new_n962), .B2(new_n757), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(KEYINPUT60), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT60), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n970), .A2(new_n974), .A3(new_n971), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n975), .ZN(G1350gat));
  NAND3_X1  g775(.A1(new_n959), .A2(new_n294), .A3(new_n744), .ZN(new_n977));
  OAI21_X1  g776(.A(G190gat), .B1(new_n962), .B2(new_n763), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n978), .A2(KEYINPUT61), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT61), .ZN(new_n980));
  OAI211_X1 g779(.A(new_n980), .B(G190gat), .C1(new_n962), .C2(new_n763), .ZN(new_n981));
  INV_X1    g780(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n977), .B1(new_n979), .B2(new_n982), .ZN(G1351gat));
  NOR3_X1   g782(.A1(new_n551), .A2(new_n586), .A3(new_n354), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n883), .A2(new_n542), .A3(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g785(.A(G197gat), .B1(new_n986), .B2(new_n267), .ZN(new_n987));
  OR2_X1    g786(.A1(new_n946), .A2(new_n947), .ZN(new_n988));
  AND2_X1   g787(.A1(new_n988), .A2(new_n984), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n268), .A2(new_n322), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n987), .B1(new_n989), .B2(new_n990), .ZN(G1352gat));
  NAND3_X1  g790(.A1(new_n988), .A2(new_n786), .A3(new_n984), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(G204gat), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n786), .A2(new_n323), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n985), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g794(.A(new_n995), .B(KEYINPUT62), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n993), .A2(new_n996), .ZN(G1353gat));
  OR3_X1    g796(.A1(new_n985), .A2(G211gat), .A3(new_n757), .ZN(new_n998));
  OAI211_X1 g797(.A(new_n623), .B(new_n984), .C1(new_n946), .C2(new_n947), .ZN(new_n999));
  AND3_X1   g798(.A1(new_n999), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1000));
  AOI21_X1  g799(.A(KEYINPUT63), .B1(new_n999), .B2(G211gat), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n998), .B1(new_n1000), .B2(new_n1001), .ZN(G1354gat));
  NAND3_X1  g801(.A1(new_n988), .A2(new_n744), .A3(new_n984), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(G218gat), .ZN(new_n1004));
  OR3_X1    g803(.A1(new_n985), .A2(G218gat), .A3(new_n763), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(new_n1005), .ZN(G1355gat));
endmodule


