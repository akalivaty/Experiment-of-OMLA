

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U552 ( .A1(n672), .A2(n671), .ZN(n518) );
  INV_X1 U553 ( .A(n682), .ZN(n519) );
  XNOR2_X1 U554 ( .A(n527), .B(KEYINPUT68), .ZN(n528) );
  NOR2_X1 U555 ( .A1(n662), .A2(n803), .ZN(n664) );
  INV_X1 U556 ( .A(KEYINPUT28), .ZN(n663) );
  NAND2_X1 U557 ( .A1(n721), .A2(n522), .ZN(n722) );
  INV_X1 U558 ( .A(KEYINPUT13), .ZN(n627) );
  NAND2_X1 U559 ( .A1(n598), .A2(n597), .ZN(n600) );
  NOR2_X2 U560 ( .A1(n536), .A2(n535), .ZN(G164) );
  XOR2_X1 U561 ( .A(n679), .B(KEYINPUT31), .Z(n520) );
  NOR2_X1 U562 ( .A1(n719), .A2(n700), .ZN(n521) );
  XOR2_X1 U563 ( .A(n720), .B(KEYINPUT100), .Z(n522) );
  XOR2_X1 U564 ( .A(KEYINPUT27), .B(n657), .Z(n523) );
  XOR2_X1 U565 ( .A(G543), .B(KEYINPUT0), .Z(n524) );
  XOR2_X1 U566 ( .A(KEYINPUT104), .B(KEYINPUT32), .Z(n525) );
  NOR2_X1 U567 ( .A1(n961), .A2(n640), .ZN(n652) );
  OR2_X1 U568 ( .A1(n652), .A2(n651), .ZN(n656) );
  XNOR2_X1 U569 ( .A(n674), .B(KEYINPUT30), .ZN(n675) );
  NOR2_X1 U570 ( .A1(n675), .A2(G168), .ZN(n678) );
  NOR2_X1 U571 ( .A1(n678), .A2(n677), .ZN(n679) );
  INV_X1 U572 ( .A(KEYINPUT103), .ZN(n680) );
  XNOR2_X1 U573 ( .A(n690), .B(n525), .ZN(n698) );
  INV_X1 U574 ( .A(KEYINPUT64), .ZN(n702) );
  XNOR2_X1 U575 ( .A(n703), .B(n702), .ZN(n705) );
  NOR2_X1 U576 ( .A1(G164), .A2(G1384), .ZN(n635) );
  INV_X1 U577 ( .A(KEYINPUT17), .ZN(n527) );
  OR2_X1 U578 ( .A1(n723), .A2(n722), .ZN(n736) );
  NOR2_X1 U579 ( .A1(n738), .A2(n737), .ZN(n754) );
  NOR2_X1 U580 ( .A1(n589), .A2(G651), .ZN(n792) );
  XNOR2_X1 U581 ( .A(n600), .B(n599), .ZN(n758) );
  NOR2_X1 U582 ( .A1(n754), .A2(n753), .ZN(n756) );
  NAND2_X1 U583 ( .A1(n633), .A2(n632), .ZN(n961) );
  XOR2_X1 U584 ( .A(KEYINPUT73), .B(n580), .Z(G171) );
  XNOR2_X2 U585 ( .A(G2104), .B(KEYINPUT65), .ZN(n532) );
  AND2_X2 U586 ( .A1(n532), .A2(G2105), .ZN(n889) );
  NAND2_X1 U587 ( .A1(n889), .A2(G126), .ZN(n526) );
  XNOR2_X1 U588 ( .A(n526), .B(KEYINPUT94), .ZN(n531) );
  NOR2_X1 U589 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  XNOR2_X2 U590 ( .A(n529), .B(n528), .ZN(n882) );
  NAND2_X1 U591 ( .A1(G138), .A2(n882), .ZN(n530) );
  NAND2_X1 U592 ( .A1(n531), .A2(n530), .ZN(n536) );
  NOR2_X4 U593 ( .A1(n532), .A2(G2105), .ZN(n881) );
  NAND2_X1 U594 ( .A1(G102), .A2(n881), .ZN(n534) );
  AND2_X1 U595 ( .A1(G2105), .A2(G2104), .ZN(n886) );
  NAND2_X1 U596 ( .A1(G114), .A2(n886), .ZN(n533) );
  NAND2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U598 ( .A1(G543), .A2(G651), .ZN(n787) );
  NAND2_X1 U599 ( .A1(n787), .A2(G89), .ZN(n537) );
  XNOR2_X1 U600 ( .A(n537), .B(KEYINPUT4), .ZN(n540) );
  XOR2_X1 U601 ( .A(KEYINPUT69), .B(n524), .Z(n589) );
  INV_X1 U602 ( .A(G651), .ZN(n542) );
  NOR2_X1 U603 ( .A1(n589), .A2(n542), .ZN(n538) );
  XNOR2_X2 U604 ( .A(n538), .B(KEYINPUT70), .ZN(n788) );
  NAND2_X1 U605 ( .A1(G76), .A2(n788), .ZN(n539) );
  NAND2_X1 U606 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n541), .B(KEYINPUT5), .ZN(n548) );
  NOR2_X1 U608 ( .A1(G543), .A2(n542), .ZN(n543) );
  XOR2_X1 U609 ( .A(KEYINPUT1), .B(n543), .Z(n791) );
  NAND2_X1 U610 ( .A1(G63), .A2(n791), .ZN(n545) );
  NAND2_X1 U611 ( .A1(G51), .A2(n792), .ZN(n544) );
  NAND2_X1 U612 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U613 ( .A(KEYINPUT6), .B(n546), .Z(n547) );
  NAND2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n549), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U616 ( .A1(n791), .A2(G60), .ZN(n550) );
  XOR2_X1 U617 ( .A(KEYINPUT71), .B(n550), .Z(n552) );
  NAND2_X1 U618 ( .A1(n792), .A2(G47), .ZN(n551) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U620 ( .A(KEYINPUT72), .B(n553), .Z(n557) );
  NAND2_X1 U621 ( .A1(n788), .A2(G72), .ZN(n555) );
  NAND2_X1 U622 ( .A1(G85), .A2(n787), .ZN(n554) );
  AND2_X1 U623 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(G290) );
  NAND2_X1 U625 ( .A1(n791), .A2(G61), .ZN(n559) );
  NAND2_X1 U626 ( .A1(n787), .A2(G86), .ZN(n558) );
  NAND2_X1 U627 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U628 ( .A(KEYINPUT88), .B(n560), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n788), .A2(G73), .ZN(n561) );
  XOR2_X1 U630 ( .A(KEYINPUT2), .B(n561), .Z(n562) );
  NOR2_X1 U631 ( .A1(n563), .A2(n562), .ZN(n565) );
  NAND2_X1 U632 ( .A1(n792), .A2(G48), .ZN(n564) );
  NAND2_X1 U633 ( .A1(n565), .A2(n564), .ZN(G305) );
  NAND2_X1 U634 ( .A1(G91), .A2(n787), .ZN(n567) );
  NAND2_X1 U635 ( .A1(G78), .A2(n788), .ZN(n566) );
  NAND2_X1 U636 ( .A1(n567), .A2(n566), .ZN(n570) );
  NAND2_X1 U637 ( .A1(n792), .A2(G53), .ZN(n568) );
  XOR2_X1 U638 ( .A(KEYINPUT74), .B(n568), .Z(n569) );
  NOR2_X1 U639 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n791), .A2(G65), .ZN(n571) );
  NAND2_X1 U641 ( .A1(n572), .A2(n571), .ZN(G299) );
  NAND2_X1 U642 ( .A1(G64), .A2(n791), .ZN(n574) );
  NAND2_X1 U643 ( .A1(G52), .A2(n792), .ZN(n573) );
  NAND2_X1 U644 ( .A1(n574), .A2(n573), .ZN(n579) );
  NAND2_X1 U645 ( .A1(G90), .A2(n787), .ZN(n576) );
  NAND2_X1 U646 ( .A1(G77), .A2(n788), .ZN(n575) );
  NAND2_X1 U647 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U648 ( .A(KEYINPUT9), .B(n577), .Z(n578) );
  NOR2_X1 U649 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U650 ( .A(G168), .B(KEYINPUT8), .Z(n581) );
  XNOR2_X1 U651 ( .A(KEYINPUT82), .B(n581), .ZN(G286) );
  NAND2_X1 U652 ( .A1(G75), .A2(n788), .ZN(n584) );
  NAND2_X1 U653 ( .A1(G88), .A2(n787), .ZN(n582) );
  XOR2_X1 U654 ( .A(KEYINPUT89), .B(n582), .Z(n583) );
  NAND2_X1 U655 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U656 ( .A1(G62), .A2(n791), .ZN(n586) );
  NAND2_X1 U657 ( .A1(G50), .A2(n792), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U659 ( .A1(n588), .A2(n587), .ZN(G166) );
  INV_X1 U660 ( .A(G166), .ZN(G303) );
  NAND2_X1 U661 ( .A1(G651), .A2(G74), .ZN(n594) );
  NAND2_X1 U662 ( .A1(G49), .A2(n792), .ZN(n591) );
  NAND2_X1 U663 ( .A1(G87), .A2(n589), .ZN(n590) );
  NAND2_X1 U664 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U665 ( .A1(n791), .A2(n592), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U667 ( .A(KEYINPUT87), .B(n595), .Z(G288) );
  NAND2_X1 U668 ( .A1(n881), .A2(G101), .ZN(n596) );
  XOR2_X1 U669 ( .A(n596), .B(KEYINPUT23), .Z(n598) );
  NAND2_X1 U670 ( .A1(n889), .A2(G125), .ZN(n597) );
  INV_X1 U671 ( .A(KEYINPUT66), .ZN(n599) );
  NAND2_X1 U672 ( .A1(G137), .A2(n882), .ZN(n757) );
  NAND2_X1 U673 ( .A1(G113), .A2(n886), .ZN(n601) );
  XOR2_X1 U674 ( .A(KEYINPUT67), .B(n601), .Z(n759) );
  AND2_X1 U675 ( .A1(n759), .A2(G40), .ZN(n602) );
  AND2_X1 U676 ( .A1(n757), .A2(n602), .ZN(n634) );
  NAND2_X1 U677 ( .A1(n758), .A2(n634), .ZN(n603) );
  NOR2_X1 U678 ( .A1(n635), .A2(n603), .ZN(n750) );
  XNOR2_X1 U679 ( .A(G1986), .B(G290), .ZN(n958) );
  NAND2_X1 U680 ( .A1(n750), .A2(n958), .ZN(n622) );
  NAND2_X1 U681 ( .A1(G119), .A2(n889), .ZN(n605) );
  NAND2_X1 U682 ( .A1(G131), .A2(n882), .ZN(n604) );
  NAND2_X1 U683 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U684 ( .A1(G95), .A2(n881), .ZN(n607) );
  NAND2_X1 U685 ( .A1(G107), .A2(n886), .ZN(n606) );
  NAND2_X1 U686 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U687 ( .A1(n609), .A2(n608), .ZN(n901) );
  INV_X1 U688 ( .A(G1991), .ZN(n1005) );
  NOR2_X1 U689 ( .A1(n901), .A2(n1005), .ZN(n619) );
  XOR2_X1 U690 ( .A(KEYINPUT38), .B(KEYINPUT98), .Z(n611) );
  NAND2_X1 U691 ( .A1(G105), .A2(n881), .ZN(n610) );
  XNOR2_X1 U692 ( .A(n611), .B(n610), .ZN(n615) );
  NAND2_X1 U693 ( .A1(G117), .A2(n886), .ZN(n613) );
  NAND2_X1 U694 ( .A1(G141), .A2(n882), .ZN(n612) );
  NAND2_X1 U695 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U696 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U697 ( .A1(n889), .A2(G129), .ZN(n616) );
  NAND2_X1 U698 ( .A1(n617), .A2(n616), .ZN(n872) );
  AND2_X1 U699 ( .A1(n872), .A2(G1996), .ZN(n618) );
  NOR2_X1 U700 ( .A1(n619), .A2(n618), .ZN(n934) );
  XNOR2_X1 U701 ( .A(KEYINPUT99), .B(n750), .ZN(n620) );
  NOR2_X1 U702 ( .A1(n934), .A2(n620), .ZN(n742) );
  INV_X1 U703 ( .A(n742), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n738) );
  XNOR2_X1 U705 ( .A(G1981), .B(G305), .ZN(n947) );
  NAND2_X1 U706 ( .A1(n791), .A2(G56), .ZN(n623) );
  XOR2_X1 U707 ( .A(KEYINPUT14), .B(n623), .Z(n630) );
  NAND2_X1 U708 ( .A1(G68), .A2(n788), .ZN(n626) );
  NAND2_X1 U709 ( .A1(n787), .A2(G81), .ZN(n624) );
  XNOR2_X1 U710 ( .A(n624), .B(KEYINPUT12), .ZN(n625) );
  NAND2_X1 U711 ( .A1(n626), .A2(n625), .ZN(n628) );
  XNOR2_X1 U712 ( .A(n628), .B(n627), .ZN(n629) );
  NOR2_X1 U713 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U714 ( .A(n631), .B(KEYINPUT78), .ZN(n633) );
  NAND2_X1 U715 ( .A1(G43), .A2(n792), .ZN(n632) );
  AND2_X1 U716 ( .A1(n758), .A2(n634), .ZN(n636) );
  NAND2_X2 U717 ( .A1(n636), .A2(n635), .ZN(n682) );
  AND2_X1 U718 ( .A1(n519), .A2(G1996), .ZN(n637) );
  XOR2_X1 U719 ( .A(n637), .B(KEYINPUT26), .Z(n639) );
  NAND2_X1 U720 ( .A1(n682), .A2(G1341), .ZN(n638) );
  NAND2_X1 U721 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U722 ( .A1(n792), .A2(G54), .ZN(n647) );
  NAND2_X1 U723 ( .A1(G92), .A2(n787), .ZN(n642) );
  NAND2_X1 U724 ( .A1(G66), .A2(n791), .ZN(n641) );
  NAND2_X1 U725 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U726 ( .A1(G79), .A2(n788), .ZN(n643) );
  XNOR2_X1 U727 ( .A(KEYINPUT81), .B(n643), .ZN(n644) );
  NOR2_X1 U728 ( .A1(n645), .A2(n644), .ZN(n646) );
  AND2_X1 U729 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U730 ( .A(KEYINPUT15), .B(n648), .ZN(n653) );
  NAND2_X1 U731 ( .A1(G1348), .A2(n682), .ZN(n650) );
  NAND2_X1 U732 ( .A1(n519), .A2(G2067), .ZN(n649) );
  NAND2_X1 U733 ( .A1(n650), .A2(n649), .ZN(n654) );
  NOR2_X1 U734 ( .A1(n653), .A2(n654), .ZN(n651) );
  INV_X1 U735 ( .A(n653), .ZN(n908) );
  NAND2_X1 U736 ( .A1(n653), .A2(n654), .ZN(n655) );
  NAND2_X1 U737 ( .A1(n656), .A2(n655), .ZN(n661) );
  INV_X1 U738 ( .A(G299), .ZN(n803) );
  NAND2_X1 U739 ( .A1(n682), .A2(G1956), .ZN(n658) );
  NAND2_X1 U740 ( .A1(n519), .A2(G2072), .ZN(n657) );
  NAND2_X1 U741 ( .A1(n658), .A2(n523), .ZN(n659) );
  XNOR2_X1 U742 ( .A(n659), .B(KEYINPUT101), .ZN(n662) );
  NAND2_X1 U743 ( .A1(n803), .A2(n662), .ZN(n660) );
  NAND2_X1 U744 ( .A1(n661), .A2(n660), .ZN(n666) );
  XNOR2_X1 U745 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U746 ( .A1(n666), .A2(n665), .ZN(n668) );
  XNOR2_X1 U747 ( .A(KEYINPUT29), .B(KEYINPUT102), .ZN(n667) );
  XNOR2_X1 U748 ( .A(n668), .B(n667), .ZN(n672) );
  XNOR2_X1 U749 ( .A(G2078), .B(KEYINPUT25), .ZN(n1001) );
  NOR2_X1 U750 ( .A1(n682), .A2(n1001), .ZN(n670) );
  AND2_X1 U751 ( .A1(n682), .A2(G1961), .ZN(n669) );
  NOR2_X1 U752 ( .A1(n670), .A2(n669), .ZN(n676) );
  AND2_X1 U753 ( .A1(G171), .A2(n676), .ZN(n671) );
  NAND2_X1 U754 ( .A1(G8), .A2(n682), .ZN(n719) );
  NOR2_X1 U755 ( .A1(G1966), .A2(n719), .ZN(n694) );
  NOR2_X1 U756 ( .A1(G2084), .A2(n682), .ZN(n691) );
  NOR2_X1 U757 ( .A1(n694), .A2(n691), .ZN(n673) );
  NAND2_X1 U758 ( .A1(G8), .A2(n673), .ZN(n674) );
  NOR2_X1 U759 ( .A1(G171), .A2(n676), .ZN(n677) );
  XNOR2_X1 U760 ( .A(n520), .B(n680), .ZN(n681) );
  NAND2_X1 U761 ( .A1(n518), .A2(n681), .ZN(n692) );
  NAND2_X1 U762 ( .A1(n692), .A2(G286), .ZN(n689) );
  INV_X1 U763 ( .A(G8), .ZN(n687) );
  NOR2_X1 U764 ( .A1(G1971), .A2(n719), .ZN(n684) );
  NOR2_X1 U765 ( .A1(G2090), .A2(n682), .ZN(n683) );
  NOR2_X1 U766 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U767 ( .A1(n685), .A2(G303), .ZN(n686) );
  OR2_X1 U768 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U769 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U770 ( .A1(n691), .A2(G8), .ZN(n696) );
  INV_X1 U771 ( .A(n692), .ZN(n693) );
  NOR2_X1 U772 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U773 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U774 ( .A1(n698), .A2(n697), .ZN(n713) );
  NOR2_X1 U775 ( .A1(G1976), .A2(G288), .ZN(n706) );
  NOR2_X1 U776 ( .A1(G1971), .A2(G303), .ZN(n699) );
  NOR2_X1 U777 ( .A1(n706), .A2(n699), .ZN(n950) );
  NAND2_X1 U778 ( .A1(n713), .A2(n950), .ZN(n701) );
  NAND2_X1 U779 ( .A1(G1976), .A2(G288), .ZN(n949) );
  INV_X1 U780 ( .A(n949), .ZN(n700) );
  NAND2_X1 U781 ( .A1(n701), .A2(n521), .ZN(n703) );
  INV_X1 U782 ( .A(KEYINPUT33), .ZN(n704) );
  NAND2_X1 U783 ( .A1(n705), .A2(n704), .ZN(n710) );
  INV_X1 U784 ( .A(n719), .ZN(n707) );
  NAND2_X1 U785 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U786 ( .A1(n708), .A2(KEYINPUT33), .ZN(n709) );
  NAND2_X1 U787 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U788 ( .A(KEYINPUT105), .B(n711), .ZN(n712) );
  NOR2_X1 U789 ( .A1(n947), .A2(n712), .ZN(n723) );
  NOR2_X1 U790 ( .A1(G2090), .A2(G303), .ZN(n714) );
  NAND2_X1 U791 ( .A1(G8), .A2(n714), .ZN(n715) );
  NAND2_X1 U792 ( .A1(n713), .A2(n715), .ZN(n716) );
  NAND2_X1 U793 ( .A1(n716), .A2(n719), .ZN(n721) );
  NOR2_X1 U794 ( .A1(G1981), .A2(G305), .ZN(n717) );
  XOR2_X1 U795 ( .A(n717), .B(KEYINPUT24), .Z(n718) );
  NOR2_X1 U796 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U797 ( .A(G2067), .B(KEYINPUT37), .ZN(n748) );
  XNOR2_X1 U798 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n728) );
  NAND2_X1 U799 ( .A1(G128), .A2(n889), .ZN(n725) );
  NAND2_X1 U800 ( .A1(G116), .A2(n886), .ZN(n724) );
  NAND2_X1 U801 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U802 ( .A(n726), .B(KEYINPUT35), .ZN(n727) );
  XNOR2_X1 U803 ( .A(n728), .B(n727), .ZN(n734) );
  NAND2_X1 U804 ( .A1(G140), .A2(n882), .ZN(n729) );
  XOR2_X1 U805 ( .A(KEYINPUT95), .B(n729), .Z(n731) );
  NAND2_X1 U806 ( .A1(n881), .A2(G104), .ZN(n730) );
  NAND2_X1 U807 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U808 ( .A(KEYINPUT34), .B(n732), .ZN(n733) );
  NOR2_X1 U809 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U810 ( .A(KEYINPUT36), .B(n735), .ZN(n904) );
  NOR2_X1 U811 ( .A1(n748), .A2(n904), .ZN(n940) );
  NAND2_X1 U812 ( .A1(n750), .A2(n940), .ZN(n747) );
  NAND2_X1 U813 ( .A1(n736), .A2(n747), .ZN(n737) );
  NOR2_X1 U814 ( .A1(G1996), .A2(n872), .ZN(n920) );
  AND2_X1 U815 ( .A1(n1005), .A2(n901), .ZN(n932) );
  NOR2_X1 U816 ( .A1(G1986), .A2(G290), .ZN(n739) );
  XNOR2_X1 U817 ( .A(KEYINPUT106), .B(n739), .ZN(n740) );
  NOR2_X1 U818 ( .A1(n932), .A2(n740), .ZN(n741) );
  NOR2_X1 U819 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U820 ( .A1(n920), .A2(n743), .ZN(n744) );
  XOR2_X1 U821 ( .A(n744), .B(KEYINPUT39), .Z(n745) );
  XNOR2_X1 U822 ( .A(KEYINPUT107), .B(n745), .ZN(n746) );
  NAND2_X1 U823 ( .A1(n747), .A2(n746), .ZN(n749) );
  NAND2_X1 U824 ( .A1(n748), .A2(n904), .ZN(n937) );
  NAND2_X1 U825 ( .A1(n749), .A2(n937), .ZN(n751) );
  NAND2_X1 U826 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U827 ( .A(KEYINPUT108), .B(n752), .Z(n753) );
  INV_X1 U828 ( .A(KEYINPUT40), .ZN(n755) );
  XNOR2_X1 U829 ( .A(n756), .B(n755), .ZN(G329) );
  AND2_X1 U830 ( .A1(n758), .A2(n757), .ZN(n760) );
  AND2_X1 U831 ( .A1(n760), .A2(n759), .ZN(G160) );
  AND2_X1 U832 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U833 ( .A1(n882), .A2(G135), .ZN(n767) );
  NAND2_X1 U834 ( .A1(G99), .A2(n881), .ZN(n762) );
  NAND2_X1 U835 ( .A1(G111), .A2(n886), .ZN(n761) );
  NAND2_X1 U836 ( .A1(n762), .A2(n761), .ZN(n765) );
  NAND2_X1 U837 ( .A1(n889), .A2(G123), .ZN(n763) );
  XOR2_X1 U838 ( .A(KEYINPUT18), .B(n763), .Z(n764) );
  NOR2_X1 U839 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U840 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U841 ( .A(n768), .B(KEYINPUT84), .ZN(n929) );
  XNOR2_X1 U842 ( .A(n929), .B(G2096), .ZN(n769) );
  OR2_X1 U843 ( .A1(G2100), .A2(n769), .ZN(G156) );
  INV_X1 U844 ( .A(G57), .ZN(G237) );
  INV_X1 U845 ( .A(G132), .ZN(G219) );
  INV_X1 U846 ( .A(G82), .ZN(G220) );
  XOR2_X1 U847 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n771) );
  NAND2_X1 U848 ( .A1(G7), .A2(G661), .ZN(n770) );
  XNOR2_X1 U849 ( .A(n771), .B(n770), .ZN(G223) );
  XOR2_X1 U850 ( .A(KEYINPUT77), .B(KEYINPUT11), .Z(n773) );
  INV_X1 U851 ( .A(G223), .ZN(n840) );
  NAND2_X1 U852 ( .A1(G567), .A2(n840), .ZN(n772) );
  XNOR2_X1 U853 ( .A(n773), .B(n772), .ZN(n774) );
  XOR2_X1 U854 ( .A(KEYINPUT76), .B(n774), .Z(G234) );
  INV_X1 U855 ( .A(G860), .ZN(n781) );
  OR2_X1 U856 ( .A1(n961), .A2(n781), .ZN(G153) );
  XNOR2_X1 U857 ( .A(G171), .B(KEYINPUT79), .ZN(G301) );
  NAND2_X1 U858 ( .A1(G868), .A2(G301), .ZN(n775) );
  XNOR2_X1 U859 ( .A(n775), .B(KEYINPUT80), .ZN(n777) );
  INV_X1 U860 ( .A(G868), .ZN(n801) );
  NAND2_X1 U861 ( .A1(n801), .A2(n653), .ZN(n776) );
  NAND2_X1 U862 ( .A1(n777), .A2(n776), .ZN(G284) );
  NOR2_X1 U863 ( .A1(G286), .A2(n801), .ZN(n778) );
  XOR2_X1 U864 ( .A(KEYINPUT83), .B(n778), .Z(n780) );
  NOR2_X1 U865 ( .A1(G868), .A2(G299), .ZN(n779) );
  NOR2_X1 U866 ( .A1(n780), .A2(n779), .ZN(G297) );
  NAND2_X1 U867 ( .A1(n781), .A2(G559), .ZN(n782) );
  NAND2_X1 U868 ( .A1(n782), .A2(n908), .ZN(n783) );
  XNOR2_X1 U869 ( .A(n783), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U870 ( .A1(G868), .A2(n961), .ZN(n786) );
  NAND2_X1 U871 ( .A1(n908), .A2(G868), .ZN(n784) );
  NOR2_X1 U872 ( .A1(G559), .A2(n784), .ZN(n785) );
  NOR2_X1 U873 ( .A1(n786), .A2(n785), .ZN(G282) );
  NAND2_X1 U874 ( .A1(G93), .A2(n787), .ZN(n790) );
  NAND2_X1 U875 ( .A1(G80), .A2(n788), .ZN(n789) );
  NAND2_X1 U876 ( .A1(n790), .A2(n789), .ZN(n796) );
  NAND2_X1 U877 ( .A1(G67), .A2(n791), .ZN(n794) );
  NAND2_X1 U878 ( .A1(G55), .A2(n792), .ZN(n793) );
  NAND2_X1 U879 ( .A1(n794), .A2(n793), .ZN(n795) );
  OR2_X1 U880 ( .A1(n796), .A2(n795), .ZN(n806) );
  NAND2_X1 U881 ( .A1(G559), .A2(n908), .ZN(n797) );
  XOR2_X1 U882 ( .A(n961), .B(n797), .Z(n810) );
  XNOR2_X1 U883 ( .A(KEYINPUT85), .B(n810), .ZN(n798) );
  NOR2_X1 U884 ( .A1(G860), .A2(n798), .ZN(n799) );
  XOR2_X1 U885 ( .A(n806), .B(n799), .Z(n800) );
  XNOR2_X1 U886 ( .A(n800), .B(KEYINPUT86), .ZN(G145) );
  NAND2_X1 U887 ( .A1(n801), .A2(n806), .ZN(n802) );
  XNOR2_X1 U888 ( .A(n802), .B(KEYINPUT90), .ZN(n813) );
  XNOR2_X1 U889 ( .A(G290), .B(KEYINPUT19), .ZN(n805) );
  XNOR2_X1 U890 ( .A(G166), .B(n803), .ZN(n804) );
  XNOR2_X1 U891 ( .A(n805), .B(n804), .ZN(n809) );
  XNOR2_X1 U892 ( .A(n806), .B(G305), .ZN(n807) );
  XNOR2_X1 U893 ( .A(G288), .B(n807), .ZN(n808) );
  XNOR2_X1 U894 ( .A(n809), .B(n808), .ZN(n907) );
  XNOR2_X1 U895 ( .A(n907), .B(n810), .ZN(n811) );
  NAND2_X1 U896 ( .A1(G868), .A2(n811), .ZN(n812) );
  NAND2_X1 U897 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U898 ( .A(KEYINPUT91), .B(n814), .Z(G295) );
  NAND2_X1 U899 ( .A1(G2078), .A2(G2084), .ZN(n816) );
  XOR2_X1 U900 ( .A(KEYINPUT92), .B(KEYINPUT20), .Z(n815) );
  XNOR2_X1 U901 ( .A(n816), .B(n815), .ZN(n817) );
  NAND2_X1 U902 ( .A1(G2090), .A2(n817), .ZN(n818) );
  XNOR2_X1 U903 ( .A(KEYINPUT21), .B(n818), .ZN(n819) );
  NAND2_X1 U904 ( .A1(n819), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U905 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U906 ( .A1(G220), .A2(G219), .ZN(n820) );
  XOR2_X1 U907 ( .A(KEYINPUT22), .B(n820), .Z(n821) );
  NOR2_X1 U908 ( .A1(G218), .A2(n821), .ZN(n822) );
  NAND2_X1 U909 ( .A1(G96), .A2(n822), .ZN(n845) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n845), .ZN(n826) );
  NAND2_X1 U911 ( .A1(G69), .A2(G120), .ZN(n823) );
  NOR2_X1 U912 ( .A1(G237), .A2(n823), .ZN(n824) );
  NAND2_X1 U913 ( .A1(G108), .A2(n824), .ZN(n846) );
  NAND2_X1 U914 ( .A1(G567), .A2(n846), .ZN(n825) );
  NAND2_X1 U915 ( .A1(n826), .A2(n825), .ZN(n847) );
  NAND2_X1 U916 ( .A1(G661), .A2(G483), .ZN(n827) );
  NOR2_X1 U917 ( .A1(n847), .A2(n827), .ZN(n844) );
  NAND2_X1 U918 ( .A1(G36), .A2(n844), .ZN(n828) );
  XOR2_X1 U919 ( .A(KEYINPUT93), .B(n828), .Z(G176) );
  XNOR2_X1 U920 ( .A(G2427), .B(G2451), .ZN(n838) );
  XOR2_X1 U921 ( .A(G2430), .B(G2443), .Z(n830) );
  XNOR2_X1 U922 ( .A(KEYINPUT109), .B(G2438), .ZN(n829) );
  XNOR2_X1 U923 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U924 ( .A(G2435), .B(G2454), .Z(n832) );
  XNOR2_X1 U925 ( .A(G1341), .B(G1348), .ZN(n831) );
  XNOR2_X1 U926 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U927 ( .A(n834), .B(n833), .Z(n836) );
  XNOR2_X1 U928 ( .A(KEYINPUT110), .B(G2446), .ZN(n835) );
  XNOR2_X1 U929 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U930 ( .A(n838), .B(n837), .ZN(n839) );
  NAND2_X1 U931 ( .A1(n839), .A2(G14), .ZN(n913) );
  XNOR2_X1 U932 ( .A(KEYINPUT111), .B(n913), .ZN(G401) );
  NAND2_X1 U933 ( .A1(n840), .A2(G2106), .ZN(n841) );
  XNOR2_X1 U934 ( .A(n841), .B(KEYINPUT112), .ZN(G217) );
  AND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n842) );
  NAND2_X1 U936 ( .A1(G661), .A2(n842), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n843) );
  NAND2_X1 U938 ( .A1(n844), .A2(n843), .ZN(G188) );
  INV_X1 U940 ( .A(G120), .ZN(G236) );
  INV_X1 U941 ( .A(G96), .ZN(G221) );
  INV_X1 U942 ( .A(G69), .ZN(G235) );
  NOR2_X1 U943 ( .A1(n846), .A2(n845), .ZN(G325) );
  INV_X1 U944 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U945 ( .A(KEYINPUT113), .B(n847), .ZN(G319) );
  XOR2_X1 U946 ( .A(G2100), .B(G2096), .Z(n849) );
  XNOR2_X1 U947 ( .A(KEYINPUT42), .B(G2678), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U949 ( .A(KEYINPUT43), .B(G2072), .Z(n851) );
  XNOR2_X1 U950 ( .A(G2090), .B(G2067), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U952 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2084), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(G227) );
  XOR2_X1 U955 ( .A(G1986), .B(G1961), .Z(n857) );
  XNOR2_X1 U956 ( .A(G1976), .B(G1971), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U958 ( .A(n858), .B(KEYINPUT41), .Z(n860) );
  XNOR2_X1 U959 ( .A(G1981), .B(G1966), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U961 ( .A(G2474), .B(G1991), .Z(n862) );
  XNOR2_X1 U962 ( .A(G1996), .B(G1956), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(G229) );
  NAND2_X1 U965 ( .A1(G112), .A2(n886), .ZN(n866) );
  NAND2_X1 U966 ( .A1(G136), .A2(n882), .ZN(n865) );
  NAND2_X1 U967 ( .A1(n866), .A2(n865), .ZN(n871) );
  NAND2_X1 U968 ( .A1(G124), .A2(n889), .ZN(n867) );
  XNOR2_X1 U969 ( .A(n867), .B(KEYINPUT44), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n881), .A2(G100), .ZN(n868) );
  NAND2_X1 U971 ( .A1(n869), .A2(n868), .ZN(n870) );
  NOR2_X1 U972 ( .A1(n871), .A2(n870), .ZN(G162) );
  XOR2_X1 U973 ( .A(G160), .B(n872), .Z(n880) );
  NAND2_X1 U974 ( .A1(G103), .A2(n881), .ZN(n874) );
  NAND2_X1 U975 ( .A1(G139), .A2(n882), .ZN(n873) );
  NAND2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n879) );
  NAND2_X1 U977 ( .A1(G127), .A2(n889), .ZN(n876) );
  NAND2_X1 U978 ( .A1(G115), .A2(n886), .ZN(n875) );
  NAND2_X1 U979 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U980 ( .A(KEYINPUT47), .B(n877), .Z(n878) );
  NOR2_X1 U981 ( .A1(n879), .A2(n878), .ZN(n922) );
  XNOR2_X1 U982 ( .A(n880), .B(n922), .ZN(n894) );
  NAND2_X1 U983 ( .A1(G106), .A2(n881), .ZN(n884) );
  NAND2_X1 U984 ( .A1(G142), .A2(n882), .ZN(n883) );
  NAND2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U986 ( .A(n885), .B(KEYINPUT45), .ZN(n888) );
  NAND2_X1 U987 ( .A1(G118), .A2(n886), .ZN(n887) );
  NAND2_X1 U988 ( .A1(n888), .A2(n887), .ZN(n892) );
  NAND2_X1 U989 ( .A1(n889), .A2(G130), .ZN(n890) );
  XOR2_X1 U990 ( .A(KEYINPUT114), .B(n890), .Z(n891) );
  NOR2_X1 U991 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U992 ( .A(n894), .B(n893), .Z(n896) );
  XNOR2_X1 U993 ( .A(G164), .B(G162), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n900) );
  XOR2_X1 U995 ( .A(KEYINPUT116), .B(KEYINPUT115), .Z(n898) );
  XNOR2_X1 U996 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n897) );
  XNOR2_X1 U997 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U998 ( .A(n900), .B(n899), .Z(n903) );
  XNOR2_X1 U999 ( .A(n901), .B(n929), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n905) );
  XOR2_X1 U1001 ( .A(n905), .B(n904), .Z(n906) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n906), .ZN(G395) );
  XNOR2_X1 U1003 ( .A(n908), .B(n907), .ZN(n910) );
  XNOR2_X1 U1004 ( .A(G286), .B(G171), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(n911), .B(n961), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n912), .ZN(G397) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n913), .ZN(n916) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(n914), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1013 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1016 ( .A(G2090), .B(G162), .Z(n919) );
  NOR2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1018 ( .A(KEYINPUT51), .B(n921), .Z(n928) );
  XNOR2_X1 U1019 ( .A(KEYINPUT117), .B(KEYINPUT50), .ZN(n926) );
  XNOR2_X1 U1020 ( .A(G2072), .B(n922), .ZN(n924) );
  XNOR2_X1 U1021 ( .A(G164), .B(G2078), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(n926), .B(n925), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n936) );
  XNOR2_X1 U1025 ( .A(G160), .B(G2084), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n938) );
  NAND2_X1 U1030 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1031 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1032 ( .A(KEYINPUT52), .B(n941), .ZN(n943) );
  INV_X1 U1033 ( .A(KEYINPUT55), .ZN(n942) );
  NAND2_X1 U1034 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1035 ( .A1(n944), .A2(G29), .ZN(n1025) );
  INV_X1 U1036 ( .A(G16), .ZN(n992) );
  XOR2_X1 U1037 ( .A(KEYINPUT56), .B(KEYINPUT124), .Z(n945) );
  XNOR2_X1 U1038 ( .A(n992), .B(n945), .ZN(n967) );
  XOR2_X1 U1039 ( .A(G168), .B(G1966), .Z(n946) );
  NOR2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1041 ( .A(KEYINPUT57), .B(n948), .Z(n965) );
  XNOR2_X1 U1042 ( .A(G171), .B(G1961), .ZN(n960) );
  AND2_X1 U1043 ( .A1(G303), .A2(G1971), .ZN(n952) );
  NAND2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n956) );
  XNOR2_X1 U1046 ( .A(n653), .B(G1348), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(G299), .B(G1956), .ZN(n953) );
  NOR2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1050 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1051 ( .A1(n960), .A2(n959), .ZN(n963) );
  XNOR2_X1 U1052 ( .A(G1341), .B(n961), .ZN(n962) );
  NOR2_X1 U1053 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1054 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1055 ( .A1(n967), .A2(n966), .ZN(n994) );
  XNOR2_X1 U1056 ( .A(G1976), .B(G23), .ZN(n969) );
  XNOR2_X1 U1057 ( .A(G1971), .B(G22), .ZN(n968) );
  NOR2_X1 U1058 ( .A1(n969), .A2(n968), .ZN(n971) );
  XOR2_X1 U1059 ( .A(G1986), .B(G24), .Z(n970) );
  NAND2_X1 U1060 ( .A1(n971), .A2(n970), .ZN(n973) );
  XOR2_X1 U1061 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n972) );
  XNOR2_X1 U1062 ( .A(n973), .B(n972), .ZN(n977) );
  XNOR2_X1 U1063 ( .A(G1961), .B(G5), .ZN(n975) );
  XNOR2_X1 U1064 ( .A(G1966), .B(G21), .ZN(n974) );
  NOR2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1066 ( .A1(n977), .A2(n976), .ZN(n988) );
  XNOR2_X1 U1067 ( .A(G1956), .B(G20), .ZN(n982) );
  XNOR2_X1 U1068 ( .A(G1981), .B(G6), .ZN(n979) );
  XNOR2_X1 U1069 ( .A(G1341), .B(G19), .ZN(n978) );
  NOR2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1071 ( .A(KEYINPUT125), .B(n980), .ZN(n981) );
  NOR2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n985) );
  XNOR2_X1 U1073 ( .A(G1348), .B(KEYINPUT59), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(n983), .B(G4), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(KEYINPUT60), .B(n986), .ZN(n987) );
  NOR2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1078 ( .A(n989), .B(KEYINPUT127), .Z(n990) );
  XNOR2_X1 U1079 ( .A(KEYINPUT61), .B(n990), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1081 ( .A1(n994), .A2(n993), .ZN(n1023) );
  XOR2_X1 U1082 ( .A(G2084), .B(G34), .Z(n995) );
  XNOR2_X1 U1083 ( .A(KEYINPUT54), .B(n995), .ZN(n1014) );
  XNOR2_X1 U1084 ( .A(G2090), .B(G35), .ZN(n1012) );
  XOR2_X1 U1085 ( .A(G2067), .B(G26), .Z(n998) );
  XOR2_X1 U1086 ( .A(G33), .B(KEYINPUT118), .Z(n996) );
  XNOR2_X1 U1087 ( .A(n996), .B(G2072), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(KEYINPUT119), .B(n999), .ZN(n1000) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(G28), .ZN(n1009) );
  XOR2_X1 U1091 ( .A(n1001), .B(G27), .Z(n1003) );
  XNOR2_X1 U1092 ( .A(G32), .B(G1996), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(KEYINPUT120), .B(n1004), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(n1005), .B(G25), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(KEYINPUT53), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(n1015), .B(KEYINPUT122), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(n1017), .B(n1016), .ZN(n1019) );
  INV_X1 U1104 ( .A(G29), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(G11), .ZN(n1021) );
  XOR2_X1 U1107 ( .A(KEYINPUT123), .B(n1021), .Z(n1022) );
  NOR2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1026), .Z(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

