//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n831, new_n832, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946;
  XNOR2_X1  g000(.A(G141gat), .B(G148gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  AOI21_X1  g002(.A(new_n202), .B1(KEYINPUT2), .B2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G155gat), .ZN(new_n205));
  INV_X1    g004(.A(G162gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(new_n203), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n204), .A2(new_n208), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n203), .B(new_n207), .C1(new_n202), .C2(KEYINPUT2), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(G113gat), .B(G120gat), .Z(new_n212));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G127gat), .B(G134gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n212), .A2(new_n213), .A3(new_n215), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n211), .B(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT5), .ZN(new_n221));
  NAND2_X1  g020(.A1(G225gat), .A2(G233gat), .ZN(new_n222));
  NOR3_X1   g021(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OR3_X1    g022(.A1(new_n211), .A2(KEYINPUT81), .A3(KEYINPUT3), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT81), .B1(new_n211), .B2(KEYINPUT3), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n219), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n227), .B1(KEYINPUT3), .B2(new_n211), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n221), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT72), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n219), .B(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n211), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT4), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n227), .ZN(new_n235));
  OAI22_X1  g034(.A1(new_n234), .A2(KEYINPUT82), .B1(KEYINPUT4), .B2(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n234), .A2(KEYINPUT82), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n229), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n222), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n226), .A2(new_n228), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n232), .A2(KEYINPUT4), .A3(new_n227), .ZN(new_n241));
  INV_X1    g040(.A(new_n233), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n240), .B(new_n241), .C1(new_n242), .C2(KEYINPUT4), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n239), .B1(new_n243), .B2(new_n221), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n223), .B1(new_n238), .B2(new_n244), .ZN(new_n245));
  XOR2_X1   g044(.A(G1gat), .B(G29gat), .Z(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(G85gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT0), .B(G57gat), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n247), .B(new_n248), .Z(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  OR2_X1    g049(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT6), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n245), .A2(new_n250), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT83), .ZN(new_n255));
  OR2_X1    g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n245), .A2(new_n250), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT6), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n255), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(G169gat), .A2(G176gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT23), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT65), .ZN(new_n263));
  INV_X1    g062(.A(G169gat), .ZN(new_n264));
  INV_X1    g063(.A(G176gat), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT23), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n265), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT24), .ZN(new_n272));
  INV_X1    g071(.A(G183gat), .ZN(new_n273));
  INV_X1    g072(.A(G190gat), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n269), .A2(new_n270), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n275), .B(new_n276), .C1(G183gat), .C2(G190gat), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n263), .B(new_n268), .C1(new_n271), .C2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT25), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n268), .A2(KEYINPUT25), .A3(new_n262), .ZN(new_n281));
  AND2_X1   g080(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n269), .B(new_n275), .C1(new_n284), .C2(G190gat), .ZN(new_n285));
  AND3_X1   g084(.A1(new_n281), .A2(KEYINPUT67), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT67), .B1(new_n281), .B2(new_n285), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n280), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT27), .ZN(new_n289));
  AOI21_X1  g088(.A(G190gat), .B1(new_n289), .B2(G183gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT66), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n273), .ZN(new_n292));
  NAND2_X1  g091(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n289), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT68), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n290), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n295), .B(KEYINPUT27), .C1(new_n282), .C2(new_n283), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT69), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT28), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT27), .B1(new_n282), .B2(new_n283), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT68), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT69), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n302), .A2(new_n303), .A3(new_n297), .A4(new_n290), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n299), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n273), .A2(new_n274), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT27), .B(G183gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(new_n274), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n306), .B1(new_n308), .B2(KEYINPUT28), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n310));
  OR3_X1    g109(.A1(new_n310), .A2(new_n261), .A3(KEYINPUT70), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT70), .B1(new_n310), .B2(new_n261), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n267), .A2(KEYINPUT26), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n305), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n288), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G226gat), .A2(G233gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n302), .A2(new_n297), .A3(new_n290), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT28), .B1(new_n321), .B2(KEYINPUT69), .ZN(new_n322));
  AOI211_X1 g121(.A(KEYINPUT71), .B(new_n315), .C1(new_n322), .C2(new_n304), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT71), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n324), .B1(new_n305), .B2(new_n316), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n288), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT79), .B(KEYINPUT29), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n327), .B1(G226gat), .B2(G233gat), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n320), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G197gat), .B(G204gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT22), .ZN(new_n331));
  INV_X1    g130(.A(G211gat), .ZN(new_n332));
  INV_X1    g131(.A(G218gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G211gat), .B(G218gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n329), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT29), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n318), .A2(new_n339), .A3(new_n319), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n340), .B1(new_n326), .B2(new_n319), .ZN(new_n341));
  INV_X1    g140(.A(new_n337), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G8gat), .B(G36gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(G64gat), .B(G92gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n348), .A2(KEYINPUT80), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(KEYINPUT80), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT30), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n348), .A2(KEYINPUT30), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n344), .A2(new_n347), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n260), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G228gat), .A2(G233gat), .ZN(new_n358));
  INV_X1    g157(.A(new_n327), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n342), .B1(new_n226), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT84), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n337), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n336), .A2(new_n330), .A3(new_n334), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n362), .B(new_n359), .C1(new_n361), .C2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT3), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n232), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n358), .B1(new_n360), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT3), .B1(new_n342), .B2(new_n339), .ZN(new_n368));
  OAI211_X1 g167(.A(G228gat), .B(G233gat), .C1(new_n368), .C2(new_n232), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n367), .B1(new_n360), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT85), .B1(new_n370), .B2(G22gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(G78gat), .B(G106gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT31), .B(G50gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n370), .B(G22gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n357), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n243), .A2(new_n239), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n250), .B1(new_n380), .B2(KEYINPUT39), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT39), .B1(new_n220), .B2(new_n239), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n382), .B1(new_n243), .B2(new_n239), .ZN(new_n383));
  OR2_X1    g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT40), .ZN(new_n385));
  OR3_X1    g184(.A1(new_n384), .A2(KEYINPUT88), .A3(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT88), .B1(new_n384), .B2(new_n385), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n384), .A2(new_n385), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n389), .A2(KEYINPUT87), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(KEYINPUT87), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n388), .A2(new_n251), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT86), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n393), .B1(new_n352), .B2(new_n355), .ZN(new_n394));
  INV_X1    g193(.A(new_n355), .ZN(new_n395));
  INV_X1    g194(.A(new_n351), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n396), .A2(new_n349), .ZN(new_n397));
  OAI211_X1 g196(.A(KEYINPUT86), .B(new_n395), .C1(new_n397), .C2(KEYINPUT30), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n392), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT38), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT37), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n401), .B1(new_n341), .B2(new_n337), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n329), .A2(new_n342), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(new_n404), .B(KEYINPUT90), .Z(new_n405));
  NAND3_X1  g204(.A1(new_n338), .A2(new_n401), .A3(new_n343), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n347), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n400), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n344), .A2(KEYINPUT37), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n409), .A2(KEYINPUT38), .A3(new_n347), .A4(new_n406), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT89), .ZN(new_n413));
  INV_X1    g212(.A(new_n253), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n252), .B1(new_n245), .B2(new_n250), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n251), .A2(KEYINPUT89), .A3(new_n252), .A4(new_n253), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n397), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT91), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n257), .B2(KEYINPUT6), .ZN(new_n421));
  NOR4_X1   g220(.A1(new_n245), .A2(KEYINPUT91), .A3(new_n252), .A4(new_n250), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n418), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n377), .B1(new_n412), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n379), .B1(new_n399), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n219), .B(KEYINPUT72), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n326), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(G227gat), .ZN(new_n429));
  INV_X1    g228(.A(G233gat), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n231), .B(new_n288), .C1(new_n323), .C2(new_n325), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n428), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  XOR2_X1   g233(.A(new_n434), .B(KEYINPUT34), .Z(new_n435));
  AOI21_X1  g234(.A(new_n432), .B1(new_n428), .B2(new_n433), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT32), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(G15gat), .B(G43gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(G71gat), .B(G99gat), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n439), .B(new_n440), .Z(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT33), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT74), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n436), .A2(KEYINPUT73), .A3(KEYINPUT33), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n441), .B1(new_n436), .B2(new_n437), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT73), .B1(new_n436), .B2(KEYINPUT33), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n444), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n441), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n317), .A2(KEYINPUT71), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n305), .A2(new_n324), .A3(new_n316), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n231), .B1(new_n453), .B2(new_n288), .ZN(new_n454));
  INV_X1    g253(.A(new_n433), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n431), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n450), .B1(new_n456), .B2(KEYINPUT32), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT73), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT33), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n456), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n457), .A2(new_n460), .A3(new_n448), .A4(new_n444), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n435), .B(new_n443), .C1(new_n449), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT75), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n457), .A2(new_n448), .A3(new_n460), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT74), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n466), .A2(new_n461), .B1(new_n438), .B2(new_n442), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n467), .A2(new_n435), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n443), .B1(new_n449), .B2(new_n462), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT75), .ZN(new_n471));
  INV_X1    g270(.A(new_n435), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT36), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT76), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n471), .B1(new_n467), .B2(new_n435), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n470), .A2(new_n472), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n473), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(KEYINPUT76), .A3(KEYINPUT36), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT77), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n479), .A2(new_n484), .A3(new_n463), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT36), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n470), .A2(KEYINPUT77), .A3(new_n472), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT78), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT78), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n485), .A2(new_n487), .A3(new_n490), .A4(new_n486), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n426), .B1(new_n483), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n377), .B1(new_n469), .B2(new_n474), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT92), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT92), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n496), .A3(new_n377), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT35), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n357), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n495), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n378), .B1(new_n485), .B2(new_n487), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n418), .A2(new_n423), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n394), .A2(new_n398), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n498), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n493), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(G229gat), .A2(G233gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(G43gat), .B(G50gat), .ZN(new_n509));
  NOR2_X1   g308(.A1(G29gat), .A2(G36gat), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT14), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XOR2_X1   g311(.A(new_n512), .B(KEYINPUT93), .Z(new_n513));
  XOR2_X1   g312(.A(KEYINPUT94), .B(G36gat), .Z(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(G29gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT95), .ZN(new_n516));
  OAI211_X1 g315(.A(KEYINPUT15), .B(new_n509), .C1(new_n513), .C2(new_n516), .ZN(new_n517));
  OR3_X1    g316(.A1(new_n509), .A2(KEYINPUT96), .A3(KEYINPUT15), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n509), .A2(KEYINPUT15), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT96), .B1(new_n509), .B2(KEYINPUT15), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n518), .A2(new_n519), .A3(new_n512), .A4(new_n520), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(G8gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT16), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n525), .B1(new_n526), .B2(G1gat), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n524), .B1(new_n527), .B2(KEYINPUT97), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n527), .B1(G1gat), .B2(new_n525), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n528), .B(new_n529), .Z(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n523), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n530), .B1(new_n523), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT17), .B1(new_n517), .B2(new_n522), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n508), .B(new_n532), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT18), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n523), .B(new_n531), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n508), .B(KEYINPUT13), .Z(new_n540));
  AOI22_X1  g339(.A1(new_n536), .A2(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G113gat), .B(G141gat), .ZN(new_n543));
  INV_X1    g342(.A(G197gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT11), .B(G169gat), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n545), .B(new_n546), .Z(new_n547));
  XOR2_X1   g346(.A(new_n547), .B(KEYINPUT12), .Z(new_n548));
  OR2_X1    g347(.A1(new_n542), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n538), .A2(new_n541), .A3(new_n548), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT98), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n538), .A2(new_n541), .A3(KEYINPUT98), .A4(new_n548), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n507), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT9), .ZN(new_n558));
  INV_X1    g357(.A(G71gat), .ZN(new_n559));
  INV_X1    g358(.A(G78gat), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT99), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n562), .ZN(new_n564));
  XOR2_X1   g363(.A(G57gat), .B(G64gat), .Z(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G71gat), .B(G78gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(KEYINPUT100), .B(KEYINPUT21), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(G127gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(new_n205), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n575));
  XNOR2_X1  g374(.A(G183gat), .B(G211gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n574), .B(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n531), .B1(KEYINPUT21), .B2(new_n568), .ZN(new_n579));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n580), .B(KEYINPUT101), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n579), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n578), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT7), .ZN(new_n584));
  NAND2_X1  g383(.A1(G85gat), .A2(G92gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  AOI22_X1  g385(.A1(new_n584), .A2(new_n585), .B1(new_n586), .B2(KEYINPUT8), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT102), .B(G85gat), .ZN(new_n588));
  OAI221_X1 g387(.A(new_n587), .B1(new_n584), .B2(new_n585), .C1(G92gat), .C2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT103), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(G99gat), .B(G106gat), .Z(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n589), .B(KEYINPUT103), .ZN(new_n594));
  INV_X1    g393(.A(new_n592), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n533), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(new_n523), .ZN(new_n599));
  AND2_X1   g398(.A1(G232gat), .A2(G233gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n599), .B1(KEYINPUT41), .B2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n600), .B(KEYINPUT41), .Z(new_n602));
  OAI21_X1  g401(.A(new_n601), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G134gat), .B(G162gat), .Z(new_n604));
  XNOR2_X1  g403(.A(G190gat), .B(G218gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n603), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n583), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n594), .A2(new_n595), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n591), .A2(new_n592), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n568), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n593), .A2(new_n596), .A3(new_n569), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(KEYINPUT104), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT104), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n611), .A2(new_n616), .A3(new_n612), .A4(new_n613), .ZN(new_n617));
  INV_X1    g416(.A(new_n611), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT10), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n615), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G230gat), .A2(G233gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n611), .A2(new_n613), .ZN(new_n623));
  INV_X1    g422(.A(new_n621), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G120gat), .B(G148gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(G176gat), .B(G204gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n629), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n622), .A2(new_n625), .A3(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n608), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n557), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n260), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G1gat), .ZN(G1324gat));
  INV_X1    g439(.A(new_n394), .ZN(new_n641));
  INV_X1    g440(.A(new_n398), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n636), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(KEYINPUT42), .B1(new_n644), .B2(new_n524), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT16), .B(G8gat), .Z(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  MUX2_X1   g446(.A(KEYINPUT42), .B(new_n645), .S(new_n647), .Z(G1325gat));
  INV_X1    g447(.A(G15gat), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n488), .A2(KEYINPUT78), .ZN(new_n650));
  INV_X1    g449(.A(new_n491), .ZN(new_n651));
  AOI21_X1  g450(.A(KEYINPUT76), .B1(new_n481), .B2(KEYINPUT36), .ZN(new_n652));
  AOI211_X1 g451(.A(new_n476), .B(new_n486), .C1(new_n480), .C2(new_n473), .ZN(new_n653));
  OAI22_X1  g452(.A1(new_n650), .A2(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n636), .A2(new_n649), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n485), .A2(new_n487), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n637), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n655), .B1(new_n649), .B2(new_n657), .ZN(G1326gat));
  OR3_X1    g457(.A1(new_n636), .A2(KEYINPUT105), .A3(new_n377), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT105), .B1(new_n636), .B2(new_n377), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT43), .B(G22gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1327gat));
  NOR3_X1   g462(.A1(new_n583), .A2(new_n634), .A3(new_n607), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n557), .A2(new_n664), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n665), .A2(G29gat), .A3(new_n260), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n666), .B(KEYINPUT45), .Z(new_n667));
  INV_X1    g466(.A(new_n607), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n668), .B1(new_n493), .B2(new_n506), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT108), .B(KEYINPUT44), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  AOI22_X1  g471(.A1(new_n477), .A2(new_n482), .B1(new_n489), .B2(new_n491), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n505), .B(new_n500), .C1(new_n673), .C2(new_n426), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(KEYINPUT108), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n674), .A2(new_n668), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n633), .B(KEYINPUT107), .Z(new_n680));
  NAND2_X1  g479(.A1(new_n555), .A2(KEYINPUT106), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n549), .A2(new_n554), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n680), .A2(new_n685), .A3(new_n583), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n679), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(G29gat), .B1(new_n687), .B2(new_n260), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n667), .A2(new_n688), .ZN(G1328gat));
  NOR3_X1   g488(.A1(new_n665), .A2(new_n514), .A3(new_n643), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT46), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n514), .B1(new_n687), .B2(new_n643), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(G1329gat));
  OAI21_X1  g492(.A(G43gat), .B1(new_n687), .B2(new_n654), .ZN(new_n694));
  INV_X1    g493(.A(new_n665), .ZN(new_n695));
  INV_X1    g494(.A(G43gat), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(new_n696), .A3(new_n656), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n694), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n698), .B1(new_n694), .B2(new_n697), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(G1330gat));
  OAI21_X1  g500(.A(G50gat), .B1(new_n687), .B2(new_n377), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n377), .A2(G50gat), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT48), .ZN(new_n704));
  AOI22_X1  g503(.A1(new_n695), .A2(new_n703), .B1(KEYINPUT110), .B2(new_n704), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n704), .A2(KEYINPUT110), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n702), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n706), .B1(new_n702), .B2(new_n705), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(G1331gat));
  INV_X1    g508(.A(new_n680), .ZN(new_n710));
  NOR4_X1   g509(.A1(new_n507), .A2(new_n608), .A3(new_n684), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n638), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(G57gat), .ZN(G1332gat));
  INV_X1    g512(.A(KEYINPUT111), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n643), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT49), .B(G64gat), .Z(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n716), .B2(new_n718), .ZN(G1333gat));
  AOI21_X1  g518(.A(G71gat), .B1(new_n711), .B2(new_n656), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n654), .A2(new_n559), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n720), .B1(new_n711), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT50), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1334gat));
  NAND2_X1  g523(.A1(new_n711), .A2(new_n378), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g525(.A1(new_n684), .A2(new_n583), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n633), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n679), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n588), .B1(new_n730), .B2(new_n260), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n668), .B(new_n727), .C1(new_n493), .C2(new_n506), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT51), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n260), .A2(new_n588), .A3(new_n633), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT112), .Z(new_n735));
  OAI21_X1  g534(.A(new_n731), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT113), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT113), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n731), .B(new_n738), .C1(new_n733), .C2(new_n735), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(G1336gat));
  INV_X1    g539(.A(new_n733), .ZN(new_n741));
  INV_X1    g540(.A(new_n715), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n742), .A2(G92gat), .A3(new_n710), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT52), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n729), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n745), .B1(new_n672), .B2(new_n678), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n746), .A2(KEYINPUT116), .A3(new_n715), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G92gat), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT116), .B1(new_n746), .B2(new_n715), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n744), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n643), .ZN(new_n751));
  INV_X1    g550(.A(new_n426), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n654), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT35), .B1(new_n501), .B2(new_n503), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n496), .B1(new_n481), .B2(new_n377), .ZN(new_n755));
  AOI211_X1 g554(.A(KEYINPUT92), .B(new_n378), .C1(new_n480), .C2(new_n473), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n754), .B1(new_n757), .B2(new_n499), .ZN(new_n758));
  AOI211_X1 g557(.A(new_n607), .B(new_n676), .C1(new_n753), .C2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n670), .B1(new_n674), .B2(new_n668), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n751), .B(new_n729), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G92gat), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT114), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n732), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n674), .A2(new_n668), .A3(new_n727), .A4(new_n764), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n743), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n762), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT115), .B1(new_n770), .B2(KEYINPUT52), .ZN(new_n771));
  AOI22_X1  g570(.A1(new_n761), .A2(G92gat), .B1(new_n743), .B2(new_n768), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n750), .B1(new_n771), .B2(new_n775), .ZN(G1337gat));
  OAI21_X1  g575(.A(G99gat), .B1(new_n730), .B2(new_n654), .ZN(new_n777));
  INV_X1    g576(.A(G99gat), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n656), .A2(new_n778), .A3(new_n634), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n777), .B1(new_n733), .B2(new_n779), .ZN(G1338gat));
  INV_X1    g579(.A(G106gat), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n746), .B2(new_n378), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n710), .A2(G106gat), .A3(new_n377), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n768), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785));
  INV_X1    g584(.A(new_n783), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n733), .B2(new_n786), .ZN(new_n787));
  OAI22_X1  g586(.A1(new_n784), .A2(new_n785), .B1(new_n787), .B2(new_n782), .ZN(G1339gat));
  INV_X1    g587(.A(new_n583), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n790));
  AOI22_X1  g589(.A1(new_n614), .A2(KEYINPUT104), .B1(new_n618), .B2(KEYINPUT10), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n624), .B1(new_n791), .B2(new_n617), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n631), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n791), .A2(new_n624), .A3(new_n617), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n622), .A2(KEYINPUT54), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n790), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n794), .A2(new_n796), .A3(KEYINPUT117), .A4(KEYINPUT55), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(new_n632), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n799), .A2(KEYINPUT118), .A3(new_n632), .A4(new_n800), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n797), .A2(new_n798), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n803), .A2(new_n684), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n534), .A2(new_n535), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n508), .B1(new_n807), .B2(new_n532), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n539), .A2(new_n540), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n554), .B1(new_n547), .B2(new_n810), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n811), .A2(new_n633), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n668), .B1(new_n806), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n811), .A2(new_n607), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n803), .A2(new_n804), .A3(new_n805), .A4(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n789), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n684), .A2(new_n608), .A3(new_n634), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n820), .A2(new_n638), .A3(new_n501), .A4(new_n742), .ZN(new_n821));
  OAI21_X1  g620(.A(G113gat), .B1(new_n821), .B2(new_n556), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n260), .B1(new_n817), .B2(new_n819), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n823), .A2(new_n757), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n742), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n685), .A2(G113gat), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n822), .B1(new_n825), .B2(new_n826), .ZN(G1340gat));
  OAI21_X1  g626(.A(G120gat), .B1(new_n821), .B2(new_n710), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n633), .A2(G120gat), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n828), .B1(new_n825), .B2(new_n829), .ZN(G1341gat));
  NOR3_X1   g629(.A1(new_n821), .A2(new_n572), .A3(new_n789), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n824), .A2(new_n583), .A3(new_n742), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n831), .B1(new_n832), .B2(new_n572), .ZN(G1342gat));
  INV_X1    g632(.A(G134gat), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n751), .A2(new_n607), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n824), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(KEYINPUT56), .ZN(new_n837));
  INV_X1    g636(.A(new_n821), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n834), .B1(new_n838), .B2(new_n668), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n836), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT119), .B1(new_n836), .B2(KEYINPUT56), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT120), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n840), .B(new_n845), .C1(new_n841), .C2(new_n842), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(G1343gat));
  INV_X1    g646(.A(G141gat), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n820), .A2(new_n849), .A3(new_n378), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n673), .A2(new_n715), .A3(new_n260), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n555), .A2(new_n805), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n812), .B1(new_n801), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n607), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n815), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n818), .B1(new_n855), .B2(new_n789), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT57), .B1(new_n856), .B2(new_n377), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n850), .A2(new_n851), .A3(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n858), .B(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n848), .B1(new_n860), .B2(new_n684), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n673), .A2(new_n377), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n823), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n863), .A2(new_n742), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n864), .A2(new_n848), .A3(new_n555), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT58), .B1(new_n861), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(KEYINPUT58), .ZN(new_n867));
  OAI21_X1  g666(.A(G141gat), .B1(new_n858), .B2(new_n556), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n869), .ZN(G1344gat));
  INV_X1    g669(.A(G148gat), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n864), .A2(new_n871), .A3(new_n634), .ZN(new_n872));
  XNOR2_X1  g671(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n855), .A2(new_n789), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n635), .A2(new_n556), .ZN(new_n875));
  AOI211_X1 g674(.A(KEYINPUT57), .B(new_n377), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n820), .A2(new_n378), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(KEYINPUT57), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n634), .A3(new_n851), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n879), .A2(KEYINPUT123), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n871), .B1(new_n879), .B2(KEYINPUT123), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n873), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n871), .A2(KEYINPUT59), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n883), .B1(new_n860), .B2(new_n634), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n872), .B1(new_n882), .B2(new_n884), .ZN(G1345gat));
  AOI21_X1  g684(.A(G155gat), .B1(new_n864), .B2(new_n583), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n789), .A2(new_n205), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n860), .B2(new_n887), .ZN(G1346gat));
  NAND3_X1  g687(.A1(new_n863), .A2(new_n206), .A3(new_n835), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n860), .A2(new_n668), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(new_n206), .ZN(G1347gat));
  AOI21_X1  g690(.A(new_n638), .B1(new_n817), .B2(new_n819), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n742), .B1(new_n893), .B2(KEYINPUT124), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n894), .A2(new_n757), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n897), .A2(new_n264), .A3(new_n684), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n820), .A2(new_n501), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n643), .A2(new_n638), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(G169gat), .B1(new_n901), .B2(new_n556), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n898), .A2(new_n902), .ZN(G1348gat));
  NOR3_X1   g702(.A1(new_n901), .A2(new_n265), .A3(new_n710), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n897), .A2(new_n634), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(new_n265), .ZN(G1349gat));
  NAND2_X1  g705(.A1(new_n583), .A2(new_n307), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n899), .A2(new_n583), .A3(new_n900), .ZN(new_n909));
  AOI22_X1  g708(.A1(new_n897), .A2(new_n908), .B1(new_n909), .B2(new_n284), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n910), .B(new_n911), .ZN(G1350gat));
  OAI21_X1  g711(.A(G190gat), .B1(new_n901), .B2(new_n607), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT61), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n607), .A2(G190gat), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n897), .A2(KEYINPUT125), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT125), .B1(new_n897), .B2(new_n915), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(G1351gat));
  NOR3_X1   g717(.A1(new_n673), .A2(new_n638), .A3(new_n643), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n878), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(G197gat), .B1(new_n920), .B2(new_n556), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n894), .A2(new_n862), .A3(new_n896), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n684), .A2(new_n544), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(G1352gat));
  AND2_X1   g723(.A1(new_n894), .A2(new_n896), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT62), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n633), .A2(G204gat), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n925), .A2(new_n926), .A3(new_n862), .A4(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G204gat), .B1(new_n920), .B2(new_n710), .ZN(new_n929));
  INV_X1    g728(.A(new_n927), .ZN(new_n930));
  OAI21_X1  g729(.A(KEYINPUT62), .B1(new_n922), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n928), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n928), .A2(KEYINPUT126), .A3(new_n931), .A4(new_n929), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1353gat));
  INV_X1    g735(.A(new_n922), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(new_n332), .A3(new_n583), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n878), .A2(new_n583), .A3(new_n919), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n939), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT63), .B1(new_n939), .B2(G211gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(G1354gat));
  NAND3_X1  g741(.A1(new_n937), .A2(new_n333), .A3(new_n668), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n920), .A2(KEYINPUT127), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n920), .A2(KEYINPUT127), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n944), .A2(new_n945), .A3(new_n607), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n943), .B1(new_n946), .B2(new_n333), .ZN(G1355gat));
endmodule


