

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837;

  XNOR2_X1 U370 ( .A(n659), .B(KEYINPUT83), .ZN(n774) );
  AND2_X1 U371 ( .A1(n418), .A2(n417), .ZN(n413) );
  NAND2_X1 U372 ( .A1(n451), .A2(n448), .ZN(n743) );
  XNOR2_X1 U373 ( .A(n629), .B(KEYINPUT42), .ZN(n837) );
  AND2_X1 U374 ( .A1(n452), .A2(n357), .ZN(n451) );
  AND2_X1 U375 ( .A1(n459), .A2(n458), .ZN(n457) );
  NAND2_X1 U376 ( .A1(n633), .A2(n632), .ZN(n646) );
  BUF_X1 U377 ( .A(G953), .Z(n349) );
  AND2_X1 U378 ( .A1(n470), .A2(G224), .ZN(n360) );
  AND2_X1 U379 ( .A1(n551), .A2(n698), .ZN(n571) );
  XNOR2_X2 U380 ( .A(n550), .B(G469), .ZN(n698) );
  XNOR2_X2 U381 ( .A(n350), .B(n504), .ZN(n712) );
  NAND2_X1 U382 ( .A1(n411), .A2(n414), .ZN(n350) );
  NOR2_X1 U383 ( .A1(n799), .A2(n798), .ZN(n430) );
  XOR2_X1 U384 ( .A(n718), .B(n719), .Z(n351) );
  OR2_X2 U385 ( .A1(n402), .A2(n368), .ZN(n371) );
  NOR2_X2 U386 ( .A1(n815), .A2(n814), .ZN(n816) );
  AND2_X2 U387 ( .A1(n387), .A2(n386), .ZN(n385) );
  NOR2_X2 U388 ( .A1(n383), .A2(n780), .ZN(n382) );
  XNOR2_X2 U389 ( .A(n507), .B(n358), .ZN(n633) );
  XNOR2_X2 U390 ( .A(n582), .B(n543), .ZN(n824) );
  NAND2_X1 U391 ( .A1(n662), .A2(n623), .ZN(n798) );
  INV_X1 U392 ( .A(n694), .ZN(n352) );
  AND2_X1 U393 ( .A1(n647), .A2(n810), .ZN(n629) );
  INV_X1 U394 ( .A(n639), .ZN(n662) );
  XNOR2_X1 U395 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U396 ( .A(G101), .B(KEYINPUT3), .ZN(n552) );
  NAND2_X1 U397 ( .A1(n382), .A2(n370), .ZN(n384) );
  AND2_X1 U398 ( .A1(n371), .A2(n510), .ZN(n370) );
  NAND2_X1 U399 ( .A1(n712), .A2(n658), .ZN(n659) );
  OR2_X1 U400 ( .A1(n809), .A2(n808), .ZN(n353) );
  AND2_X1 U401 ( .A1(n489), .A2(n486), .ZN(n405) );
  NAND2_X1 U402 ( .A1(n416), .A2(n415), .ZN(n412) );
  AND2_X1 U403 ( .A1(n397), .A2(n398), .ZN(n396) );
  AND2_X1 U404 ( .A1(n491), .A2(n490), .ZN(n489) );
  NOR2_X1 U405 ( .A1(n395), .A2(n394), .ZN(n393) );
  AND2_X1 U406 ( .A1(n391), .A2(n390), .ZN(n397) );
  INV_X1 U407 ( .A(n400), .ZN(n399) );
  AND2_X1 U408 ( .A1(n495), .A2(n690), .ZN(n494) );
  AND2_X1 U409 ( .A1(n492), .A2(n488), .ZN(n487) );
  NAND2_X1 U410 ( .A1(n457), .A2(n454), .ZN(n657) );
  NAND2_X1 U411 ( .A1(n481), .A2(n623), .ZN(n480) );
  NAND2_X1 U412 ( .A1(n431), .A2(n632), .ZN(n799) );
  BUF_X1 U413 ( .A(n678), .Z(n783) );
  XNOR2_X1 U414 ( .A(n557), .B(n579), .ZN(n740) );
  XNOR2_X1 U415 ( .A(n557), .B(n579), .ZN(n356) );
  XNOR2_X1 U416 ( .A(n552), .B(G119), .ZN(n501) );
  INV_X1 U417 ( .A(G122), .ZN(n553) );
  XNOR2_X1 U418 ( .A(G116), .B(G113), .ZN(n500) );
  XNOR2_X1 U419 ( .A(KEYINPUT118), .B(n353), .ZN(n812) );
  NAND2_X1 U420 ( .A1(n385), .A2(n384), .ZN(n354) );
  NAND2_X1 U421 ( .A1(n385), .A2(n384), .ZN(n355) );
  NAND2_X1 U422 ( .A1(n385), .A2(n384), .ZN(n818) );
  INV_X4 U423 ( .A(G953), .ZN(n470) );
  AND2_X1 U424 ( .A1(n429), .A2(n645), .ZN(n445) );
  XNOR2_X1 U425 ( .A(n587), .B(KEYINPUT30), .ZN(n640) );
  XNOR2_X1 U426 ( .A(n527), .B(n526), .ZN(n678) );
  NAND2_X1 U427 ( .A1(n432), .A2(n435), .ZN(n400) );
  INV_X1 U428 ( .A(KEYINPUT66), .ZN(n514) );
  AND2_X1 U429 ( .A1(n506), .A2(n505), .ZN(n414) );
  XNOR2_X1 U430 ( .A(KEYINPUT15), .B(G902), .ZN(n710) );
  XOR2_X1 U431 ( .A(KEYINPUT100), .B(KEYINPUT12), .Z(n594) );
  XNOR2_X1 U432 ( .A(G140), .B(G131), .ZN(n593) );
  XOR2_X1 U433 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n592) );
  INV_X1 U434 ( .A(n688), .ZN(n496) );
  XNOR2_X1 U435 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n608) );
  XNOR2_X1 U436 ( .A(G101), .B(G146), .ZN(n546) );
  NAND2_X1 U437 ( .A1(n456), .A2(n455), .ZN(n454) );
  NOR2_X1 U438 ( .A1(n640), .A2(n460), .ZN(n455) );
  INV_X1 U439 ( .A(KEYINPUT1), .ZN(n424) );
  AND2_X1 U440 ( .A1(n475), .A2(n479), .ZN(n474) );
  INV_X1 U441 ( .A(n480), .ZN(n477) );
  NOR2_X1 U442 ( .A1(n372), .A2(n640), .ZN(n641) );
  XNOR2_X1 U443 ( .A(n675), .B(KEYINPUT22), .ZN(n676) );
  XNOR2_X1 U444 ( .A(n620), .B(n619), .ZN(n660) );
  XNOR2_X1 U445 ( .A(n605), .B(n604), .ZN(n639) );
  XNOR2_X1 U446 ( .A(n603), .B(n602), .ZN(n604) );
  NOR2_X1 U447 ( .A1(n783), .A2(n784), .ZN(n515) );
  BUF_X1 U448 ( .A(n692), .Z(n410) );
  XNOR2_X1 U449 ( .A(n482), .B(n522), .ZN(n726) );
  XNOR2_X1 U450 ( .A(n485), .B(n483), .ZN(n482) );
  XNOR2_X1 U451 ( .A(n427), .B(n426), .ZN(n521) );
  NAND2_X1 U452 ( .A1(n381), .A2(n377), .ZN(n386) );
  INV_X1 U453 ( .A(KEYINPUT46), .ZN(n419) );
  AND2_X1 U454 ( .A1(n442), .A2(n441), .ZN(n437) );
  INV_X1 U455 ( .A(n766), .ZN(n440) );
  NOR2_X1 U456 ( .A1(n837), .A2(n419), .ZN(n415) );
  NOR2_X1 U457 ( .A1(KEYINPUT73), .A2(G237), .ZN(n471) );
  NAND2_X1 U458 ( .A1(G953), .A2(KEYINPUT73), .ZN(n467) );
  NAND2_X1 U459 ( .A1(G237), .A2(G234), .ZN(n528) );
  XOR2_X1 U460 ( .A(KEYINPUT14), .B(KEYINPUT91), .Z(n529) );
  INV_X1 U461 ( .A(G237), .ZN(n568) );
  XOR2_X1 U462 ( .A(G137), .B(G140), .Z(n543) );
  NAND2_X1 U463 ( .A1(n710), .A2(n514), .ZN(n513) );
  NAND2_X1 U464 ( .A1(n711), .A2(n512), .ZN(n511) );
  NAND2_X1 U465 ( .A1(KEYINPUT2), .A2(n514), .ZN(n512) );
  NAND2_X1 U466 ( .A1(n469), .A2(n466), .ZN(n597) );
  AND2_X1 U467 ( .A1(n468), .A2(n467), .ZN(n466) );
  NAND2_X1 U468 ( .A1(n471), .A2(n470), .ZN(n469) );
  NAND2_X1 U469 ( .A1(G237), .A2(KEYINPUT73), .ZN(n468) );
  INV_X1 U470 ( .A(KEYINPUT39), .ZN(n460) );
  NAND2_X1 U471 ( .A1(n640), .A2(n460), .ZN(n458) );
  AND2_X1 U472 ( .A1(n634), .A2(n639), .ZN(n481) );
  NAND2_X1 U473 ( .A1(n497), .A2(n496), .ZN(n495) );
  INV_X1 U474 ( .A(n687), .ZN(n497) );
  NOR2_X1 U475 ( .A1(n783), .A2(n541), .ZN(n551) );
  INV_X1 U476 ( .A(G902), .ZN(n617) );
  INV_X1 U477 ( .A(G475), .ZN(n602) );
  INV_X1 U478 ( .A(KEYINPUT6), .ZN(n446) );
  XNOR2_X1 U479 ( .A(G134), .B(G131), .ZN(n542) );
  AND2_X1 U480 ( .A1(n597), .A2(G210), .ZN(n575) );
  XNOR2_X1 U481 ( .A(n428), .B(KEYINPUT24), .ZN(n427) );
  XNOR2_X1 U482 ( .A(KEYINPUT95), .B(G128), .ZN(n428) );
  XNOR2_X1 U483 ( .A(G119), .B(G110), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n543), .B(n484), .ZN(n483) );
  XNOR2_X1 U485 ( .A(KEYINPUT75), .B(KEYINPUT23), .ZN(n484) );
  NOR2_X1 U486 ( .A1(n378), .A2(n717), .ZN(n377) );
  NOR2_X1 U487 ( .A1(n380), .A2(n379), .ZN(n378) );
  INV_X1 U488 ( .A(n368), .ZN(n380) );
  INV_X1 U489 ( .A(n510), .ZN(n379) );
  XOR2_X1 U490 ( .A(KEYINPUT11), .B(G122), .Z(n589) );
  XNOR2_X1 U491 ( .A(G104), .B(G143), .ZN(n591) );
  XNOR2_X1 U492 ( .A(n430), .B(n624), .ZN(n810) );
  INV_X1 U493 ( .A(KEYINPUT35), .ZN(n488) );
  NOR2_X1 U494 ( .A1(n679), .A2(n363), .ZN(n434) );
  NOR2_X1 U495 ( .A1(n696), .A2(n447), .ZN(n790) );
  XNOR2_X1 U496 ( .A(n436), .B(n614), .ZN(n819) );
  XNOR2_X1 U497 ( .A(n613), .B(n616), .ZN(n436) );
  AND2_X1 U498 ( .A1(n654), .A2(n502), .ZN(n656) );
  NAND2_X1 U499 ( .A1(n450), .A2(n449), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n637), .B(KEYINPUT111), .ZN(n465) );
  NAND2_X1 U501 ( .A1(n636), .A2(n423), .ZN(n637) );
  NAND2_X1 U502 ( .A1(n679), .A2(n363), .ZN(n435) );
  XNOR2_X1 U503 ( .A(n408), .B(n643), .ZN(n429) );
  NOR2_X1 U504 ( .A1(n689), .A2(n502), .ZN(n642) );
  NAND2_X1 U505 ( .A1(n682), .A2(n681), .ZN(n432) );
  AND2_X1 U506 ( .A1(n362), .A2(n410), .ZN(n681) );
  NAND2_X1 U507 ( .A1(n515), .A2(n447), .ZN(n699) );
  INV_X1 U508 ( .A(n726), .ZN(n464) );
  XNOR2_X1 U509 ( .A(n432), .B(G110), .ZN(G12) );
  INV_X1 U510 ( .A(n796), .ZN(n632) );
  OR2_X1 U511 ( .A1(n453), .A2(KEYINPUT40), .ZN(n357) );
  XOR2_X1 U512 ( .A(n570), .B(n569), .Z(n358) );
  XOR2_X1 U513 ( .A(KEYINPUT71), .B(KEYINPUT38), .Z(n359) );
  AND2_X1 U514 ( .A1(n434), .A2(KEYINPUT85), .ZN(n361) );
  INV_X1 U515 ( .A(n622), .ZN(n431) );
  AND2_X1 U516 ( .A1(n678), .A2(n625), .ZN(n630) );
  AND2_X1 U517 ( .A1(n783), .A2(n447), .ZN(n362) );
  INV_X1 U518 ( .A(n769), .ZN(n453) );
  XNOR2_X1 U519 ( .A(KEYINPUT79), .B(KEYINPUT32), .ZN(n363) );
  AND2_X1 U520 ( .A1(n648), .A2(KEYINPUT70), .ZN(n364) );
  AND2_X1 U521 ( .A1(n363), .A2(KEYINPUT85), .ZN(n365) );
  AND2_X1 U522 ( .A1(n496), .A2(KEYINPUT35), .ZN(n366) );
  XOR2_X1 U523 ( .A(n723), .B(n722), .Z(n367) );
  NAND2_X1 U524 ( .A1(n777), .A2(KEYINPUT66), .ZN(n368) );
  AND2_X1 U525 ( .A1(n711), .A2(n514), .ZN(n369) );
  XNOR2_X1 U526 ( .A(n405), .B(G122), .ZN(G24) );
  NAND2_X1 U527 ( .A1(n405), .A2(n406), .ZN(n404) );
  NAND2_X1 U528 ( .A1(n393), .A2(n399), .ZN(n392) );
  NAND2_X1 U529 ( .A1(n513), .A2(n511), .ZN(n510) );
  NAND2_X1 U530 ( .A1(n698), .A2(n551), .ZN(n372) );
  XNOR2_X2 U531 ( .A(n373), .B(n583), .ZN(n788) );
  NOR2_X1 U532 ( .A1(n723), .A2(G902), .ZN(n373) );
  NAND2_X1 U533 ( .A1(n403), .A2(n706), .ZN(n708) );
  XNOR2_X1 U534 ( .A(n404), .B(n691), .ZN(n403) );
  INV_X1 U535 ( .A(n657), .ZN(n450) );
  NOR2_X2 U536 ( .A1(n692), .A2(n421), .ZN(n695) );
  AND2_X2 U537 ( .A1(n709), .A2(n731), .ZN(n402) );
  XNOR2_X1 U538 ( .A(n508), .B(n356), .ZN(n374) );
  XNOR2_X1 U539 ( .A(n508), .B(n740), .ZN(n752) );
  AND2_X1 U540 ( .A1(n498), .A2(n494), .ZN(n375) );
  INV_X1 U541 ( .A(n804), .ZN(n376) );
  XNOR2_X1 U542 ( .A(n685), .B(KEYINPUT33), .ZN(n420) );
  NAND2_X1 U543 ( .A1(n402), .A2(n510), .ZN(n381) );
  INV_X1 U544 ( .A(n389), .ZN(n780) );
  NAND2_X1 U545 ( .A1(n389), .A2(n407), .ZN(n388) );
  XNOR2_X2 U546 ( .A(n716), .B(KEYINPUT74), .ZN(n389) );
  NAND2_X1 U547 ( .A1(n407), .A2(n717), .ZN(n383) );
  NAND2_X1 U548 ( .A1(n388), .A2(KEYINPUT65), .ZN(n387) );
  NAND2_X1 U549 ( .A1(n694), .A2(n363), .ZN(n401) );
  NAND2_X1 U550 ( .A1(n352), .A2(n434), .ZN(n425) );
  NAND2_X1 U551 ( .A1(n694), .A2(n365), .ZN(n390) );
  NAND2_X1 U552 ( .A1(n352), .A2(n361), .ZN(n391) );
  NAND2_X1 U553 ( .A1(n396), .A2(n392), .ZN(n406) );
  NAND2_X1 U554 ( .A1(n401), .A2(n683), .ZN(n394) );
  INV_X1 U555 ( .A(n425), .ZN(n395) );
  NAND2_X1 U556 ( .A1(n400), .A2(KEYINPUT85), .ZN(n398) );
  AND2_X1 U557 ( .A1(n401), .A2(n435), .ZN(n433) );
  NAND2_X1 U558 ( .A1(n402), .A2(n369), .ZN(n407) );
  NAND2_X1 U559 ( .A1(n837), .A2(n419), .ZN(n417) );
  NAND2_X1 U560 ( .A1(n612), .A2(G221), .ZN(n485) );
  XNOR2_X2 U561 ( .A(n708), .B(n707), .ZN(n731) );
  NAND2_X1 U562 ( .A1(n641), .A2(n642), .ZN(n408) );
  NAND2_X1 U563 ( .A1(n375), .A2(n487), .ZN(n486) );
  OR2_X1 U564 ( .A1(n420), .A2(n688), .ZN(n492) );
  NAND2_X1 U565 ( .A1(n413), .A2(n412), .ZN(n411) );
  INV_X1 U566 ( .A(n743), .ZN(n416) );
  NAND2_X1 U567 ( .A1(n743), .A2(n419), .ZN(n418) );
  INV_X1 U568 ( .A(n420), .ZN(n804) );
  NAND2_X1 U569 ( .A1(n499), .A2(n420), .ZN(n498) );
  NAND2_X1 U570 ( .A1(n376), .A2(n810), .ZN(n811) );
  AND2_X1 U571 ( .A1(n421), .A2(n692), .ZN(n782) );
  INV_X1 U572 ( .A(n515), .ZN(n421) );
  OR2_X1 U573 ( .A1(n692), .A2(n422), .ZN(n679) );
  INV_X1 U574 ( .A(n783), .ZN(n422) );
  INV_X1 U575 ( .A(n692), .ZN(n423) );
  XNOR2_X2 U576 ( .A(n698), .B(n424), .ZN(n692) );
  NAND2_X1 U577 ( .A1(n433), .A2(n425), .ZN(n744) );
  XNOR2_X1 U578 ( .A(n429), .B(G143), .ZN(G45) );
  NAND2_X1 U579 ( .A1(n657), .A2(n621), .ZN(n452) );
  NAND2_X1 U580 ( .A1(n438), .A2(n437), .ZN(n444) );
  NAND2_X1 U581 ( .A1(n439), .A2(n440), .ZN(n438) );
  NOR2_X1 U582 ( .A1(n800), .A2(n364), .ZN(n439) );
  NAND2_X1 U583 ( .A1(n800), .A2(n364), .ZN(n441) );
  NAND2_X1 U584 ( .A1(n766), .A2(n364), .ZN(n442) );
  XNOR2_X1 U585 ( .A(n443), .B(KEYINPUT69), .ZN(n506) );
  NAND2_X1 U586 ( .A1(n445), .A2(n444), .ZN(n443) );
  NAND2_X1 U587 ( .A1(n788), .A2(n632), .ZN(n587) );
  XNOR2_X1 U588 ( .A(n788), .B(n446), .ZN(n684) );
  INV_X1 U589 ( .A(n788), .ZN(n447) );
  NAND2_X2 U590 ( .A1(n671), .A2(n670), .ZN(n509) );
  XNOR2_X2 U591 ( .A(n646), .B(KEYINPUT19), .ZN(n671) );
  NOR2_X1 U592 ( .A1(n769), .A2(n621), .ZN(n449) );
  INV_X1 U593 ( .A(n588), .ZN(n456) );
  NAND2_X1 U594 ( .A1(n588), .A2(n460), .ZN(n459) );
  XNOR2_X1 U595 ( .A(n461), .B(n367), .ZN(n517) );
  NAND2_X1 U596 ( .A1(n354), .A2(G472), .ZN(n461) );
  XNOR2_X1 U597 ( .A(n462), .B(n351), .ZN(n518) );
  NAND2_X1 U598 ( .A1(n355), .A2(G469), .ZN(n462) );
  NAND2_X1 U599 ( .A1(n463), .A2(n724), .ZN(n728) );
  XNOR2_X1 U600 ( .A(n727), .B(n464), .ZN(n463) );
  XNOR2_X1 U601 ( .A(n465), .B(n638), .ZN(n505) );
  XNOR2_X1 U602 ( .A(n465), .B(G125), .ZN(n835) );
  NAND2_X1 U603 ( .A1(n474), .A2(n472), .ZN(n636) );
  NAND2_X1 U604 ( .A1(n473), .A2(n477), .ZN(n472) );
  AND2_X1 U605 ( .A1(n476), .A2(n684), .ZN(n473) );
  NAND2_X1 U606 ( .A1(n478), .A2(n635), .ZN(n475) );
  NAND2_X1 U607 ( .A1(n630), .A2(n684), .ZN(n478) );
  NOR2_X1 U608 ( .A1(n631), .A2(n635), .ZN(n476) );
  NAND2_X1 U609 ( .A1(n480), .A2(n635), .ZN(n479) );
  NOR2_X1 U610 ( .A1(n631), .A2(n769), .ZN(n649) );
  NAND2_X1 U611 ( .A1(n623), .A2(n639), .ZN(n769) );
  NAND2_X1 U612 ( .A1(n804), .A2(n366), .ZN(n490) );
  NAND2_X1 U613 ( .A1(n493), .A2(KEYINPUT35), .ZN(n491) );
  NAND2_X1 U614 ( .A1(n498), .A2(n494), .ZN(n493) );
  AND2_X1 U615 ( .A1(n687), .A2(n688), .ZN(n499) );
  XNOR2_X2 U616 ( .A(n501), .B(n500), .ZN(n579) );
  XNOR2_X1 U617 ( .A(n633), .B(n359), .ZN(n622) );
  INV_X1 U618 ( .A(n633), .ZN(n502) );
  XNOR2_X2 U619 ( .A(n503), .B(G143), .ZN(n615) );
  XNOR2_X2 U620 ( .A(G128), .B(KEYINPUT80), .ZN(n503) );
  INV_X1 U621 ( .A(KEYINPUT48), .ZN(n504) );
  NAND2_X1 U622 ( .A1(n752), .A2(n710), .ZN(n507) );
  NAND2_X1 U623 ( .A1(n566), .A2(n567), .ZN(n508) );
  NAND2_X1 U624 ( .A1(n686), .A2(n674), .ZN(n677) );
  XNOR2_X2 U625 ( .A(n509), .B(n673), .ZN(n686) );
  XNOR2_X1 U626 ( .A(n360), .B(n520), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n520), .B(KEYINPUT10), .ZN(n825) );
  NOR2_X2 U628 ( .A1(n749), .A2(n823), .ZN(n750) );
  NOR2_X2 U629 ( .A1(n755), .A2(n823), .ZN(n757) );
  XNOR2_X1 U630 ( .A(n560), .B(n561), .ZN(n562) );
  XNOR2_X2 U631 ( .A(n563), .B(n542), .ZN(n582) );
  XNOR2_X2 U632 ( .A(n544), .B(G104), .ZN(n556) );
  XNOR2_X2 U633 ( .A(G110), .B(G107), .ZN(n544) );
  NAND2_X1 U634 ( .A1(n712), .A2(n836), .ZN(n516) );
  XNOR2_X1 U635 ( .A(n589), .B(G113), .ZN(n590) );
  BUF_X1 U636 ( .A(n731), .Z(n776) );
  INV_X1 U637 ( .A(n823), .ZN(n724) );
  NAND2_X1 U638 ( .A1(G234), .A2(n470), .ZN(n519) );
  XOR2_X1 U639 ( .A(KEYINPUT8), .B(n519), .Z(n612) );
  XNOR2_X2 U640 ( .A(G125), .B(G146), .ZN(n520) );
  XNOR2_X1 U641 ( .A(n825), .B(n521), .ZN(n522) );
  NAND2_X1 U642 ( .A1(n726), .A2(n617), .ZN(n527) );
  NAND2_X1 U643 ( .A1(G234), .A2(n710), .ZN(n523) );
  XNOR2_X1 U644 ( .A(KEYINPUT20), .B(n523), .ZN(n536) );
  NAND2_X1 U645 ( .A1(n536), .A2(G217), .ZN(n524) );
  XNOR2_X1 U646 ( .A(n524), .B(KEYINPUT25), .ZN(n525) );
  XNOR2_X1 U647 ( .A(n525), .B(KEYINPUT96), .ZN(n526) );
  XNOR2_X1 U648 ( .A(n529), .B(n528), .ZN(n531) );
  NAND2_X1 U649 ( .A1(G952), .A2(n531), .ZN(n809) );
  NOR2_X1 U650 ( .A1(n349), .A2(n809), .ZN(n530) );
  XNOR2_X1 U651 ( .A(n530), .B(KEYINPUT92), .ZN(n669) );
  NAND2_X1 U652 ( .A1(G902), .A2(n531), .ZN(n665) );
  NOR2_X1 U653 ( .A1(G900), .A2(n665), .ZN(n532) );
  AND2_X1 U654 ( .A1(n349), .A2(n532), .ZN(n533) );
  OR2_X1 U655 ( .A1(n669), .A2(n533), .ZN(n535) );
  INV_X1 U656 ( .A(KEYINPUT81), .ZN(n534) );
  XNOR2_X1 U657 ( .A(n535), .B(n534), .ZN(n540) );
  NAND2_X1 U658 ( .A1(n536), .A2(G221), .ZN(n538) );
  XOR2_X1 U659 ( .A(KEYINPUT21), .B(KEYINPUT97), .Z(n537) );
  XNOR2_X1 U660 ( .A(n538), .B(n537), .ZN(n784) );
  INV_X1 U661 ( .A(n784), .ZN(n539) );
  AND2_X1 U662 ( .A1(n540), .A2(n539), .ZN(n625) );
  INV_X1 U663 ( .A(n625), .ZN(n541) );
  XNOR2_X2 U664 ( .A(n615), .B(KEYINPUT4), .ZN(n563) );
  NAND2_X1 U665 ( .A1(G227), .A2(n470), .ZN(n545) );
  XNOR2_X1 U666 ( .A(n545), .B(KEYINPUT94), .ZN(n547) );
  XNOR2_X1 U667 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U668 ( .A(n556), .B(n548), .ZN(n549) );
  XNOR2_X1 U669 ( .A(n824), .B(n549), .ZN(n718) );
  OR2_X2 U670 ( .A1(n718), .A2(G902), .ZN(n550) );
  XNOR2_X1 U671 ( .A(KEYINPUT68), .B(KEYINPUT16), .ZN(n554) );
  XNOR2_X1 U672 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U673 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n559) );
  XNOR2_X1 U674 ( .A(KEYINPUT88), .B(KEYINPUT76), .ZN(n558) );
  XNOR2_X1 U675 ( .A(n559), .B(n558), .ZN(n561) );
  NAND2_X1 U676 ( .A1(n562), .A2(n563), .ZN(n567) );
  INV_X1 U677 ( .A(n562), .ZN(n565) );
  INV_X1 U678 ( .A(n563), .ZN(n564) );
  NAND2_X1 U679 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U680 ( .A1(n617), .A2(n568), .ZN(n584) );
  NAND2_X1 U681 ( .A1(n584), .A2(G210), .ZN(n570) );
  INV_X1 U682 ( .A(KEYINPUT89), .ZN(n569) );
  NAND2_X1 U683 ( .A1(n571), .A2(n431), .ZN(n588) );
  XNOR2_X1 U684 ( .A(KEYINPUT5), .B(G137), .ZN(n572) );
  XNOR2_X1 U685 ( .A(n572), .B(G146), .ZN(n574) );
  NAND2_X1 U686 ( .A1(n597), .A2(G210), .ZN(n573) );
  NAND2_X1 U687 ( .A1(n574), .A2(n573), .ZN(n578) );
  INV_X1 U688 ( .A(n574), .ZN(n576) );
  NAND2_X1 U689 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U690 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U691 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U692 ( .A(n582), .B(n581), .ZN(n723) );
  INV_X1 U693 ( .A(G472), .ZN(n583) );
  NAND2_X1 U694 ( .A1(n584), .A2(G214), .ZN(n586) );
  INV_X1 U695 ( .A(KEYINPUT90), .ZN(n585) );
  XNOR2_X1 U696 ( .A(n586), .B(n585), .ZN(n796) );
  XNOR2_X1 U697 ( .A(n825), .B(n590), .ZN(n601) );
  XNOR2_X1 U698 ( .A(n592), .B(n591), .ZN(n596) );
  XNOR2_X1 U699 ( .A(n594), .B(n593), .ZN(n595) );
  XOR2_X1 U700 ( .A(n596), .B(n595), .Z(n599) );
  NAND2_X1 U701 ( .A1(n597), .A2(G214), .ZN(n598) );
  XNOR2_X1 U702 ( .A(n599), .B(n598), .ZN(n600) );
  XNOR2_X1 U703 ( .A(n601), .B(n600), .ZN(n745) );
  NOR2_X1 U704 ( .A1(G902), .A2(n745), .ZN(n605) );
  INV_X1 U705 ( .A(KEYINPUT13), .ZN(n603) );
  XOR2_X1 U706 ( .A(G134), .B(G122), .Z(n607) );
  XNOR2_X1 U707 ( .A(G116), .B(G107), .ZN(n606) );
  XNOR2_X1 U708 ( .A(n607), .B(n606), .ZN(n611) );
  XOR2_X1 U709 ( .A(KEYINPUT102), .B(KEYINPUT101), .Z(n609) );
  XNOR2_X1 U710 ( .A(n609), .B(n608), .ZN(n610) );
  XOR2_X1 U711 ( .A(n611), .B(n610), .Z(n614) );
  NAND2_X1 U712 ( .A1(G217), .A2(n612), .ZN(n613) );
  INV_X1 U713 ( .A(n615), .ZN(n616) );
  NAND2_X1 U714 ( .A1(n819), .A2(n617), .ZN(n620) );
  INV_X1 U715 ( .A(KEYINPUT103), .ZN(n618) );
  XNOR2_X1 U716 ( .A(n618), .B(G478), .ZN(n619) );
  INV_X1 U717 ( .A(n660), .ZN(n623) );
  INV_X1 U718 ( .A(KEYINPUT40), .ZN(n621) );
  XNOR2_X1 U719 ( .A(KEYINPUT41), .B(KEYINPUT109), .ZN(n624) );
  NAND2_X1 U720 ( .A1(n630), .A2(n788), .ZN(n627) );
  XOR2_X1 U721 ( .A(KEYINPUT28), .B(KEYINPUT108), .Z(n626) );
  XNOR2_X1 U722 ( .A(n627), .B(n626), .ZN(n628) );
  AND2_X1 U723 ( .A1(n698), .A2(n628), .ZN(n647) );
  INV_X1 U724 ( .A(n630), .ZN(n631) );
  INV_X1 U725 ( .A(n646), .ZN(n634) );
  XOR2_X1 U726 ( .A(KEYINPUT36), .B(KEYINPUT110), .Z(n635) );
  INV_X1 U727 ( .A(KEYINPUT84), .ZN(n638) );
  NAND2_X1 U728 ( .A1(n639), .A2(n660), .ZN(n689) );
  INV_X1 U729 ( .A(KEYINPUT107), .ZN(n643) );
  INV_X1 U730 ( .A(KEYINPUT70), .ZN(n644) );
  NAND2_X1 U731 ( .A1(n644), .A2(KEYINPUT47), .ZN(n645) );
  NAND2_X1 U732 ( .A1(n647), .A2(n671), .ZN(n766) );
  NAND2_X1 U733 ( .A1(n662), .A2(n660), .ZN(n772) );
  AND2_X1 U734 ( .A1(n772), .A2(n769), .ZN(n800) );
  INV_X1 U735 ( .A(KEYINPUT47), .ZN(n648) );
  AND2_X1 U736 ( .A1(n649), .A2(n684), .ZN(n650) );
  NAND2_X1 U737 ( .A1(n692), .A2(n650), .ZN(n651) );
  NOR2_X1 U738 ( .A1(n796), .A2(n651), .ZN(n653) );
  XNOR2_X1 U739 ( .A(KEYINPUT43), .B(KEYINPUT105), .ZN(n652) );
  XNOR2_X1 U740 ( .A(n653), .B(n652), .ZN(n654) );
  INV_X1 U741 ( .A(KEYINPUT106), .ZN(n655) );
  XNOR2_X1 U742 ( .A(n656), .B(n655), .ZN(n836) );
  OR2_X1 U743 ( .A1(n657), .A2(n772), .ZN(n730) );
  AND2_X1 U744 ( .A1(n836), .A2(n730), .ZN(n658) );
  XNOR2_X1 U745 ( .A(n774), .B(KEYINPUT72), .ZN(n709) );
  NOR2_X1 U746 ( .A1(n660), .A2(n784), .ZN(n661) );
  NAND2_X1 U747 ( .A1(n662), .A2(n661), .ZN(n664) );
  INV_X1 U748 ( .A(KEYINPUT104), .ZN(n663) );
  XNOR2_X1 U749 ( .A(n664), .B(n663), .ZN(n674) );
  INV_X1 U750 ( .A(n665), .ZN(n666) );
  NOR2_X1 U751 ( .A1(G898), .A2(n470), .ZN(n738) );
  NAND2_X1 U752 ( .A1(n666), .A2(n738), .ZN(n667) );
  XNOR2_X1 U753 ( .A(n667), .B(KEYINPUT93), .ZN(n668) );
  OR2_X1 U754 ( .A1(n669), .A2(n668), .ZN(n670) );
  INV_X1 U755 ( .A(KEYINPUT86), .ZN(n672) );
  XNOR2_X1 U756 ( .A(n672), .B(KEYINPUT0), .ZN(n673) );
  INV_X1 U757 ( .A(KEYINPUT67), .ZN(n675) );
  XNOR2_X1 U758 ( .A(n677), .B(n676), .ZN(n680) );
  OR2_X2 U759 ( .A1(n680), .A2(n684), .ZN(n694) );
  INV_X1 U760 ( .A(n680), .ZN(n682) );
  INV_X1 U761 ( .A(KEYINPUT85), .ZN(n683) );
  NAND2_X1 U762 ( .A1(n695), .A2(n684), .ZN(n685) );
  BUF_X1 U763 ( .A(n686), .Z(n687) );
  XOR2_X1 U764 ( .A(KEYINPUT34), .B(KEYINPUT78), .Z(n688) );
  XNOR2_X1 U765 ( .A(n689), .B(KEYINPUT77), .ZN(n690) );
  INV_X1 U766 ( .A(KEYINPUT44), .ZN(n691) );
  NAND2_X1 U767 ( .A1(n410), .A2(n422), .ZN(n693) );
  NOR2_X1 U768 ( .A1(n694), .A2(n693), .ZN(n758) );
  INV_X1 U769 ( .A(n758), .ZN(n705) );
  INV_X1 U770 ( .A(n695), .ZN(n696) );
  NAND2_X1 U771 ( .A1(n790), .A2(n687), .ZN(n697) );
  XOR2_X1 U772 ( .A(KEYINPUT31), .B(n697), .Z(n771) );
  INV_X1 U773 ( .A(n698), .ZN(n700) );
  NOR2_X1 U774 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U775 ( .A1(n687), .A2(n701), .ZN(n760) );
  NAND2_X1 U776 ( .A1(n771), .A2(n760), .ZN(n703) );
  INV_X1 U777 ( .A(n800), .ZN(n702) );
  NAND2_X1 U778 ( .A1(n703), .A2(n702), .ZN(n704) );
  AND2_X1 U779 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U780 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n707) );
  INV_X1 U781 ( .A(KEYINPUT2), .ZN(n777) );
  INV_X1 U782 ( .A(n710), .ZN(n711) );
  NAND2_X1 U783 ( .A1(n730), .A2(KEYINPUT2), .ZN(n713) );
  XNOR2_X1 U784 ( .A(n713), .B(KEYINPUT82), .ZN(n714) );
  NOR2_X1 U785 ( .A1(n516), .A2(n714), .ZN(n715) );
  NAND2_X1 U786 ( .A1(n731), .A2(n715), .ZN(n716) );
  INV_X1 U787 ( .A(KEYINPUT65), .ZN(n717) );
  XOR2_X1 U788 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n719) );
  INV_X1 U789 ( .A(G952), .ZN(n720) );
  AND2_X1 U790 ( .A1(n720), .A2(n349), .ZN(n823) );
  NAND2_X1 U791 ( .A1(n518), .A2(n724), .ZN(n721) );
  XNOR2_X1 U792 ( .A(n721), .B(KEYINPUT121), .ZN(G54) );
  XNOR2_X1 U793 ( .A(KEYINPUT112), .B(KEYINPUT62), .ZN(n722) );
  NAND2_X1 U794 ( .A1(n517), .A2(n724), .ZN(n725) );
  XNOR2_X1 U795 ( .A(n725), .B(KEYINPUT63), .ZN(G57) );
  AND2_X2 U796 ( .A1(n355), .A2(G217), .ZN(n727) );
  XNOR2_X1 U797 ( .A(n728), .B(KEYINPUT123), .ZN(G66) );
  XNOR2_X1 U798 ( .A(G134), .B(KEYINPUT114), .ZN(n729) );
  XNOR2_X1 U799 ( .A(n730), .B(n729), .ZN(G36) );
  INV_X1 U800 ( .A(n776), .ZN(n732) );
  NOR2_X1 U801 ( .A1(n732), .A2(n349), .ZN(n737) );
  NAND2_X1 U802 ( .A1(n349), .A2(G224), .ZN(n733) );
  XNOR2_X1 U803 ( .A(KEYINPUT61), .B(n733), .ZN(n734) );
  NAND2_X1 U804 ( .A1(n734), .A2(G898), .ZN(n735) );
  XOR2_X1 U805 ( .A(KEYINPUT124), .B(n735), .Z(n736) );
  NOR2_X1 U806 ( .A1(n737), .A2(n736), .ZN(n742) );
  INV_X1 U807 ( .A(n738), .ZN(n739) );
  NAND2_X1 U808 ( .A1(n356), .A2(n739), .ZN(n741) );
  XNOR2_X1 U809 ( .A(n742), .B(n741), .ZN(G69) );
  XOR2_X1 U810 ( .A(n743), .B(G131), .Z(G33) );
  XOR2_X1 U811 ( .A(G119), .B(n744), .Z(G21) );
  NAND2_X1 U812 ( .A1(n818), .A2(G475), .ZN(n748) );
  XNOR2_X1 U813 ( .A(KEYINPUT87), .B(KEYINPUT59), .ZN(n746) );
  XNOR2_X1 U814 ( .A(n745), .B(n746), .ZN(n747) );
  XNOR2_X1 U815 ( .A(n748), .B(n747), .ZN(n749) );
  XNOR2_X1 U816 ( .A(n750), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U817 ( .A1(n818), .A2(G210), .ZN(n754) );
  XNOR2_X1 U818 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n751) );
  XNOR2_X1 U819 ( .A(n374), .B(n751), .ZN(n753) );
  XNOR2_X1 U820 ( .A(n754), .B(n753), .ZN(n755) );
  XNOR2_X1 U821 ( .A(KEYINPUT120), .B(KEYINPUT56), .ZN(n756) );
  XNOR2_X1 U822 ( .A(n757), .B(n756), .ZN(G51) );
  XOR2_X1 U823 ( .A(G101), .B(n758), .Z(G3) );
  NOR2_X1 U824 ( .A1(n769), .A2(n760), .ZN(n759) );
  XOR2_X1 U825 ( .A(G104), .B(n759), .Z(G6) );
  NOR2_X1 U826 ( .A1(n772), .A2(n760), .ZN(n762) );
  XNOR2_X1 U827 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n761) );
  XNOR2_X1 U828 ( .A(n762), .B(n761), .ZN(n763) );
  XNOR2_X1 U829 ( .A(G107), .B(n763), .ZN(G9) );
  XOR2_X1 U830 ( .A(G128), .B(KEYINPUT29), .Z(n765) );
  OR2_X1 U831 ( .A1(n772), .A2(n766), .ZN(n764) );
  XNOR2_X1 U832 ( .A(n765), .B(n764), .ZN(G30) );
  XOR2_X1 U833 ( .A(G146), .B(KEYINPUT113), .Z(n768) );
  OR2_X1 U834 ( .A1(n769), .A2(n766), .ZN(n767) );
  XNOR2_X1 U835 ( .A(n768), .B(n767), .ZN(G48) );
  NOR2_X1 U836 ( .A1(n769), .A2(n771), .ZN(n770) );
  XOR2_X1 U837 ( .A(G113), .B(n770), .Z(G15) );
  NOR2_X1 U838 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U839 ( .A(G116), .B(n773), .Z(G18) );
  BUF_X1 U840 ( .A(n774), .Z(n775) );
  NAND2_X1 U841 ( .A1(n775), .A2(n776), .ZN(n778) );
  AND2_X1 U842 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U843 ( .A1(n780), .A2(n779), .ZN(n815) );
  XNOR2_X1 U844 ( .A(KEYINPUT115), .B(KEYINPUT50), .ZN(n781) );
  XNOR2_X1 U845 ( .A(n782), .B(n781), .ZN(n787) );
  NAND2_X1 U846 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U847 ( .A(KEYINPUT49), .B(n785), .Z(n786) );
  NAND2_X1 U848 ( .A1(n787), .A2(n786), .ZN(n789) );
  NOR2_X1 U849 ( .A1(n789), .A2(n788), .ZN(n791) );
  NOR2_X1 U850 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U851 ( .A(n792), .B(KEYINPUT116), .ZN(n793) );
  XNOR2_X1 U852 ( .A(n793), .B(KEYINPUT51), .ZN(n794) );
  NAND2_X1 U853 ( .A1(n794), .A2(n810), .ZN(n795) );
  XNOR2_X1 U854 ( .A(n795), .B(KEYINPUT117), .ZN(n806) );
  AND2_X1 U855 ( .A1(n622), .A2(n796), .ZN(n797) );
  NOR2_X1 U856 ( .A1(n798), .A2(n797), .ZN(n802) );
  NOR2_X1 U857 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U858 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U859 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U860 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U861 ( .A(n807), .B(KEYINPUT52), .ZN(n808) );
  NAND2_X1 U862 ( .A1(n812), .A2(n811), .ZN(n813) );
  XOR2_X1 U863 ( .A(KEYINPUT119), .B(n813), .Z(n814) );
  NAND2_X1 U864 ( .A1(n470), .A2(n816), .ZN(n817) );
  XOR2_X1 U865 ( .A(KEYINPUT53), .B(n817), .Z(G75) );
  NAND2_X1 U866 ( .A1(n354), .A2(G478), .ZN(n821) );
  XOR2_X1 U867 ( .A(KEYINPUT122), .B(n819), .Z(n820) );
  XNOR2_X1 U868 ( .A(n821), .B(n820), .ZN(n822) );
  NOR2_X1 U869 ( .A1(n823), .A2(n822), .ZN(G63) );
  XNOR2_X1 U870 ( .A(n824), .B(n825), .ZN(n828) );
  XNOR2_X1 U871 ( .A(n828), .B(KEYINPUT125), .ZN(n826) );
  XNOR2_X1 U872 ( .A(n775), .B(n826), .ZN(n827) );
  NAND2_X1 U873 ( .A1(n827), .A2(n470), .ZN(n834) );
  XNOR2_X1 U874 ( .A(G227), .B(KEYINPUT126), .ZN(n829) );
  XNOR2_X1 U875 ( .A(n829), .B(n828), .ZN(n830) );
  NAND2_X1 U876 ( .A1(G900), .A2(n830), .ZN(n831) );
  XOR2_X1 U877 ( .A(KEYINPUT127), .B(n831), .Z(n832) );
  NAND2_X1 U878 ( .A1(n349), .A2(n832), .ZN(n833) );
  NAND2_X1 U879 ( .A1(n834), .A2(n833), .ZN(G72) );
  XNOR2_X1 U880 ( .A(n835), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U881 ( .A(G140), .B(n836), .ZN(G42) );
  XOR2_X1 U882 ( .A(n837), .B(G137), .Z(G39) );
endmodule

