

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U553 ( .A(n742), .B(n741), .ZN(n764) );
  BUF_X1 U554 ( .A(n720), .Z(n732) );
  INV_X1 U555 ( .A(n732), .ZN(n714) );
  NOR2_X1 U556 ( .A1(G164), .A2(G1384), .ZN(n777) );
  NOR2_X2 U557 ( .A1(G2104), .A2(G2105), .ZN(n525) );
  NAND2_X1 U558 ( .A1(n683), .A2(n777), .ZN(n720) );
  AND2_X2 U559 ( .A1(n740), .A2(n739), .ZN(n742) );
  XOR2_X2 U560 ( .A(KEYINPUT66), .B(n526), .Z(n611) );
  NOR2_X1 U561 ( .A1(n720), .A2(n989), .ZN(n685) );
  NOR2_X1 U562 ( .A1(n709), .A2(G299), .ZN(n688) );
  INV_X1 U563 ( .A(G2105), .ZN(n522) );
  NOR2_X1 U564 ( .A1(n648), .A2(G651), .ZN(n653) );
  NOR2_X2 U565 ( .A1(n531), .A2(n530), .ZN(G160) );
  INV_X1 U566 ( .A(KEYINPUT31), .ZN(n727) );
  XNOR2_X1 U567 ( .A(n727), .B(KEYINPUT97), .ZN(n728) );
  XNOR2_X1 U568 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U569 ( .A(KEYINPUT100), .B(KEYINPUT32), .ZN(n741) );
  INV_X1 U570 ( .A(KEYINPUT103), .ZN(n761) );
  NAND2_X1 U571 ( .A1(G8), .A2(n720), .ZN(n775) );
  INV_X1 U572 ( .A(G651), .ZN(n535) );
  XNOR2_X1 U573 ( .A(KEYINPUT68), .B(n537), .ZN(n652) );
  NOR2_X1 U574 ( .A1(n829), .A2(n828), .ZN(n830) );
  AND2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n894) );
  NAND2_X1 U576 ( .A1(G113), .A2(n894), .ZN(n521) );
  NOR2_X2 U577 ( .A1(G2104), .A2(n522), .ZN(n895) );
  NAND2_X1 U578 ( .A1(G125), .A2(n895), .ZN(n520) );
  NAND2_X1 U579 ( .A1(n521), .A2(n520), .ZN(n531) );
  NAND2_X1 U580 ( .A1(n522), .A2(G2104), .ZN(n523) );
  XNOR2_X2 U581 ( .A(n523), .B(KEYINPUT65), .ZN(n898) );
  NAND2_X1 U582 ( .A1(G101), .A2(n898), .ZN(n524) );
  XOR2_X1 U583 ( .A(KEYINPUT23), .B(n524), .Z(n529) );
  XNOR2_X1 U584 ( .A(n525), .B(KEYINPUT17), .ZN(n526) );
  NAND2_X1 U585 ( .A1(G137), .A2(n611), .ZN(n527) );
  XOR2_X1 U586 ( .A(n527), .B(KEYINPUT67), .Z(n528) );
  NAND2_X1 U587 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U588 ( .A(KEYINPUT0), .B(G543), .Z(n648) );
  NOR2_X1 U589 ( .A1(n648), .A2(n535), .ZN(n639) );
  NAND2_X1 U590 ( .A1(G78), .A2(n639), .ZN(n534) );
  NOR2_X1 U591 ( .A1(G651), .A2(G543), .ZN(n532) );
  XNOR2_X1 U592 ( .A(n532), .B(KEYINPUT64), .ZN(n640) );
  NAND2_X1 U593 ( .A1(G91), .A2(n640), .ZN(n533) );
  NAND2_X1 U594 ( .A1(n534), .A2(n533), .ZN(n541) );
  NAND2_X1 U595 ( .A1(n653), .A2(G53), .ZN(n539) );
  NOR2_X1 U596 ( .A1(G543), .A2(n535), .ZN(n536) );
  XOR2_X1 U597 ( .A(KEYINPUT1), .B(n536), .Z(n537) );
  NAND2_X1 U598 ( .A1(G65), .A2(n652), .ZN(n538) );
  NAND2_X1 U599 ( .A1(n539), .A2(n538), .ZN(n540) );
  OR2_X1 U600 ( .A1(n541), .A2(n540), .ZN(G299) );
  NAND2_X1 U601 ( .A1(G126), .A2(n895), .ZN(n543) );
  NAND2_X1 U602 ( .A1(n611), .A2(G138), .ZN(n542) );
  NAND2_X1 U603 ( .A1(n543), .A2(n542), .ZN(n547) );
  NAND2_X1 U604 ( .A1(G114), .A2(n894), .ZN(n545) );
  NAND2_X1 U605 ( .A1(G102), .A2(n898), .ZN(n544) );
  NAND2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U607 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U608 ( .A(KEYINPUT87), .B(n548), .Z(G164) );
  NAND2_X1 U609 ( .A1(G72), .A2(n639), .ZN(n550) );
  NAND2_X1 U610 ( .A1(G85), .A2(n640), .ZN(n549) );
  NAND2_X1 U611 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n653), .A2(G47), .ZN(n552) );
  NAND2_X1 U613 ( .A1(G60), .A2(n652), .ZN(n551) );
  NAND2_X1 U614 ( .A1(n552), .A2(n551), .ZN(n553) );
  OR2_X1 U615 ( .A1(n554), .A2(n553), .ZN(G290) );
  INV_X1 U616 ( .A(G132), .ZN(G219) );
  INV_X1 U617 ( .A(G82), .ZN(G220) );
  INV_X1 U618 ( .A(G69), .ZN(G235) );
  INV_X1 U619 ( .A(G57), .ZN(G237) );
  NAND2_X1 U620 ( .A1(n653), .A2(G52), .ZN(n556) );
  NAND2_X1 U621 ( .A1(G64), .A2(n652), .ZN(n555) );
  NAND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n561) );
  NAND2_X1 U623 ( .A1(G77), .A2(n639), .ZN(n558) );
  NAND2_X1 U624 ( .A1(G90), .A2(n640), .ZN(n557) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U626 ( .A(KEYINPUT9), .B(n559), .Z(n560) );
  NOR2_X1 U627 ( .A1(n561), .A2(n560), .ZN(G171) );
  XNOR2_X1 U628 ( .A(KEYINPUT7), .B(KEYINPUT76), .ZN(n575) );
  XOR2_X1 U629 ( .A(KEYINPUT4), .B(KEYINPUT74), .Z(n563) );
  NAND2_X1 U630 ( .A1(G89), .A2(n640), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U632 ( .A(KEYINPUT73), .B(n564), .ZN(n566) );
  NAND2_X1 U633 ( .A1(n639), .A2(G76), .ZN(n565) );
  NAND2_X1 U634 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n567), .B(KEYINPUT5), .ZN(n573) );
  XNOR2_X1 U636 ( .A(KEYINPUT75), .B(KEYINPUT6), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n653), .A2(G51), .ZN(n569) );
  NAND2_X1 U638 ( .A1(G63), .A2(n652), .ZN(n568) );
  NAND2_X1 U639 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U640 ( .A(n571), .B(n570), .ZN(n572) );
  NAND2_X1 U641 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n575), .B(n574), .ZN(G168) );
  XOR2_X1 U643 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U644 ( .A1(G94), .A2(G452), .ZN(n576) );
  XNOR2_X1 U645 ( .A(n576), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U646 ( .A1(G7), .A2(G661), .ZN(n577) );
  XNOR2_X1 U647 ( .A(n577), .B(KEYINPUT70), .ZN(n578) );
  XNOR2_X1 U648 ( .A(KEYINPUT10), .B(n578), .ZN(G223) );
  INV_X1 U649 ( .A(G223), .ZN(n841) );
  NAND2_X1 U650 ( .A1(n841), .A2(G567), .ZN(n579) );
  XOR2_X1 U651 ( .A(KEYINPUT11), .B(n579), .Z(G234) );
  NAND2_X1 U652 ( .A1(G81), .A2(n640), .ZN(n580) );
  XNOR2_X1 U653 ( .A(n580), .B(KEYINPUT12), .ZN(n582) );
  NAND2_X1 U654 ( .A1(G68), .A2(n639), .ZN(n581) );
  NAND2_X1 U655 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U656 ( .A(KEYINPUT13), .B(n583), .ZN(n589) );
  NAND2_X1 U657 ( .A1(n652), .A2(G56), .ZN(n584) );
  XOR2_X1 U658 ( .A(KEYINPUT14), .B(n584), .Z(n587) );
  NAND2_X1 U659 ( .A1(G43), .A2(n653), .ZN(n585) );
  XNOR2_X1 U660 ( .A(KEYINPUT71), .B(n585), .ZN(n586) );
  NOR2_X1 U661 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U662 ( .A1(n589), .A2(n588), .ZN(n1013) );
  INV_X1 U663 ( .A(G860), .ZN(n623) );
  OR2_X1 U664 ( .A1(n1013), .A2(n623), .ZN(G153) );
  INV_X1 U665 ( .A(G171), .ZN(G301) );
  NAND2_X1 U666 ( .A1(G79), .A2(n639), .ZN(n591) );
  NAND2_X1 U667 ( .A1(G92), .A2(n640), .ZN(n590) );
  NAND2_X1 U668 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U669 ( .A1(n653), .A2(G54), .ZN(n593) );
  NAND2_X1 U670 ( .A1(G66), .A2(n652), .ZN(n592) );
  NAND2_X1 U671 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U672 ( .A1(n595), .A2(n594), .ZN(n597) );
  XNOR2_X1 U673 ( .A(KEYINPUT72), .B(KEYINPUT15), .ZN(n596) );
  XNOR2_X2 U674 ( .A(n597), .B(n596), .ZN(n1018) );
  NOR2_X1 U675 ( .A1(n1018), .A2(G868), .ZN(n599) );
  INV_X1 U676 ( .A(G868), .ZN(n600) );
  NOR2_X1 U677 ( .A1(n600), .A2(G301), .ZN(n598) );
  NOR2_X1 U678 ( .A1(n599), .A2(n598), .ZN(G284) );
  NAND2_X1 U679 ( .A1(G868), .A2(G286), .ZN(n602) );
  NAND2_X1 U680 ( .A1(G299), .A2(n600), .ZN(n601) );
  NAND2_X1 U681 ( .A1(n602), .A2(n601), .ZN(G297) );
  NAND2_X1 U682 ( .A1(n623), .A2(G559), .ZN(n603) );
  INV_X1 U683 ( .A(n1018), .ZN(n621) );
  NAND2_X1 U684 ( .A1(n603), .A2(n621), .ZN(n604) );
  XNOR2_X1 U685 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U686 ( .A1(G868), .A2(n1013), .ZN(n607) );
  NAND2_X1 U687 ( .A1(n621), .A2(G868), .ZN(n605) );
  NOR2_X1 U688 ( .A1(G559), .A2(n605), .ZN(n606) );
  NOR2_X1 U689 ( .A1(n607), .A2(n606), .ZN(G282) );
  NAND2_X1 U690 ( .A1(G111), .A2(n894), .ZN(n609) );
  NAND2_X1 U691 ( .A1(G99), .A2(n898), .ZN(n608) );
  NAND2_X1 U692 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U693 ( .A(n610), .B(KEYINPUT77), .ZN(n613) );
  BUF_X1 U694 ( .A(n611), .Z(n899) );
  NAND2_X1 U695 ( .A1(G135), .A2(n899), .ZN(n612) );
  NAND2_X1 U696 ( .A1(n613), .A2(n612), .ZN(n616) );
  NAND2_X1 U697 ( .A1(n895), .A2(G123), .ZN(n614) );
  XOR2_X1 U698 ( .A(KEYINPUT18), .B(n614), .Z(n615) );
  NOR2_X1 U699 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U700 ( .A(KEYINPUT78), .B(n617), .ZN(n978) );
  XOR2_X1 U701 ( .A(G2096), .B(KEYINPUT79), .Z(n618) );
  XNOR2_X1 U702 ( .A(n978), .B(n618), .ZN(n620) );
  INV_X1 U703 ( .A(G2100), .ZN(n619) );
  NAND2_X1 U704 ( .A1(n620), .A2(n619), .ZN(G156) );
  NAND2_X1 U705 ( .A1(n621), .A2(G559), .ZN(n622) );
  XOR2_X1 U706 ( .A(n1013), .B(n622), .Z(n662) );
  NAND2_X1 U707 ( .A1(n623), .A2(n662), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n653), .A2(G55), .ZN(n625) );
  NAND2_X1 U709 ( .A1(G67), .A2(n652), .ZN(n624) );
  NAND2_X1 U710 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U711 ( .A1(G80), .A2(n639), .ZN(n627) );
  NAND2_X1 U712 ( .A1(G93), .A2(n640), .ZN(n626) );
  NAND2_X1 U713 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U714 ( .A1(n629), .A2(n628), .ZN(n664) );
  XOR2_X1 U715 ( .A(n630), .B(n664), .Z(G145) );
  NAND2_X1 U716 ( .A1(n653), .A2(G48), .ZN(n637) );
  NAND2_X1 U717 ( .A1(G86), .A2(n640), .ZN(n632) );
  NAND2_X1 U718 ( .A1(G61), .A2(n652), .ZN(n631) );
  NAND2_X1 U719 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U720 ( .A1(G73), .A2(n639), .ZN(n633) );
  XOR2_X1 U721 ( .A(KEYINPUT2), .B(n633), .Z(n634) );
  NOR2_X1 U722 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U723 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U724 ( .A(n638), .B(KEYINPUT80), .ZN(G305) );
  NAND2_X1 U725 ( .A1(G75), .A2(n639), .ZN(n642) );
  NAND2_X1 U726 ( .A1(G88), .A2(n640), .ZN(n641) );
  NAND2_X1 U727 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n653), .A2(G50), .ZN(n644) );
  NAND2_X1 U729 ( .A1(G62), .A2(n652), .ZN(n643) );
  NAND2_X1 U730 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U731 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U732 ( .A(KEYINPUT81), .B(n647), .Z(G166) );
  NAND2_X1 U733 ( .A1(G74), .A2(G651), .ZN(n650) );
  NAND2_X1 U734 ( .A1(G87), .A2(n648), .ZN(n649) );
  NAND2_X1 U735 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U736 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U737 ( .A1(n653), .A2(G49), .ZN(n654) );
  NAND2_X1 U738 ( .A1(n655), .A2(n654), .ZN(G288) );
  XNOR2_X1 U739 ( .A(KEYINPUT19), .B(KEYINPUT82), .ZN(n656) );
  XNOR2_X1 U740 ( .A(n656), .B(n664), .ZN(n659) );
  XNOR2_X1 U741 ( .A(G166), .B(G299), .ZN(n657) );
  XNOR2_X1 U742 ( .A(n657), .B(G290), .ZN(n658) );
  XNOR2_X1 U743 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U744 ( .A(n660), .B(G288), .ZN(n661) );
  XNOR2_X1 U745 ( .A(G305), .B(n661), .ZN(n914) );
  XNOR2_X1 U746 ( .A(n662), .B(n914), .ZN(n663) );
  NAND2_X1 U747 ( .A1(n663), .A2(G868), .ZN(n666) );
  OR2_X1 U748 ( .A1(G868), .A2(n664), .ZN(n665) );
  NAND2_X1 U749 ( .A1(n666), .A2(n665), .ZN(G295) );
  NAND2_X1 U750 ( .A1(G2078), .A2(G2084), .ZN(n667) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n667), .Z(n668) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n668), .ZN(n670) );
  XOR2_X1 U753 ( .A(KEYINPUT21), .B(KEYINPUT83), .Z(n669) );
  XNOR2_X1 U754 ( .A(n670), .B(n669), .ZN(n671) );
  NAND2_X1 U755 ( .A1(G2072), .A2(n671), .ZN(G158) );
  XNOR2_X1 U756 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U757 ( .A1(G237), .A2(G235), .ZN(n672) );
  NAND2_X1 U758 ( .A1(G120), .A2(n672), .ZN(n673) );
  XNOR2_X1 U759 ( .A(KEYINPUT85), .B(n673), .ZN(n674) );
  NAND2_X1 U760 ( .A1(n674), .A2(G108), .ZN(n845) );
  NAND2_X1 U761 ( .A1(n845), .A2(G567), .ZN(n680) );
  NOR2_X1 U762 ( .A1(G220), .A2(G219), .ZN(n675) );
  XNOR2_X1 U763 ( .A(KEYINPUT22), .B(n675), .ZN(n676) );
  NAND2_X1 U764 ( .A1(n676), .A2(G96), .ZN(n677) );
  NOR2_X1 U765 ( .A1(G218), .A2(n677), .ZN(n678) );
  XOR2_X1 U766 ( .A(KEYINPUT84), .B(n678), .Z(n846) );
  NAND2_X1 U767 ( .A1(n846), .A2(G2106), .ZN(n679) );
  NAND2_X1 U768 ( .A1(n680), .A2(n679), .ZN(n847) );
  NAND2_X1 U769 ( .A1(G661), .A2(G483), .ZN(n681) );
  XNOR2_X1 U770 ( .A(KEYINPUT86), .B(n681), .ZN(n682) );
  NOR2_X1 U771 ( .A1(n847), .A2(n682), .ZN(n844) );
  NAND2_X1 U772 ( .A1(n844), .A2(G36), .ZN(G176) );
  XOR2_X1 U773 ( .A(KEYINPUT88), .B(G166), .Z(G303) );
  NAND2_X1 U774 ( .A1(G160), .A2(G40), .ZN(n776) );
  INV_X1 U775 ( .A(n776), .ZN(n683) );
  INV_X1 U776 ( .A(G2072), .ZN(n989) );
  XNOR2_X1 U777 ( .A(KEYINPUT27), .B(KEYINPUT94), .ZN(n684) );
  XNOR2_X1 U778 ( .A(n685), .B(n684), .ZN(n687) );
  NAND2_X1 U779 ( .A1(n732), .A2(G1956), .ZN(n686) );
  NAND2_X1 U780 ( .A1(n687), .A2(n686), .ZN(n709) );
  XNOR2_X1 U781 ( .A(n688), .B(KEYINPUT96), .ZN(n693) );
  NAND2_X1 U782 ( .A1(G1348), .A2(n732), .ZN(n690) );
  NAND2_X1 U783 ( .A1(n714), .A2(G2067), .ZN(n689) );
  NAND2_X1 U784 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U785 ( .A1(n691), .A2(n1018), .ZN(n692) );
  NOR2_X1 U786 ( .A1(n693), .A2(n692), .ZN(n708) );
  INV_X1 U787 ( .A(G1341), .ZN(n694) );
  NAND2_X1 U788 ( .A1(n1018), .A2(G1348), .ZN(n1011) );
  NAND2_X1 U789 ( .A1(n694), .A2(n1011), .ZN(n695) );
  NAND2_X1 U790 ( .A1(n732), .A2(n695), .ZN(n698) );
  NAND2_X1 U791 ( .A1(n714), .A2(G1996), .ZN(n696) );
  XNOR2_X1 U792 ( .A(KEYINPUT26), .B(KEYINPUT95), .ZN(n700) );
  NAND2_X1 U793 ( .A1(n696), .A2(n700), .ZN(n697) );
  NAND2_X1 U794 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U795 ( .A1(n1013), .A2(n699), .ZN(n706) );
  NAND2_X1 U796 ( .A1(n1018), .A2(G2067), .ZN(n703) );
  INV_X1 U797 ( .A(n700), .ZN(n701) );
  NAND2_X1 U798 ( .A1(n701), .A2(G1996), .ZN(n702) );
  NAND2_X1 U799 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U800 ( .A1(n704), .A2(n714), .ZN(n705) );
  NAND2_X1 U801 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U802 ( .A1(n708), .A2(n707), .ZN(n712) );
  NAND2_X1 U803 ( .A1(G299), .A2(n709), .ZN(n710) );
  XNOR2_X1 U804 ( .A(KEYINPUT28), .B(n710), .ZN(n711) );
  NAND2_X1 U805 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U806 ( .A(n713), .B(KEYINPUT29), .ZN(n718) );
  NAND2_X1 U807 ( .A1(G1961), .A2(n732), .ZN(n716) );
  XOR2_X1 U808 ( .A(KEYINPUT25), .B(G2078), .Z(n956) );
  NAND2_X1 U809 ( .A1(n714), .A2(n956), .ZN(n715) );
  NAND2_X1 U810 ( .A1(n716), .A2(n715), .ZN(n719) );
  NOR2_X1 U811 ( .A1(G301), .A2(n719), .ZN(n717) );
  NOR2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n731) );
  AND2_X1 U813 ( .A1(G301), .A2(n719), .ZN(n726) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n775), .ZN(n746) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n720), .ZN(n743) );
  INV_X1 U816 ( .A(G8), .ZN(n721) );
  OR2_X1 U817 ( .A1(n743), .A2(n721), .ZN(n722) );
  OR2_X1 U818 ( .A1(n746), .A2(n722), .ZN(n723) );
  XNOR2_X1 U819 ( .A(n723), .B(KEYINPUT30), .ZN(n724) );
  NOR2_X1 U820 ( .A1(n724), .A2(G168), .ZN(n725) );
  NOR2_X1 U821 ( .A1(n726), .A2(n725), .ZN(n729) );
  OR2_X2 U822 ( .A1(n731), .A2(n730), .ZN(n744) );
  NAND2_X1 U823 ( .A1(n744), .A2(G286), .ZN(n740) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n732), .ZN(n733) );
  XOR2_X1 U825 ( .A(KEYINPUT99), .B(n733), .Z(n736) );
  NOR2_X1 U826 ( .A1(G1971), .A2(n775), .ZN(n734) );
  XNOR2_X1 U827 ( .A(n734), .B(KEYINPUT98), .ZN(n735) );
  NOR2_X1 U828 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U829 ( .A1(G303), .A2(n737), .ZN(n738) );
  OR2_X1 U830 ( .A1(n721), .A2(n738), .ZN(n739) );
  NAND2_X1 U831 ( .A1(n743), .A2(G8), .ZN(n748) );
  INV_X1 U832 ( .A(n744), .ZN(n745) );
  NOR2_X1 U833 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U834 ( .A1(n748), .A2(n747), .ZN(n765) );
  NAND2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n1023) );
  AND2_X1 U836 ( .A1(n765), .A2(n1023), .ZN(n749) );
  NAND2_X1 U837 ( .A1(n764), .A2(n749), .ZN(n754) );
  INV_X1 U838 ( .A(n1023), .ZN(n752) );
  NOR2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n1021) );
  NOR2_X1 U840 ( .A1(G303), .A2(G1971), .ZN(n1020) );
  XOR2_X1 U841 ( .A(n1020), .B(KEYINPUT101), .Z(n750) );
  NOR2_X1 U842 ( .A1(n1021), .A2(n750), .ZN(n751) );
  OR2_X1 U843 ( .A1(n752), .A2(n751), .ZN(n753) );
  AND2_X1 U844 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U845 ( .A1(n775), .A2(n755), .ZN(n756) );
  NOR2_X1 U846 ( .A1(KEYINPUT33), .A2(n756), .ZN(n760) );
  NAND2_X1 U847 ( .A1(KEYINPUT33), .A2(n1021), .ZN(n757) );
  NOR2_X1 U848 ( .A1(n775), .A2(n757), .ZN(n758) );
  XNOR2_X1 U849 ( .A(n758), .B(KEYINPUT102), .ZN(n759) );
  NOR2_X2 U850 ( .A1(n760), .A2(n759), .ZN(n762) );
  XNOR2_X1 U851 ( .A(n762), .B(n761), .ZN(n763) );
  XOR2_X1 U852 ( .A(G305), .B(G1981), .Z(n1004) );
  NAND2_X1 U853 ( .A1(n763), .A2(n1004), .ZN(n771) );
  NAND2_X1 U854 ( .A1(n765), .A2(n764), .ZN(n768) );
  NOR2_X1 U855 ( .A1(G2090), .A2(G303), .ZN(n766) );
  NAND2_X1 U856 ( .A1(G8), .A2(n766), .ZN(n767) );
  NAND2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U858 ( .A1(n769), .A2(n775), .ZN(n770) );
  NAND2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U860 ( .A(n772), .B(KEYINPUT104), .ZN(n818) );
  NOR2_X1 U861 ( .A1(G305), .A2(G1981), .ZN(n773) );
  XOR2_X1 U862 ( .A(n773), .B(KEYINPUT24), .Z(n774) );
  NOR2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n816) );
  NOR2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n823) );
  NAND2_X1 U865 ( .A1(n898), .A2(G104), .ZN(n779) );
  NAND2_X1 U866 ( .A1(G140), .A2(n899), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U868 ( .A(KEYINPUT34), .B(n780), .ZN(n785) );
  NAND2_X1 U869 ( .A1(G116), .A2(n894), .ZN(n782) );
  NAND2_X1 U870 ( .A1(G128), .A2(n895), .ZN(n781) );
  NAND2_X1 U871 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U872 ( .A(n783), .B(KEYINPUT35), .Z(n784) );
  NOR2_X1 U873 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U874 ( .A(KEYINPUT36), .B(n786), .Z(n787) );
  XNOR2_X1 U875 ( .A(KEYINPUT89), .B(n787), .ZN(n891) );
  XNOR2_X1 U876 ( .A(G2067), .B(KEYINPUT37), .ZN(n812) );
  NOR2_X1 U877 ( .A1(n891), .A2(n812), .ZN(n983) );
  NAND2_X1 U878 ( .A1(n823), .A2(n983), .ZN(n820) );
  NAND2_X1 U879 ( .A1(G129), .A2(n895), .ZN(n789) );
  NAND2_X1 U880 ( .A1(G141), .A2(n899), .ZN(n788) );
  NAND2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U882 ( .A1(n898), .A2(G105), .ZN(n790) );
  XOR2_X1 U883 ( .A(KEYINPUT38), .B(n790), .Z(n791) );
  NOR2_X1 U884 ( .A1(n792), .A2(n791), .ZN(n794) );
  NAND2_X1 U885 ( .A1(n894), .A2(G117), .ZN(n793) );
  NAND2_X1 U886 ( .A1(n794), .A2(n793), .ZN(n905) );
  NOR2_X1 U887 ( .A1(G1996), .A2(n905), .ZN(n974) );
  NAND2_X1 U888 ( .A1(G1996), .A2(n905), .ZN(n804) );
  NAND2_X1 U889 ( .A1(G95), .A2(n898), .ZN(n795) );
  XNOR2_X1 U890 ( .A(n795), .B(KEYINPUT90), .ZN(n802) );
  NAND2_X1 U891 ( .A1(G107), .A2(n894), .ZN(n797) );
  NAND2_X1 U892 ( .A1(G119), .A2(n895), .ZN(n796) );
  NAND2_X1 U893 ( .A1(n797), .A2(n796), .ZN(n800) );
  NAND2_X1 U894 ( .A1(G131), .A2(n899), .ZN(n798) );
  XNOR2_X1 U895 ( .A(KEYINPUT91), .B(n798), .ZN(n799) );
  NOR2_X1 U896 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U897 ( .A1(n802), .A2(n801), .ZN(n887) );
  NAND2_X1 U898 ( .A1(G1991), .A2(n887), .ZN(n803) );
  NAND2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n979) );
  NAND2_X1 U900 ( .A1(n979), .A2(n823), .ZN(n805) );
  XOR2_X1 U901 ( .A(KEYINPUT92), .B(n805), .Z(n819) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n806) );
  NOR2_X1 U903 ( .A1(G1991), .A2(n887), .ZN(n977) );
  NOR2_X1 U904 ( .A1(n806), .A2(n977), .ZN(n807) );
  NOR2_X1 U905 ( .A1(n819), .A2(n807), .ZN(n808) );
  NOR2_X1 U906 ( .A1(n974), .A2(n808), .ZN(n809) );
  XOR2_X1 U907 ( .A(n809), .B(KEYINPUT105), .Z(n810) );
  XNOR2_X1 U908 ( .A(KEYINPUT39), .B(n810), .ZN(n811) );
  NAND2_X1 U909 ( .A1(n820), .A2(n811), .ZN(n813) );
  NAND2_X1 U910 ( .A1(n891), .A2(n812), .ZN(n994) );
  NAND2_X1 U911 ( .A1(n813), .A2(n994), .ZN(n814) );
  NAND2_X1 U912 ( .A1(n814), .A2(n823), .ZN(n815) );
  XOR2_X1 U913 ( .A(KEYINPUT106), .B(n815), .Z(n827) );
  OR2_X1 U914 ( .A1(n816), .A2(n827), .ZN(n817) );
  NOR2_X1 U915 ( .A1(n818), .A2(n817), .ZN(n829) );
  INV_X1 U916 ( .A(n819), .ZN(n821) );
  NAND2_X1 U917 ( .A1(n821), .A2(n820), .ZN(n822) );
  XOR2_X1 U918 ( .A(KEYINPUT93), .B(n822), .Z(n825) );
  XNOR2_X1 U919 ( .A(G1986), .B(G290), .ZN(n1010) );
  AND2_X1 U920 ( .A1(n1010), .A2(n823), .ZN(n824) );
  NOR2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U923 ( .A(n830), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U924 ( .A(G2454), .B(G2435), .Z(n832) );
  XNOR2_X1 U925 ( .A(G2438), .B(G2427), .ZN(n831) );
  XNOR2_X1 U926 ( .A(n832), .B(n831), .ZN(n839) );
  XOR2_X1 U927 ( .A(KEYINPUT107), .B(G2446), .Z(n834) );
  XNOR2_X1 U928 ( .A(G2443), .B(G2430), .ZN(n833) );
  XNOR2_X1 U929 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U930 ( .A(n835), .B(G2451), .Z(n837) );
  XNOR2_X1 U931 ( .A(G1341), .B(G1348), .ZN(n836) );
  XNOR2_X1 U932 ( .A(n837), .B(n836), .ZN(n838) );
  XNOR2_X1 U933 ( .A(n839), .B(n838), .ZN(n840) );
  NAND2_X1 U934 ( .A1(n840), .A2(G14), .ZN(n919) );
  XOR2_X1 U935 ( .A(KEYINPUT108), .B(n919), .Z(G401) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n841), .ZN(G217) );
  AND2_X1 U937 ( .A1(G15), .A2(G2), .ZN(n842) );
  NAND2_X1 U938 ( .A1(G661), .A2(n842), .ZN(G259) );
  NAND2_X1 U939 ( .A1(G3), .A2(G1), .ZN(n843) );
  NAND2_X1 U940 ( .A1(n844), .A2(n843), .ZN(G188) );
  XNOR2_X1 U941 ( .A(G120), .B(KEYINPUT109), .ZN(G236) );
  INV_X1 U943 ( .A(G108), .ZN(G238) );
  INV_X1 U944 ( .A(G96), .ZN(G221) );
  NOR2_X1 U945 ( .A1(n846), .A2(n845), .ZN(G325) );
  INV_X1 U946 ( .A(G325), .ZN(G261) );
  INV_X1 U947 ( .A(n847), .ZN(G319) );
  XOR2_X1 U948 ( .A(G1966), .B(G1956), .Z(n849) );
  XNOR2_X1 U949 ( .A(G1981), .B(G1971), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n859) );
  XOR2_X1 U951 ( .A(KEYINPUT111), .B(KEYINPUT41), .Z(n851) );
  XNOR2_X1 U952 ( .A(G1996), .B(KEYINPUT113), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U954 ( .A(G1991), .B(G1986), .Z(n853) );
  XNOR2_X1 U955 ( .A(G1976), .B(G1961), .ZN(n852) );
  XNOR2_X1 U956 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U957 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U958 ( .A(KEYINPUT112), .B(G2474), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U960 ( .A(n859), .B(n858), .Z(G229) );
  XOR2_X1 U961 ( .A(G2096), .B(KEYINPUT43), .Z(n861) );
  XNOR2_X1 U962 ( .A(G2090), .B(KEYINPUT110), .ZN(n860) );
  XNOR2_X1 U963 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U964 ( .A(n862), .B(G2678), .Z(n864) );
  XNOR2_X1 U965 ( .A(G2067), .B(G2072), .ZN(n863) );
  XNOR2_X1 U966 ( .A(n864), .B(n863), .ZN(n868) );
  XOR2_X1 U967 ( .A(KEYINPUT42), .B(G2100), .Z(n866) );
  XNOR2_X1 U968 ( .A(G2078), .B(G2084), .ZN(n865) );
  XNOR2_X1 U969 ( .A(n866), .B(n865), .ZN(n867) );
  XNOR2_X1 U970 ( .A(n868), .B(n867), .ZN(G227) );
  NAND2_X1 U971 ( .A1(G124), .A2(n895), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n869), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n894), .A2(G112), .ZN(n870) );
  NAND2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n875) );
  NAND2_X1 U975 ( .A1(n898), .A2(G100), .ZN(n873) );
  NAND2_X1 U976 ( .A1(G136), .A2(n899), .ZN(n872) );
  NAND2_X1 U977 ( .A1(n873), .A2(n872), .ZN(n874) );
  NOR2_X1 U978 ( .A1(n875), .A2(n874), .ZN(G162) );
  XOR2_X1 U979 ( .A(KEYINPUT116), .B(KEYINPUT48), .Z(n877) );
  XNOR2_X1 U980 ( .A(G160), .B(KEYINPUT46), .ZN(n876) );
  XNOR2_X1 U981 ( .A(n877), .B(n876), .ZN(n890) );
  NAND2_X1 U982 ( .A1(G115), .A2(n894), .ZN(n879) );
  NAND2_X1 U983 ( .A1(G127), .A2(n895), .ZN(n878) );
  NAND2_X1 U984 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U985 ( .A(KEYINPUT47), .B(n880), .ZN(n886) );
  NAND2_X1 U986 ( .A1(n899), .A2(G139), .ZN(n881) );
  XNOR2_X1 U987 ( .A(n881), .B(KEYINPUT115), .ZN(n884) );
  NAND2_X1 U988 ( .A1(G103), .A2(n898), .ZN(n882) );
  XOR2_X1 U989 ( .A(KEYINPUT114), .B(n882), .Z(n883) );
  NOR2_X1 U990 ( .A1(n884), .A2(n883), .ZN(n885) );
  NAND2_X1 U991 ( .A1(n886), .A2(n885), .ZN(n987) );
  XOR2_X1 U992 ( .A(n887), .B(n987), .Z(n888) );
  XNOR2_X1 U993 ( .A(n978), .B(n888), .ZN(n889) );
  XNOR2_X1 U994 ( .A(n890), .B(n889), .ZN(n893) );
  XNOR2_X1 U995 ( .A(n891), .B(G162), .ZN(n892) );
  XNOR2_X1 U996 ( .A(n893), .B(n892), .ZN(n909) );
  NAND2_X1 U997 ( .A1(G118), .A2(n894), .ZN(n897) );
  NAND2_X1 U998 ( .A1(G130), .A2(n895), .ZN(n896) );
  NAND2_X1 U999 ( .A1(n897), .A2(n896), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(n898), .A2(G106), .ZN(n901) );
  NAND2_X1 U1001 ( .A1(G142), .A2(n899), .ZN(n900) );
  NAND2_X1 U1002 ( .A1(n901), .A2(n900), .ZN(n902) );
  XOR2_X1 U1003 ( .A(n902), .B(KEYINPUT45), .Z(n903) );
  NOR2_X1 U1004 ( .A1(n904), .A2(n903), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1006 ( .A(G164), .B(n907), .Z(n908) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n910), .ZN(n911) );
  XOR2_X1 U1009 ( .A(KEYINPUT117), .B(n911), .Z(G395) );
  XNOR2_X1 U1010 ( .A(n1018), .B(KEYINPUT118), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(G286), .B(G171), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(n913), .B(n912), .ZN(n916) );
  XOR2_X1 U1013 ( .A(n1013), .B(n914), .Z(n915) );
  XNOR2_X1 U1014 ( .A(n916), .B(n915), .ZN(n917) );
  NOR2_X1 U1015 ( .A1(G37), .A2(n917), .ZN(n918) );
  XOR2_X1 U1016 ( .A(KEYINPUT119), .B(n918), .Z(G397) );
  NAND2_X1 U1017 ( .A1(G319), .A2(n919), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(G229), .A2(G227), .ZN(n920) );
  XNOR2_X1 U1019 ( .A(KEYINPUT49), .B(n920), .ZN(n921) );
  NOR2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1024 ( .A(G1971), .B(G22), .Z(n927) );
  XNOR2_X1 U1025 ( .A(G1976), .B(KEYINPUT127), .ZN(n925) );
  XNOR2_X1 U1026 ( .A(n925), .B(G23), .ZN(n926) );
  NAND2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n929) );
  XNOR2_X1 U1028 ( .A(G24), .B(G1986), .ZN(n928) );
  NOR2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1030 ( .A(KEYINPUT58), .B(n930), .Z(n947) );
  XOR2_X1 U1031 ( .A(G1966), .B(G21), .Z(n941) );
  XOR2_X1 U1032 ( .A(KEYINPUT125), .B(G4), .Z(n932) );
  XNOR2_X1 U1033 ( .A(G1348), .B(KEYINPUT59), .ZN(n931) );
  XNOR2_X1 U1034 ( .A(n932), .B(n931), .ZN(n936) );
  XNOR2_X1 U1035 ( .A(G1981), .B(G6), .ZN(n934) );
  XNOR2_X1 U1036 ( .A(G1341), .B(G19), .ZN(n933) );
  NOR2_X1 U1037 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1038 ( .A1(n936), .A2(n935), .ZN(n938) );
  XNOR2_X1 U1039 ( .A(G20), .B(G1956), .ZN(n937) );
  NOR2_X1 U1040 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1041 ( .A(KEYINPUT60), .B(n939), .ZN(n940) );
  NAND2_X1 U1042 ( .A1(n941), .A2(n940), .ZN(n944) );
  XNOR2_X1 U1043 ( .A(KEYINPUT124), .B(G1961), .ZN(n942) );
  XNOR2_X1 U1044 ( .A(G5), .B(n942), .ZN(n943) );
  NOR2_X1 U1045 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1046 ( .A(KEYINPUT126), .B(n945), .Z(n946) );
  NOR2_X1 U1047 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1048 ( .A(KEYINPUT61), .B(n948), .Z(n949) );
  NOR2_X1 U1049 ( .A1(G16), .A2(n949), .ZN(n972) );
  INV_X1 U1050 ( .A(KEYINPUT55), .ZN(n999) );
  XNOR2_X1 U1051 ( .A(G2084), .B(G34), .ZN(n950) );
  XNOR2_X1 U1052 ( .A(n950), .B(KEYINPUT54), .ZN(n952) );
  XNOR2_X1 U1053 ( .A(G35), .B(G2090), .ZN(n951) );
  NOR2_X1 U1054 ( .A1(n952), .A2(n951), .ZN(n966) );
  XOR2_X1 U1055 ( .A(KEYINPUT53), .B(KEYINPUT123), .Z(n964) );
  XOR2_X1 U1056 ( .A(G1991), .B(G25), .Z(n953) );
  NAND2_X1 U1057 ( .A1(n953), .A2(G28), .ZN(n962) );
  XNOR2_X1 U1058 ( .A(G1996), .B(G32), .ZN(n955) );
  XNOR2_X1 U1059 ( .A(G33), .B(G2072), .ZN(n954) );
  NOR2_X1 U1060 ( .A1(n955), .A2(n954), .ZN(n960) );
  XNOR2_X1 U1061 ( .A(n956), .B(G27), .ZN(n958) );
  XNOR2_X1 U1062 ( .A(G2067), .B(G26), .ZN(n957) );
  NOR2_X1 U1063 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1064 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1065 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1066 ( .A(n964), .B(n963), .Z(n965) );
  NAND2_X1 U1067 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1068 ( .A(n999), .B(n967), .ZN(n969) );
  INV_X1 U1069 ( .A(G29), .ZN(n968) );
  NAND2_X1 U1070 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1071 ( .A1(G11), .A2(n970), .ZN(n971) );
  NOR2_X1 U1072 ( .A1(n972), .A2(n971), .ZN(n1003) );
  XOR2_X1 U1073 ( .A(G2090), .B(G162), .Z(n973) );
  NOR2_X1 U1074 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1075 ( .A(KEYINPUT51), .B(n975), .Z(n986) );
  XOR2_X1 U1076 ( .A(G2084), .B(G160), .Z(n976) );
  NOR2_X1 U1077 ( .A1(n977), .A2(n976), .ZN(n981) );
  NOR2_X1 U1078 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1079 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1080 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1081 ( .A(n984), .B(KEYINPUT120), .ZN(n985) );
  NAND2_X1 U1082 ( .A1(n986), .A2(n985), .ZN(n997) );
  XOR2_X1 U1083 ( .A(G164), .B(G2078), .Z(n991) );
  XNOR2_X1 U1084 ( .A(KEYINPUT121), .B(n987), .ZN(n988) );
  XNOR2_X1 U1085 ( .A(n989), .B(n988), .ZN(n990) );
  NOR2_X1 U1086 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1087 ( .A(KEYINPUT122), .B(n992), .ZN(n993) );
  XNOR2_X1 U1088 ( .A(n993), .B(KEYINPUT50), .ZN(n995) );
  NAND2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1091 ( .A(KEYINPUT52), .B(n998), .ZN(n1000) );
  NAND2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1001), .A2(G29), .ZN(n1002) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1033) );
  XOR2_X1 U1095 ( .A(G16), .B(KEYINPUT56), .Z(n1031) );
  XNOR2_X1 U1096 ( .A(G168), .B(G1966), .ZN(n1005) );
  NAND2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1098 ( .A(n1006), .B(KEYINPUT57), .ZN(n1017) );
  XNOR2_X1 U1099 ( .A(G1961), .B(G171), .ZN(n1008) );
  NAND2_X1 U1100 ( .A1(G1971), .A2(G303), .ZN(n1007) );
  NAND2_X1 U1101 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  NAND2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1015) );
  XNOR2_X1 U1104 ( .A(G1341), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1029) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(G1348), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1027) );
  INV_X1 U1109 ( .A(n1021), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1025) );
  XNOR2_X1 U1111 ( .A(G1956), .B(G299), .ZN(n1024) );
  NOR2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1115 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1116 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1117 ( .A(n1034), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1118 ( .A(G311), .ZN(G150) );
endmodule

