//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT65), .Z(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT66), .B(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G107), .A2(G264), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n209), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT67), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n222), .A2(new_n207), .ZN(new_n223));
  NOR2_X1   g0023(.A1(G58), .A2(G68), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n225), .A3(G50), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n209), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT0), .ZN(new_n229));
  NAND4_X1  g0029(.A1(new_n220), .A2(new_n221), .A3(new_n226), .A4(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT68), .Z(G361));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT69), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G13), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n248), .A2(G1), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G20), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n222), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n207), .A2(G1), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(G50), .A3(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G50), .B2(new_n250), .ZN(new_n258));
  INV_X1    g0058(.A(new_n253), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n202), .A2(G20), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT8), .B(G58), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G20), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n262), .A2(new_n264), .B1(G150), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n259), .B1(new_n260), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n258), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT70), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  INV_X1    g0072(.A(new_n222), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n273), .A2(new_n274), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n278), .A2(new_n269), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n277), .B1(G226), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT71), .ZN(new_n281));
  AND2_X1   g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NOR2_X1   g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT3), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n263), .ZN(new_n286));
  NAND2_X1  g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(KEYINPUT71), .A3(new_n287), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(KEYINPUT72), .A2(G1698), .ZN(new_n290));
  NOR2_X1   g0090(.A1(KEYINPUT72), .A2(G1698), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n289), .A2(G222), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G77), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n293), .B1(new_n294), .B2(new_n289), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n289), .A2(KEYINPUT73), .A3(G1698), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n284), .A2(new_n288), .A3(G1698), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT73), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n295), .B1(G223), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n280), .B1(new_n301), .B2(new_n278), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n268), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AND2_X1   g0104(.A1(KEYINPUT74), .A2(G179), .ZN(new_n305));
  NOR2_X1   g0105(.A1(KEYINPUT74), .A2(G179), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n304), .B1(new_n308), .B2(new_n302), .ZN(new_n309));
  AND3_X1   g0109(.A1(new_n251), .A2(KEYINPUT75), .A3(new_n294), .ZN(new_n310));
  AOI21_X1  g0110(.A(KEYINPUT75), .B1(new_n251), .B2(new_n294), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n262), .A2(new_n265), .B1(G20), .B2(G77), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT15), .B(G87), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n264), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n259), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  NOR4_X1   g0117(.A1(new_n251), .A2(new_n253), .A3(new_n294), .A4(new_n255), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n312), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n210), .B1(new_n296), .B2(new_n299), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n284), .A2(new_n288), .A3(G232), .A4(new_n292), .ZN(new_n322));
  INV_X1    g0122(.A(G107), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n322), .B1(new_n289), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n320), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n277), .B1(G244), .B2(new_n279), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n319), .B1(new_n327), .B2(new_n303), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n325), .A2(new_n307), .A3(new_n326), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G190), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n319), .B1(new_n327), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G200), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n325), .B2(new_n326), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g0136(.A(G190), .B(new_n280), .C1(new_n301), .C2(new_n278), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT76), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n268), .B(KEYINPUT9), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n339), .B1(new_n302), .B2(G200), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n341), .A2(KEYINPUT10), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT10), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(new_n338), .B2(new_n340), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n309), .B(new_n336), .C1(new_n342), .C2(new_n344), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n271), .A2(new_n275), .B1(new_n279), .B2(G232), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n282), .A2(new_n283), .ZN(new_n347));
  OR2_X1    g0147(.A1(KEYINPUT72), .A2(G1698), .ZN(new_n348));
  NAND2_X1  g0148(.A1(KEYINPUT72), .A2(G1698), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(G223), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G226), .A2(G1698), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n347), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G87), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n263), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n320), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n346), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n356), .A2(new_n333), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(G190), .B2(new_n356), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n284), .A2(new_n288), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT7), .B1(new_n359), .B2(new_n207), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n286), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n287), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT79), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n347), .A2(KEYINPUT79), .A3(KEYINPUT7), .A4(new_n207), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(G68), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G58), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n367), .A2(new_n211), .ZN(new_n368));
  OAI21_X1  g0168(.A(G20), .B1(new_n368), .B2(new_n224), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n265), .A2(G159), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT16), .B1(new_n366), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT80), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(G20), .B1(new_n284), .B2(new_n288), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n363), .B(new_n364), .C1(new_n376), .C2(KEYINPUT7), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n371), .B1(new_n377), .B2(G68), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT80), .B1(new_n378), .B2(KEYINPUT16), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT7), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n286), .A2(new_n287), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n380), .B1(new_n381), .B2(G20), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n361), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n371), .B1(new_n383), .B2(G68), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n259), .B1(new_n384), .B2(KEYINPUT16), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n375), .A2(new_n379), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n262), .A2(KEYINPUT81), .A3(new_n256), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n254), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT81), .B1(new_n262), .B2(new_n256), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n388), .A2(new_n389), .B1(new_n250), .B2(new_n262), .ZN(new_n390));
  XNOR2_X1  g0190(.A(new_n390), .B(KEYINPUT82), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n358), .A2(new_n386), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT17), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n358), .A2(new_n386), .A3(KEYINPUT17), .A4(new_n391), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n385), .B1(new_n373), .B2(new_n374), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n378), .A2(KEYINPUT80), .A3(KEYINPUT16), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n391), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT83), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n346), .A2(new_n355), .A3(new_n308), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n400), .B(new_n401), .C1(new_n356), .C2(new_n303), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n346), .A2(new_n355), .A3(new_n308), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n303), .B1(new_n346), .B2(new_n355), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT83), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT18), .B1(new_n399), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n399), .A2(KEYINPUT18), .A3(new_n406), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n407), .B1(KEYINPUT84), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT84), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n399), .A2(new_n410), .A3(new_n406), .A4(KEYINPUT18), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n396), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n265), .A2(G50), .ZN(new_n414));
  XOR2_X1   g0214(.A(new_n414), .B(KEYINPUT78), .Z(new_n415));
  INV_X1    g0215(.A(new_n264), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n416), .A2(new_n294), .B1(new_n207), .B2(G68), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n253), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT11), .ZN(new_n419));
  OR2_X1    g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n419), .ZN(new_n421));
  OR3_X1    g0221(.A1(new_n250), .A2(KEYINPUT12), .A3(G68), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT12), .B1(new_n250), .B2(G68), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n255), .A2(new_n211), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n422), .A2(new_n423), .B1(new_n254), .B2(new_n424), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n420), .A2(new_n421), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT14), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT77), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n289), .A2(new_n429), .A3(G232), .A4(G1698), .ZN(new_n430));
  INV_X1    g0230(.A(G97), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n263), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n284), .A2(new_n288), .A3(G232), .A4(G1698), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT77), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n284), .A2(new_n288), .A3(G226), .A4(new_n292), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n430), .A2(new_n433), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n437), .A2(new_n320), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n279), .A2(G238), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n276), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT13), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n440), .B1(new_n437), .B2(new_n320), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT13), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n428), .B1(new_n445), .B2(G169), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n442), .A2(new_n443), .ZN(new_n447));
  AOI211_X1 g0247(.A(KEYINPUT13), .B(new_n440), .C1(new_n437), .C2(new_n320), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n428), .B(G169), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n441), .A2(G179), .A3(new_n444), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n427), .B1(new_n446), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n441), .A2(G190), .A3(new_n444), .ZN(new_n453));
  OAI21_X1  g0253(.A(G200), .B1(new_n447), .B2(new_n448), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n453), .A2(new_n454), .A3(new_n426), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n345), .A2(new_n413), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT87), .ZN(new_n459));
  AND2_X1   g0259(.A1(KEYINPUT4), .A2(G244), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n284), .A2(new_n288), .A3(new_n292), .A4(new_n460), .ZN(new_n461));
  XOR2_X1   g0261(.A(KEYINPUT85), .B(KEYINPUT4), .Z(new_n462));
  OAI21_X1  g0262(.A(G244), .B1(new_n282), .B2(new_n283), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n348), .A2(new_n349), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G283), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n461), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G250), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n297), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n320), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n206), .A2(G45), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT5), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(G41), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT86), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G41), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n474), .B1(new_n476), .B2(KEYINPUT5), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(KEYINPUT5), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n320), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT86), .B1(new_n472), .B2(G41), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(new_n473), .ZN(new_n482));
  INV_X1    g0282(.A(G45), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(G1), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(new_n478), .B2(KEYINPUT86), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g0286(.A1(G257), .A2(new_n480), .B1(new_n486), .B2(new_n275), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n470), .A2(new_n487), .A3(new_n307), .ZN(new_n488));
  OAI21_X1  g0288(.A(G107), .B1(new_n360), .B2(new_n365), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT6), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n490), .A2(new_n431), .A3(G107), .ZN(new_n491));
  XNOR2_X1  g0291(.A(G97), .B(G107), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n491), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n265), .ZN(new_n494));
  OAI22_X1  g0294(.A1(new_n493), .A2(new_n207), .B1(new_n294), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n259), .B1(new_n489), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n250), .A2(G97), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n206), .A2(G33), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n254), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n499), .B1(new_n501), .B2(new_n431), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n488), .B1(new_n497), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(G169), .B1(new_n470), .B2(new_n487), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n459), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n497), .A2(new_n502), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n470), .A2(new_n487), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G200), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n506), .B(new_n508), .C1(new_n331), .C2(new_n507), .ZN(new_n509));
  INV_X1    g0309(.A(new_n504), .ZN(new_n510));
  INV_X1    g0310(.A(new_n502), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n495), .B1(new_n377), .B2(G107), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n511), .B1(new_n512), .B2(new_n259), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n510), .A2(new_n513), .A3(KEYINPUT87), .A4(new_n488), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n505), .A2(new_n509), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n501), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT25), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n250), .B2(G107), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n251), .A2(KEYINPUT25), .A3(new_n323), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n516), .A2(G107), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n353), .A2(KEYINPUT22), .A3(G20), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n284), .A2(new_n288), .A3(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n207), .B(G87), .C1(new_n282), .C2(new_n283), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT22), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT90), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT23), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n527), .A2(new_n323), .A3(G20), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT89), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G116), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n527), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n207), .ZN(new_n533));
  NAND2_X1  g0333(.A1(KEYINPUT23), .A2(G107), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n527), .A2(new_n323), .A3(KEYINPUT89), .A4(G20), .ZN(new_n535));
  AND4_X1   g0335(.A1(new_n530), .A2(new_n533), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n525), .A2(new_n526), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n526), .B1(new_n525), .B2(new_n536), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT24), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n525), .A2(new_n536), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(KEYINPUT90), .A3(new_n539), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n253), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n520), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT91), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n530), .A2(new_n533), .A3(new_n534), .A4(new_n535), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n524), .B2(new_n522), .ZN(new_n547));
  OAI21_X1  g0347(.A(KEYINPUT24), .B1(new_n547), .B2(new_n526), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n253), .B(new_n542), .C1(new_n548), .C2(new_n537), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT91), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(new_n520), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n292), .A2(G250), .ZN(new_n552));
  NAND2_X1  g0352(.A1(G257), .A2(G1698), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n347), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(G294), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n263), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n320), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n475), .A2(new_n275), .A3(new_n479), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n480), .A2(G264), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G169), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n557), .A2(G179), .A3(new_n558), .A4(new_n559), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n545), .A2(new_n551), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n560), .A2(new_n333), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n557), .A2(new_n331), .A3(new_n558), .A4(new_n559), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(KEYINPUT92), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT92), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n560), .A2(new_n568), .A3(new_n333), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n567), .A2(new_n549), .A3(new_n520), .A4(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT19), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n416), .B2(new_n431), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n381), .A2(new_n207), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n353), .A2(new_n431), .A3(new_n323), .ZN(new_n574));
  XNOR2_X1  g0374(.A(new_n574), .B(KEYINPUT88), .ZN(new_n575));
  AOI21_X1  g0375(.A(G20), .B1(new_n432), .B2(KEYINPUT19), .ZN(new_n576));
  OAI221_X1 g0376(.A(new_n572), .B1(new_n211), .B2(new_n573), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n577), .A2(new_n253), .B1(new_n251), .B2(new_n314), .ZN(new_n578));
  OAI211_X1 g0378(.A(G244), .B(G1698), .C1(new_n282), .C2(new_n283), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n579), .A2(new_n531), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n381), .A2(new_n292), .A3(G238), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n278), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n275), .A2(new_n484), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n278), .A2(G250), .A3(new_n471), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(G200), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n516), .A2(G87), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n581), .A2(new_n531), .A3(new_n579), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n320), .ZN(new_n589));
  INV_X1    g0389(.A(new_n585), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(G190), .A3(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n578), .A2(new_n586), .A3(new_n587), .A4(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n575), .A2(new_n576), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n572), .B1(new_n573), .B2(new_n211), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n253), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n251), .A2(new_n314), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n595), .B(new_n596), .C1(new_n501), .C2(new_n314), .ZN(new_n597));
  OAI21_X1  g0397(.A(G169), .B1(new_n582), .B2(new_n585), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n589), .A2(new_n308), .A3(new_n590), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n592), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n359), .A2(G303), .ZN(new_n603));
  INV_X1    g0403(.A(G257), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n290), .A2(new_n291), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G264), .A2(G1698), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n381), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n278), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(G270), .B(new_n278), .C1(new_n482), .C2(new_n485), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n558), .ZN(new_n611));
  OAI21_X1  g0411(.A(G200), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g0412(.A1(G270), .A2(new_n480), .B1(new_n486), .B2(new_n275), .ZN(new_n613));
  INV_X1    g0413(.A(G303), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n284), .B2(new_n288), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n348), .A2(G257), .A3(new_n349), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n347), .B1(new_n616), .B2(new_n606), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n320), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n613), .A2(G190), .A3(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(G116), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n251), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n259), .A2(new_n250), .A3(G116), .A4(new_n500), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n252), .A2(new_n222), .B1(G20), .B2(new_n620), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n466), .B(new_n207), .C1(G33), .C2(new_n431), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n623), .A2(KEYINPUT20), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT20), .B1(new_n623), .B2(new_n624), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n621), .B(new_n622), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n612), .A2(new_n619), .A3(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(G169), .B(new_n627), .C1(new_n609), .C2(new_n611), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT21), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n613), .A2(new_n627), .A3(G179), .A4(new_n618), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n613), .A2(new_n618), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n634), .A2(KEYINPUT21), .A3(G169), .A4(new_n627), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n629), .A2(new_n632), .A3(new_n633), .A4(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n602), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n515), .A2(new_n564), .A3(new_n570), .A4(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n458), .A2(new_n638), .ZN(G372));
  XNOR2_X1  g0439(.A(new_n341), .B(KEYINPUT10), .ZN(new_n640));
  OAI21_X1  g0440(.A(G169), .B1(new_n447), .B2(new_n448), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT14), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n642), .A2(new_n450), .A3(new_n449), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n643), .A2(new_n427), .B1(new_n455), .B2(new_n330), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n644), .A2(new_n396), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n399), .A2(KEYINPUT18), .A3(new_n406), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(new_n407), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n640), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n648), .A2(new_n309), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n600), .A2(KEYINPUT93), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT93), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n651), .B1(new_n598), .B2(new_n599), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n597), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n503), .A2(new_n504), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n653), .A2(new_n654), .A3(new_n655), .A4(new_n592), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n602), .B1(new_n505), .B2(new_n514), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n653), .B(new_n656), .C1(new_n657), .C2(new_n655), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n570), .A2(new_n653), .A3(new_n592), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(new_n515), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT94), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n549), .A2(new_n520), .B1(new_n561), .B2(new_n562), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n544), .A2(new_n563), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n633), .B1(new_n630), .B2(new_n631), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n303), .B1(new_n613), .B2(new_n618), .ZN(new_n667));
  AOI21_X1  g0467(.A(KEYINPUT21), .B1(new_n667), .B2(new_n627), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n665), .A2(KEYINPUT94), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n664), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n658), .B1(new_n660), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n649), .B1(new_n458), .B2(new_n672), .ZN(G369));
  AND2_X1   g0473(.A1(new_n564), .A2(new_n570), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n249), .A2(new_n675), .A3(new_n207), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n676), .A2(new_n678), .A3(G213), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT95), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n676), .A2(new_n678), .A3(KEYINPUT95), .A4(G213), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT96), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(G343), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(G343), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n683), .A2(KEYINPUT97), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n681), .A2(new_n682), .A3(new_n687), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT97), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n545), .A2(new_n551), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n674), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n692), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n564), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n628), .B1(new_n688), .B2(new_n691), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n666), .B2(new_n668), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n636), .B2(new_n698), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT98), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT98), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n699), .B(new_n702), .C1(new_n636), .C2(new_n698), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n701), .A2(KEYINPUT99), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT99), .B1(new_n701), .B2(new_n703), .ZN(new_n705));
  OAI21_X1  g0505(.A(G330), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n706), .A2(KEYINPUT100), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT100), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n708), .B(G330), .C1(new_n704), .C2(new_n705), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n697), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n669), .A2(new_n692), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n564), .A2(new_n570), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n662), .A2(new_n695), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT101), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n713), .A2(KEYINPUT101), .A3(new_n714), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n711), .A2(new_n719), .ZN(G399));
  INV_X1    g0520(.A(new_n227), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G41), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n575), .A2(new_n620), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n723), .A2(G1), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n225), .A2(G50), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n726), .B1(new_n727), .B2(new_n723), .ZN(new_n728));
  XOR2_X1   g0528(.A(new_n728), .B(KEYINPUT28), .Z(new_n729));
  NAND4_X1  g0529(.A1(new_n557), .A2(new_n559), .A3(new_n589), .A4(new_n590), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n613), .A2(G179), .A3(new_n618), .ZN(new_n731));
  OR3_X1    g0531(.A1(new_n507), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n308), .B1(new_n589), .B2(new_n590), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n507), .A2(new_n560), .A3(new_n634), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n732), .A2(new_n733), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n692), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT31), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n564), .A2(new_n570), .A3(new_n637), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n505), .A2(new_n509), .A3(new_n514), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(KEYINPUT102), .B1(new_n743), .B2(new_n695), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT102), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n638), .A2(new_n745), .A3(new_n692), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n740), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT29), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(new_n672), .B2(new_n692), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n657), .A2(new_n655), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n653), .A2(new_n592), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n751), .A2(new_n504), .A3(new_n503), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n750), .B(new_n653), .C1(new_n752), .C2(new_n655), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n564), .A2(new_n669), .ZN(new_n754));
  AND3_X1   g0554(.A1(new_n754), .A2(new_n659), .A3(new_n515), .ZN(new_n755));
  OAI211_X1 g0555(.A(KEYINPUT29), .B(new_n695), .C1(new_n753), .C2(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(G330), .A2(new_n747), .B1(new_n749), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n729), .B1(new_n758), .B2(new_n206), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT103), .ZN(G364));
  NOR2_X1   g0560(.A1(new_n248), .A2(G20), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n206), .B1(new_n761), .B2(G45), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n722), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n701), .A2(new_n703), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n222), .B1(G20), .B2(new_n303), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n207), .A2(new_n333), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n308), .A2(G190), .A3(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n207), .A2(G190), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n308), .A2(new_n333), .A3(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(G326), .A2(new_n772), .B1(new_n775), .B2(G311), .ZN(new_n776));
  INV_X1    g0576(.A(G322), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n207), .A2(new_n331), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n308), .A2(new_n333), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n308), .A2(new_n331), .A3(new_n770), .ZN(new_n780));
  XOR2_X1   g0580(.A(KEYINPUT33), .B(G317), .Z(new_n781));
  OAI221_X1 g0581(.A(new_n776), .B1(new_n777), .B2(new_n779), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n333), .A2(G179), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G179), .A2(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n773), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G303), .A2(new_n785), .B1(new_n788), .B2(G329), .ZN(new_n789));
  INV_X1    g0589(.A(G283), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n773), .A2(new_n783), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n786), .A2(G190), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G20), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n359), .B1(new_n795), .B2(new_n555), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n782), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n780), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G50), .A2(new_n772), .B1(new_n798), .B2(G68), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n367), .B2(new_n779), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT104), .B(G159), .ZN(new_n801));
  OR3_X1    g0601(.A1(new_n787), .A2(new_n801), .A3(KEYINPUT32), .ZN(new_n802));
  OAI21_X1  g0602(.A(KEYINPUT32), .B1(new_n787), .B2(new_n801), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n794), .A2(G97), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n774), .A2(new_n294), .ZN(new_n806));
  INV_X1    g0606(.A(new_n791), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G107), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n808), .B(new_n289), .C1(new_n353), .C2(new_n784), .ZN(new_n809));
  NOR4_X1   g0609(.A1(new_n800), .A2(new_n805), .A3(new_n806), .A4(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n769), .B1(new_n797), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n767), .A2(new_n769), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n721), .A2(new_n381), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(G45), .B2(new_n727), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G45), .B2(new_n246), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n289), .A2(new_n227), .ZN(new_n816));
  INV_X1    g0616(.A(G355), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n816), .A2(new_n817), .B1(G116), .B2(new_n227), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n812), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  AND4_X1   g0619(.A1(new_n764), .A2(new_n768), .A3(new_n811), .A4(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n707), .A2(new_n710), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n704), .A2(new_n705), .ZN(new_n822));
  INV_X1    g0622(.A(G330), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n764), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n820), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G396));
  INV_X1    g0626(.A(new_n658), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n671), .A2(new_n515), .A3(new_n659), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n692), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n328), .A2(new_n329), .ZN(new_n830));
  INV_X1    g0630(.A(new_n319), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n692), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(KEYINPUT105), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT105), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n831), .A2(new_n692), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n830), .B1(new_n335), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n330), .A2(new_n695), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n829), .B(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n743), .A2(KEYINPUT102), .A3(new_n695), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n745), .B1(new_n638), .B2(new_n692), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n823), .B1(new_n844), .B2(new_n740), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n764), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n841), .A2(new_n845), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT106), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n791), .A2(new_n211), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(G132), .B2(new_n788), .ZN(new_n852));
  INV_X1    g0652(.A(G50), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n852), .B(new_n381), .C1(new_n853), .C2(new_n784), .ZN(new_n854));
  INV_X1    g0654(.A(new_n779), .ZN(new_n855));
  INV_X1    g0655(.A(new_n801), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G143), .A2(new_n855), .B1(new_n775), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(G137), .ZN(new_n858));
  INV_X1    g0658(.A(G150), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n857), .B1(new_n858), .B2(new_n771), .C1(new_n859), .C2(new_n780), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT34), .Z(new_n861));
  AOI211_X1 g0661(.A(new_n854), .B(new_n861), .C1(G58), .C2(new_n794), .ZN(new_n862));
  AOI22_X1  g0662(.A1(G107), .A2(new_n785), .B1(new_n788), .B2(G311), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n807), .A2(G87), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n863), .A2(new_n359), .A3(new_n804), .A4(new_n864), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n555), .A2(new_n779), .B1(new_n771), .B2(new_n614), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n620), .A2(new_n774), .B1(new_n780), .B2(new_n790), .ZN(new_n867));
  NOR3_X1   g0667(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n769), .B1(new_n862), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n769), .A2(new_n765), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n869), .B1(G77), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n840), .A2(new_n766), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n764), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n849), .A2(new_n850), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n850), .B1(new_n849), .B2(new_n874), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n875), .A2(new_n876), .ZN(G384));
  INV_X1    g0677(.A(new_n493), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n878), .A2(KEYINPUT35), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(KEYINPUT35), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n879), .A2(G116), .A3(new_n223), .A4(new_n880), .ZN(new_n881));
  XNOR2_X1  g0681(.A(KEYINPUT107), .B(KEYINPUT36), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n881), .B(new_n882), .ZN(new_n883));
  OR3_X1    g0683(.A1(new_n727), .A2(new_n294), .A3(new_n368), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n853), .A2(G68), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n206), .B(G13), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT39), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n385), .B1(KEYINPUT16), .B2(new_n384), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n391), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n683), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n408), .A2(KEYINPUT84), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n399), .A2(new_n406), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT18), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n892), .A2(new_n411), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n396), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n891), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n406), .A2(new_n890), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n392), .A2(new_n899), .A3(new_n891), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(KEYINPUT37), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n399), .A2(new_n683), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT37), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n893), .A2(new_n902), .A3(new_n903), .A4(new_n392), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT38), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n898), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n902), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n647), .B2(new_n396), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n893), .A2(new_n902), .A3(new_n392), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT37), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n904), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT38), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n888), .B1(new_n908), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n643), .A2(new_n427), .A3(new_n695), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n907), .B1(new_n898), .B2(new_n906), .ZN(new_n918));
  OAI211_X1 g0718(.A(KEYINPUT38), .B(new_n905), .C1(new_n412), .C2(new_n891), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n918), .A2(new_n919), .A3(KEYINPUT39), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n915), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n427), .A2(new_n692), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n452), .A2(new_n455), .A3(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n455), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n427), .B(new_n692), .C1(new_n643), .C2(new_n924), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n828), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n840), .B(new_n695), .C1(new_n927), .C2(new_n658), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n926), .B1(new_n928), .B2(new_n838), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n918), .A2(new_n919), .ZN(new_n930));
  INV_X1    g0730(.A(new_n683), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n929), .A2(new_n930), .B1(new_n647), .B2(new_n931), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n921), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n457), .A2(new_n749), .A3(new_n756), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n649), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n933), .B(new_n935), .Z(new_n936));
  INV_X1    g0736(.A(KEYINPUT31), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(KEYINPUT108), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n739), .A2(new_n938), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n739), .A2(new_n938), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n842), .A2(new_n843), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n923), .A2(new_n925), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n840), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT40), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n941), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n910), .A2(new_n913), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n907), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n919), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n941), .A2(new_n943), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT40), .B1(new_n951), .B2(new_n930), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n950), .A2(new_n952), .B1(new_n458), .B2(new_n941), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n930), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n944), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n940), .A2(new_n939), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n844), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n955), .A2(new_n457), .A3(new_n957), .A4(new_n949), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n953), .A2(G330), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n936), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n206), .B2(new_n761), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n936), .A2(new_n959), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n887), .B1(new_n961), .B2(new_n962), .ZN(G367));
  INV_X1    g0763(.A(KEYINPUT113), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT45), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT111), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n515), .B1(new_n506), .B2(new_n695), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n654), .A2(new_n692), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n966), .B1(new_n719), .B2(new_n969), .ZN(new_n970));
  AND3_X1   g0770(.A1(new_n713), .A2(KEYINPUT101), .A3(new_n714), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT101), .B1(new_n713), .B2(new_n714), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n966), .B(new_n969), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n965), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(KEYINPUT111), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n977), .A2(KEYINPUT45), .A3(new_n973), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n971), .A2(new_n972), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n979), .A2(KEYINPUT44), .A3(new_n967), .A4(new_n968), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT44), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n719), .B2(new_n969), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n975), .A2(new_n978), .A3(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n711), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n706), .A2(KEYINPUT100), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n987), .A2(KEYINPUT112), .A3(new_n709), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n713), .B1(new_n697), .B2(new_n712), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n987), .A2(new_n989), .A3(KEYINPUT112), .A4(new_n709), .ZN(new_n992));
  AND3_X1   g0792(.A1(new_n991), .A2(new_n757), .A3(new_n992), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n711), .A2(new_n975), .A3(new_n978), .A4(new_n983), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n986), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n757), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n722), .B(KEYINPUT41), .Z(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n964), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  AOI211_X1 g0799(.A(KEYINPUT113), .B(new_n997), .C1(new_n995), .C2(new_n757), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n762), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n578), .A2(new_n587), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n692), .ZN(new_n1003));
  MUX2_X1   g0803(.A(new_n653), .B(new_n751), .S(new_n1003), .Z(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT109), .ZN(new_n1005));
  AOI21_X1  g0805(.A(KEYINPUT43), .B1(new_n1005), .B2(KEYINPUT110), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(KEYINPUT110), .B2(new_n1005), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n713), .B1(new_n967), .B2(new_n968), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT42), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n564), .B1(new_n967), .B2(new_n968), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n505), .A2(new_n514), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n695), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1005), .A2(KEYINPUT43), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1007), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n1013), .B2(new_n1007), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n985), .A2(new_n969), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1016), .B(new_n1017), .Z(new_n1018));
  NAND2_X1  g0818(.A1(new_n1001), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n807), .A2(G77), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n367), .B2(new_n784), .C1(new_n858), .C2(new_n787), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n795), .A2(new_n211), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n1021), .A2(new_n359), .A3(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G150), .A2(new_n855), .B1(new_n798), .B2(new_n856), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G143), .A2(new_n772), .B1(new_n775), .B2(G50), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT114), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n807), .A2(G97), .ZN(new_n1029));
  INV_X1    g0829(.A(G317), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1029), .B(new_n347), .C1(new_n1030), .C2(new_n787), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n785), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT46), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n784), .B2(new_n620), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1032), .B(new_n1034), .C1(new_n323), .C2(new_n795), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n1031), .B(new_n1035), .C1(G303), .C2(new_n855), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G294), .A2(new_n798), .B1(new_n775), .B2(G283), .ZN(new_n1037));
  INV_X1    g0837(.A(G311), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1036), .B(new_n1037), .C1(new_n1038), .C2(new_n771), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1028), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  XOR2_X1   g0841(.A(KEYINPUT115), .B(KEYINPUT47), .Z(new_n1042));
  XNOR2_X1  g0842(.A(new_n1041), .B(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n769), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n812), .B1(new_n227), .B2(new_n314), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n813), .B2(new_n234), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n847), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n767), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1044), .B(new_n1047), .C1(new_n1005), .C2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1019), .A2(new_n1049), .ZN(G387));
  NAND3_X1  g0850(.A1(new_n991), .A2(new_n763), .A3(new_n992), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n813), .B1(new_n239), .B2(new_n483), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n725), .B2(new_n816), .ZN(new_n1053));
  OR3_X1    g0853(.A1(new_n261), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1054));
  OAI21_X1  g0854(.A(KEYINPUT50), .B1(new_n261), .B2(G50), .ZN(new_n1055));
  AOI21_X1  g0855(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n725), .A2(new_n1054), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1053), .A2(new_n1057), .B1(new_n323), .B2(new_n721), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n812), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n764), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n211), .A2(new_n774), .B1(new_n780), .B2(new_n261), .ZN(new_n1061));
  INV_X1    g0861(.A(G159), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n853), .A2(new_n779), .B1(new_n771), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n785), .A2(G77), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n788), .A2(G150), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1064), .A2(new_n1029), .A3(new_n1065), .A4(new_n381), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n795), .A2(new_n314), .ZN(new_n1067));
  NOR4_X1   g0867(.A1(new_n1061), .A2(new_n1063), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT116), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n381), .B1(new_n788), .B2(G326), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n795), .A2(new_n790), .B1(new_n784), .B2(new_n555), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT117), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G311), .A2(new_n798), .B1(new_n772), .B2(G322), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n614), .B2(new_n774), .C1(new_n1030), .C2(new_n779), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT48), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1072), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n1075), .B2(new_n1074), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT49), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1070), .B1(new_n620), .B2(new_n791), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1069), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1060), .B1(new_n1081), .B2(new_n769), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n697), .B2(new_n1048), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n993), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n722), .B(KEYINPUT118), .Z(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n757), .B1(new_n991), .B2(new_n992), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1051), .B(new_n1083), .C1(new_n1086), .C2(new_n1087), .ZN(G393));
  NAND3_X1  g0888(.A1(new_n986), .A2(new_n763), .A3(new_n994), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n969), .A2(new_n1048), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT119), .Z(new_n1091));
  OAI21_X1  g0891(.A(new_n812), .B1(new_n431), .B2(new_n227), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n813), .B2(new_n243), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n798), .A2(G303), .B1(G116), .B2(new_n794), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n555), .B2(new_n774), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT122), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n1038), .A2(new_n779), .B1(new_n771), .B2(new_n1030), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT52), .Z(new_n1098));
  OAI221_X1 g0898(.A(new_n808), .B1(new_n790), .B2(new_n784), .C1(new_n777), .C2(new_n787), .ZN(new_n1099));
  OR4_X1    g0899(.A1(new_n289), .A2(new_n1096), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n859), .A2(new_n771), .B1(new_n779), .B2(new_n1062), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(KEYINPUT120), .B(KEYINPUT51), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1101), .B(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n795), .A2(new_n294), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G68), .A2(new_n785), .B1(new_n788), .B2(G143), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1105), .A2(new_n381), .A3(new_n864), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n853), .A2(new_n780), .B1(new_n774), .B2(new_n261), .ZN(new_n1107));
  NOR4_X1   g0907(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1109), .A2(KEYINPUT121), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(KEYINPUT121), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1100), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n847), .B(new_n1093), .C1(new_n1112), .C2(new_n769), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1091), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1089), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT123), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1089), .A2(KEYINPUT123), .A3(new_n1114), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n995), .A2(new_n1085), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n986), .A2(new_n994), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n1084), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1117), .A2(new_n1118), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(G390));
  INV_X1    g0923(.A(new_n838), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n829), .B2(new_n840), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n916), .B1(new_n1125), .B2(new_n926), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n918), .A2(new_n919), .A3(KEYINPUT39), .ZN(new_n1127));
  AOI21_X1  g0927(.A(KEYINPUT39), .B1(new_n947), .B2(new_n919), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n695), .B(new_n837), .C1(new_n753), .C2(new_n755), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1130), .A2(new_n838), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n948), .B(new_n916), .C1(new_n1131), .C2(new_n926), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n845), .A2(new_n840), .A3(new_n942), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1129), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n941), .A2(new_n823), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n839), .B1(new_n923), .B2(new_n925), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n763), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n765), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n847), .B1(new_n261), .B2(new_n870), .ZN(new_n1142));
  INV_X1    g0942(.A(G125), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n791), .A2(new_n853), .B1(new_n787), .B2(new_n1143), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n359), .B(new_n1144), .C1(G159), .C2(new_n794), .ZN(new_n1145));
  XOR2_X1   g0945(.A(KEYINPUT54), .B(G143), .Z(new_n1146));
  AOI22_X1  g0946(.A1(G128), .A2(new_n772), .B1(new_n775), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n798), .A2(G137), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n785), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT53), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n784), .B2(new_n859), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n855), .A2(G132), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1145), .A2(new_n1147), .A3(new_n1148), .A4(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(G107), .A2(new_n798), .B1(new_n855), .B2(G116), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(G283), .A2(new_n772), .B1(new_n775), .B2(G97), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n787), .A2(new_n555), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1156), .B(new_n851), .C1(G87), .C2(new_n785), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1104), .A2(new_n289), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1154), .A2(new_n1155), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1153), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1160), .A2(KEYINPUT124), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(KEYINPUT124), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n769), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1141), .B(new_n1142), .C1(new_n1161), .C2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n957), .A2(G330), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n926), .B1(new_n1165), .B2(new_n839), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1166), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1125), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1165), .A2(new_n943), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n942), .B1(new_n845), .B2(new_n840), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1168), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1167), .A2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n934), .B(new_n649), .C1(new_n458), .C2(new_n1165), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n692), .B(new_n839), .C1(new_n827), .C2(new_n828), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n942), .B1(new_n1176), .B2(new_n1124), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n915), .A2(new_n920), .B1(new_n1177), .B2(new_n916), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n898), .A2(new_n906), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n914), .B1(new_n1179), .B2(KEYINPUT38), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n926), .B1(new_n1130), .B2(new_n838), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1180), .A2(new_n1181), .A3(new_n917), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1169), .B1(new_n1178), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1129), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1085), .B1(new_n1175), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1173), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1139), .A2(new_n1187), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1140), .B(new_n1164), .C1(new_n1186), .C2(new_n1188), .ZN(G378));
  AOI21_X1  g0989(.A(new_n823), .B1(new_n945), .B2(new_n948), .ZN(new_n1190));
  XOR2_X1   g0990(.A(KEYINPUT125), .B(KEYINPUT56), .Z(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n268), .A2(new_n931), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT55), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n640), .B2(new_n309), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n309), .B(new_n1195), .C1(new_n342), .C2(new_n344), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1192), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n309), .B1(new_n342), .B2(new_n344), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n1194), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1201), .A2(new_n1191), .A3(new_n1197), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1190), .A2(new_n955), .A3(new_n1203), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n957), .A2(KEYINPUT40), .A3(new_n1136), .ZN(new_n1206));
  OAI21_X1  g1006(.A(G330), .B1(new_n1206), .B2(new_n1180), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1205), .B1(new_n1207), .B2(new_n952), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1204), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n933), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1204), .A2(new_n933), .A3(new_n1208), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1205), .A2(new_n765), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n871), .A2(G50), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n263), .B(new_n476), .C1(new_n791), .C2(new_n801), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n785), .A2(new_n1146), .B1(new_n794), .B2(G150), .ZN(new_n1217));
  INV_X1    g1017(.A(G132), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1217), .B1(new_n1218), .B2(new_n780), .ZN(new_n1219));
  INV_X1    g1019(.A(G128), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n1143), .A2(new_n771), .B1(new_n779), .B2(new_n1220), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1219), .B(new_n1221), .C1(G137), .C2(new_n775), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1216), .B(new_n1224), .C1(G124), .C2(new_n788), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(KEYINPUT59), .B2(new_n1223), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1064), .B1(new_n790), .B2(new_n787), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n347), .A2(new_n476), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n791), .A2(new_n367), .ZN(new_n1229));
  NOR4_X1   g1029(.A1(new_n1227), .A2(new_n1022), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(G116), .A2(new_n772), .B1(new_n775), .B2(new_n315), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(G97), .A2(new_n798), .B1(new_n855), .B2(G107), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT58), .ZN(new_n1234));
  AOI21_X1  g1034(.A(G50), .B1(new_n263), .B2(new_n476), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1233), .A2(new_n1234), .B1(new_n1228), .B2(new_n1235), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1226), .B(new_n1236), .C1(new_n1234), .C2(new_n1233), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n847), .B(new_n1215), .C1(new_n1237), .C2(new_n769), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1213), .A2(new_n763), .B1(new_n1214), .B2(new_n1238), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1204), .A2(new_n933), .A3(new_n1208), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n933), .B1(new_n1204), .B2(new_n1208), .ZN(new_n1241));
  OAI21_X1  g1041(.A(KEYINPUT57), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1173), .B1(new_n1139), .B2(new_n1172), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1085), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1174), .B1(new_n1175), .B2(new_n1185), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT57), .B1(new_n1213), .B2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1239), .B1(new_n1244), .B2(new_n1246), .ZN(G375));
  NAND3_X1  g1047(.A1(new_n1167), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1175), .A2(new_n998), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n926), .A2(new_n765), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n764), .B1(G68), .B2(new_n871), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(G283), .A2(new_n855), .B1(new_n772), .B2(G294), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n1252), .B1(new_n323), .B2(new_n774), .C1(new_n620), .C2(new_n780), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1020), .B1(new_n431), .B2(new_n784), .C1(new_n614), .C2(new_n787), .ZN(new_n1254));
  NOR4_X1   g1054(.A1(new_n1253), .A2(new_n289), .A3(new_n1067), .A4(new_n1254), .ZN(new_n1255));
  OR2_X1    g1055(.A1(new_n1255), .A2(KEYINPUT126), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(KEYINPUT126), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(G132), .A2(new_n772), .B1(new_n855), .B2(G137), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n798), .A2(new_n1146), .B1(new_n775), .B2(G150), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n795), .A2(new_n853), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n784), .A2(new_n1062), .B1(new_n787), .B2(new_n1220), .ZN(new_n1261));
  NOR4_X1   g1061(.A1(new_n1260), .A2(new_n1261), .A3(new_n347), .A4(new_n1229), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1258), .A2(new_n1259), .A3(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1256), .A2(new_n1257), .A3(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1251), .B1(new_n1264), .B2(new_n769), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n1172), .A2(new_n763), .B1(new_n1250), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1249), .A2(new_n1266), .ZN(G381));
  NOR2_X1   g1067(.A1(G393), .A2(G396), .ZN(new_n1268));
  INV_X1    g1068(.A(G384), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NOR4_X1   g1070(.A1(G390), .A2(new_n1270), .A3(G378), .A4(G381), .ZN(new_n1271));
  INV_X1    g1071(.A(G375), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1271), .A2(new_n1019), .A3(new_n1049), .A4(new_n1272), .ZN(G407));
  OAI21_X1  g1073(.A(new_n1164), .B1(new_n1185), .B2(new_n762), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1085), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(new_n1139), .B2(new_n1187), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1175), .A2(new_n1185), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1274), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n685), .A2(new_n686), .A3(G213), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1272), .A2(new_n1278), .A3(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(G407), .A2(G213), .A3(new_n1281), .ZN(G409));
  INV_X1    g1082(.A(KEYINPUT127), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G390), .B1(new_n1019), .B2(new_n1049), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1049), .ZN(new_n1285));
  AOI211_X1 g1085(.A(new_n1285), .B(new_n1122), .C1(new_n1001), .C2(new_n1018), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1283), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(G393), .A2(G396), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1289), .A2(new_n1268), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1287), .A2(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1287), .A2(new_n1290), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  OAI211_X1 g1093(.A(G378), .B(new_n1239), .C1(new_n1244), .C2(new_n1246), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1213), .A2(new_n1245), .A3(new_n998), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1214), .A2(new_n1238), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1296), .B1(new_n1297), .B2(new_n762), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1278), .B1(new_n1295), .B2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1280), .B1(new_n1294), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT60), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1248), .A2(new_n1301), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1167), .A2(new_n1171), .A3(KEYINPUT60), .A4(new_n1173), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1302), .A2(new_n1175), .A3(new_n1085), .A4(new_n1303), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1304), .A2(G384), .A3(new_n1266), .ZN(new_n1305));
  AOI21_X1  g1105(.A(G384), .B1(new_n1304), .B2(new_n1266), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1300), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT61), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1300), .A2(KEYINPUT63), .A3(new_n1307), .ZN(new_n1312));
  OAI211_X1 g1112(.A(G2897), .B(new_n1280), .C1(new_n1305), .C2(new_n1306), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1306), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1304), .A2(G384), .A3(new_n1266), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1280), .A2(G2897), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1314), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  AND2_X1   g1117(.A1(new_n1313), .A2(new_n1317), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1294), .A2(new_n1299), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1318), .B1(new_n1319), .B2(new_n1280), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1310), .A2(new_n1311), .A3(new_n1312), .A4(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1313), .A2(new_n1317), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1311), .B1(new_n1300), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1287), .A2(new_n1290), .ZN(new_n1324));
  OAI221_X1 g1124(.A(new_n1283), .B1(new_n1268), .B2(new_n1289), .C1(new_n1284), .C2(new_n1286), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1323), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT62), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1308), .A2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1300), .A2(KEYINPUT62), .A3(new_n1307), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  AOI22_X1  g1130(.A1(new_n1293), .A2(new_n1321), .B1(new_n1326), .B2(new_n1330), .ZN(G405));
  NAND2_X1  g1131(.A1(G375), .A2(new_n1278), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1294), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1307), .ZN(new_n1334));
  OAI211_X1 g1134(.A(new_n1332), .B(new_n1294), .C1(new_n1306), .C2(new_n1305), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1336), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1324), .A2(new_n1325), .A3(new_n1334), .A4(new_n1335), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(G402));
endmodule


