//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 1 0 1 1 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n187));
  OR2_X1    g001(.A1(G475), .A2(G902), .ZN(new_n188));
  INV_X1    g002(.A(G131), .ZN(new_n189));
  INV_X1    g003(.A(G214), .ZN(new_n190));
  NOR3_X1   g004(.A1(new_n190), .A2(G237), .A3(G953), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT64), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT81), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n191), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(G237), .A2(G953), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT64), .A2(KEYINPUT81), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n199), .A2(new_n192), .A3(new_n200), .A4(G214), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n189), .B1(new_n198), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT17), .ZN(new_n204));
  AOI21_X1  g018(.A(KEYINPUT81), .B1(new_n193), .B2(new_n195), .ZN(new_n205));
  OAI211_X1 g019(.A(G131), .B(new_n201), .C1(new_n205), .C2(new_n191), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n206), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT17), .ZN(new_n209));
  INV_X1    g023(.A(G125), .ZN(new_n210));
  NOR3_X1   g024(.A1(new_n210), .A2(KEYINPUT16), .A3(G140), .ZN(new_n211));
  INV_X1    g025(.A(G140), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(G125), .A2(G140), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n211), .B1(new_n215), .B2(KEYINPUT16), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(G146), .ZN(new_n217));
  AND2_X1   g031(.A1(G125), .A2(G140), .ZN(new_n218));
  NOR2_X1   g032(.A1(G125), .A2(G140), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT16), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  OR3_X1    g034(.A1(new_n210), .A2(KEYINPUT16), .A3(G140), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(G146), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n207), .A2(new_n209), .A3(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G113), .B(G122), .ZN(new_n226));
  INV_X1    g040(.A(G104), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n226), .B(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT18), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n198), .B2(new_n202), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n199), .A2(G214), .ZN(new_n231));
  XNOR2_X1  g045(.A(KEYINPUT64), .B(G143), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(KEYINPUT81), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n233), .A2(KEYINPUT18), .A3(G131), .A4(new_n201), .ZN(new_n234));
  INV_X1    g048(.A(G146), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n215), .B(new_n235), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n230), .A2(new_n203), .A3(new_n234), .A4(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n225), .A2(new_n228), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT83), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT83), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n225), .A2(new_n240), .A3(new_n228), .A4(new_n237), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT19), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n243), .B1(new_n218), .B2(new_n219), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n213), .A2(KEYINPUT19), .A3(new_n214), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n245), .A3(new_n235), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n246), .A2(new_n222), .ZN(new_n247));
  AOI21_X1  g061(.A(G131), .B1(new_n233), .B2(new_n201), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n247), .B1(new_n208), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n237), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n228), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT82), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT82), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n250), .A2(new_n254), .A3(new_n251), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n188), .B1(new_n242), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT20), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n187), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n241), .A2(new_n239), .B1(new_n253), .B2(new_n255), .ZN(new_n260));
  OAI211_X1 g074(.A(KEYINPUT84), .B(KEYINPUT20), .C1(new_n260), .C2(new_n188), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n257), .A2(new_n258), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G902), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n228), .B1(new_n225), .B2(new_n237), .ZN(new_n265));
  XOR2_X1   g079(.A(new_n265), .B(KEYINPUT85), .Z(new_n266));
  INV_X1    g080(.A(new_n242), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n264), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G475), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n263), .A2(KEYINPUT86), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT86), .B1(new_n263), .B2(new_n269), .ZN(new_n271));
  XOR2_X1   g085(.A(KEYINPUT9), .B(G234), .Z(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G217), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n273), .A2(new_n274), .A3(G953), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n196), .A2(G128), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n277), .B1(G128), .B2(new_n192), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(G134), .ZN(new_n279));
  XNOR2_X1  g093(.A(G116), .B(G122), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n280), .B(G107), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT13), .B1(new_n192), .B2(G128), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n283), .B(KEYINPUT87), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n196), .A2(KEYINPUT13), .A3(G128), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n285), .B(KEYINPUT88), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  AOI211_X1 g101(.A(new_n279), .B(new_n281), .C1(new_n287), .C2(G134), .ZN(new_n288));
  INV_X1    g102(.A(G116), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT14), .A3(G122), .ZN(new_n290));
  INV_X1    g104(.A(new_n280), .ZN(new_n291));
  OAI211_X1 g105(.A(G107), .B(new_n290), .C1(new_n291), .C2(KEYINPUT14), .ZN(new_n292));
  XOR2_X1   g106(.A(new_n292), .B(KEYINPUT89), .Z(new_n293));
  INV_X1    g107(.A(G107), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n280), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G134), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n278), .B(new_n297), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n293), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n276), .B1(new_n288), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n287), .A2(G134), .ZN(new_n301));
  INV_X1    g115(.A(new_n279), .ZN(new_n302));
  INV_X1    g116(.A(new_n281), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n299), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(new_n275), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT91), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n308), .A3(new_n264), .ZN(new_n309));
  INV_X1    g123(.A(G478), .ZN(new_n310));
  NOR2_X1   g124(.A1(KEYINPUT90), .A2(KEYINPUT15), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(KEYINPUT90), .A2(KEYINPUT15), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n310), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(G902), .B1(new_n300), .B2(new_n306), .ZN(new_n316));
  INV_X1    g130(.A(new_n314), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n308), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G953), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G952), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n321), .B1(G234), .B2(G237), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  XOR2_X1   g137(.A(KEYINPUT21), .B(G898), .Z(new_n324));
  NAND2_X1  g138(.A1(G234), .A2(G237), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(G902), .A3(G953), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n323), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NOR4_X1   g142(.A1(new_n270), .A2(new_n271), .A3(new_n319), .A4(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G472), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT11), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n297), .B2(G137), .ZN(new_n332));
  INV_X1    g146(.A(G137), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(KEYINPUT11), .A3(G134), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n297), .A2(G137), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n332), .A2(new_n334), .A3(new_n189), .A4(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n333), .A2(G134), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n297), .A2(G137), .ZN(new_n338));
  OAI21_X1  g152(.A(G131), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n235), .B1(new_n193), .B2(new_n195), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT66), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n342), .B1(new_n192), .B2(G146), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n235), .A2(KEYINPUT66), .A3(G143), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G128), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(KEYINPUT1), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n341), .A2(new_n345), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT65), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n350), .B1(new_n235), .B2(G143), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n192), .A2(KEYINPUT65), .A3(G146), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n193), .A2(new_n195), .A3(new_n235), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n353), .A2(new_n354), .B1(G128), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n340), .B1(new_n349), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n332), .A2(new_n335), .A3(new_n334), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G131), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n336), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n196), .A2(G146), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n343), .A2(new_n344), .ZN(new_n362));
  AND2_X1   g176(.A1(KEYINPUT0), .A2(G128), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n353), .A2(new_n354), .ZN(new_n365));
  NOR2_X1   g179(.A1(KEYINPUT0), .A2(G128), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n360), .A2(new_n364), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n357), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT67), .ZN(new_n371));
  XOR2_X1   g185(.A(G116), .B(G119), .Z(new_n372));
  XNOR2_X1  g186(.A(KEYINPUT2), .B(G113), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G113), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT2), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT2), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G113), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G116), .B(G119), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n371), .B1(new_n374), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n372), .A2(new_n373), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(new_n380), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(KEYINPUT67), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n370), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n369), .A3(new_n357), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  XOR2_X1   g204(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n391));
  INV_X1    g205(.A(KEYINPUT28), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n390), .A2(new_n391), .B1(new_n392), .B2(new_n389), .ZN(new_n393));
  XNOR2_X1  g207(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n394), .B(G101), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n199), .A2(G210), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n395), .B(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(KEYINPUT29), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n357), .A2(new_n369), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n399), .B1(new_n357), .B2(new_n369), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n387), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT68), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g218(.A(KEYINPUT68), .B(new_n387), .C1(new_n400), .C2(new_n401), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n389), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n398), .B1(new_n408), .B2(new_n397), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n390), .A2(KEYINPUT28), .ZN(new_n410));
  INV_X1    g224(.A(new_n389), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n411), .A2(KEYINPUT28), .ZN(new_n412));
  INV_X1    g226(.A(new_n397), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT29), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n410), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n416), .A2(KEYINPUT72), .A3(new_n264), .ZN(new_n417));
  AOI21_X1  g231(.A(KEYINPUT72), .B1(new_n416), .B2(new_n264), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n330), .B1(new_n409), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n393), .A2(new_n397), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n389), .A2(new_n397), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT69), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT69), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n389), .A2(new_n425), .A3(new_n397), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n406), .A2(KEYINPUT70), .A3(KEYINPUT31), .A4(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n404), .A2(new_n405), .B1(new_n424), .B2(new_n426), .ZN(new_n430));
  AOI21_X1  g244(.A(KEYINPUT31), .B1(new_n430), .B2(KEYINPUT70), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n422), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT32), .ZN(new_n433));
  NOR2_X1   g247(.A1(G472), .A2(G902), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n360), .A2(new_n364), .A3(new_n368), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n336), .A2(new_n339), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n355), .A2(G128), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n365), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n361), .A2(new_n362), .A3(new_n347), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT30), .B1(new_n436), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n357), .A2(new_n369), .A3(new_n399), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(KEYINPUT68), .B1(new_n444), .B2(new_n387), .ZN(new_n445));
  AOI211_X1 g259(.A(new_n403), .B(new_n386), .C1(new_n442), .C2(new_n443), .ZN(new_n446));
  OAI211_X1 g260(.A(KEYINPUT70), .B(new_n427), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT31), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n421), .B1(new_n449), .B2(new_n428), .ZN(new_n450));
  INV_X1    g264(.A(new_n434), .ZN(new_n451));
  OAI21_X1  g265(.A(KEYINPUT32), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n420), .B1(new_n435), .B2(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(G110), .B(G140), .ZN(new_n454));
  INV_X1    g268(.A(G227), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(G953), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n454), .B(new_n456), .Z(new_n457));
  NAND2_X1  g271(.A1(new_n439), .A2(new_n440), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n227), .A2(G107), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n227), .A2(G107), .ZN(new_n461));
  OAI21_X1  g275(.A(G101), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(KEYINPUT3), .B1(new_n227), .B2(G107), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT3), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(new_n294), .A3(G104), .ZN(new_n465));
  INV_X1    g279(.A(G101), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n463), .A2(new_n465), .A3(new_n466), .A4(new_n459), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n458), .A2(KEYINPUT10), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n463), .A2(new_n465), .A3(new_n459), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(KEYINPUT4), .A3(new_n467), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT4), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n471), .A2(new_n474), .A3(G101), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n473), .A2(new_n475), .A3(new_n364), .A4(new_n368), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT1), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n477), .B1(new_n232), .B2(new_n235), .ZN(new_n478));
  OAI22_X1  g292(.A1(new_n478), .A2(new_n346), .B1(new_n341), .B2(new_n345), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n468), .B1(new_n479), .B2(new_n440), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n470), .B(new_n476), .C1(new_n480), .C2(KEYINPUT10), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n457), .B1(new_n481), .B2(new_n360), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT74), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n479), .A2(new_n440), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n469), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT10), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n360), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n487), .A2(new_n488), .A3(new_n476), .A4(new_n470), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT74), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n489), .A2(new_n490), .A3(new_n457), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n481), .A2(new_n360), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n483), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n439), .A2(new_n440), .A3(new_n468), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n485), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(KEYINPUT12), .B1(new_n495), .B2(new_n360), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT12), .ZN(new_n497));
  AOI211_X1 g311(.A(new_n497), .B(new_n488), .C1(new_n485), .C2(new_n494), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n489), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n457), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n493), .A2(new_n501), .A3(G469), .ZN(new_n502));
  INV_X1    g316(.A(G469), .ZN(new_n503));
  INV_X1    g317(.A(new_n498), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n495), .A2(new_n360), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n497), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n482), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n457), .B1(new_n489), .B2(new_n492), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n503), .B(new_n264), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n503), .A2(new_n264), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n502), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(G221), .B1(new_n273), .B2(G902), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n453), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(G214), .B1(G237), .B2(G902), .ZN(new_n516));
  XOR2_X1   g330(.A(new_n516), .B(KEYINPUT75), .Z(new_n517));
  NAND4_X1  g331(.A1(new_n382), .A2(new_n473), .A3(new_n385), .A4(new_n475), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT5), .ZN(new_n519));
  INV_X1    g333(.A(G119), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n520), .A3(G116), .ZN(new_n521));
  OAI211_X1 g335(.A(G113), .B(new_n521), .C1(new_n372), .C2(new_n519), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n469), .A2(new_n384), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT76), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(G110), .B(G122), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT77), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n518), .A2(KEYINPUT76), .A3(new_n523), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n526), .A2(KEYINPUT6), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n518), .A2(KEYINPUT76), .A3(new_n523), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT76), .B1(new_n518), .B2(new_n523), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n532), .A2(new_n533), .A3(new_n528), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n518), .A2(new_n523), .A3(new_n527), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT6), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n531), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n458), .A2(new_n210), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n368), .A2(new_n364), .A3(G125), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(G224), .A3(new_n320), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n320), .A2(G224), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n539), .A2(new_n543), .A3(new_n540), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n538), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT78), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n522), .A2(new_n384), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT80), .B1(new_n550), .B2(new_n468), .ZN(new_n551));
  OR2_X1    g365(.A1(new_n551), .A2(new_n523), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n523), .ZN(new_n553));
  XOR2_X1   g367(.A(KEYINPUT79), .B(KEYINPUT8), .Z(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(new_n527), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n535), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n543), .A2(KEYINPUT7), .ZN(new_n558));
  XOR2_X1   g372(.A(new_n541), .B(new_n558), .Z(new_n559));
  OAI21_X1  g373(.A(new_n264), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n538), .A2(KEYINPUT78), .A3(new_n546), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n549), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(G210), .B1(G237), .B2(G902), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n526), .A2(new_n529), .A3(new_n530), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n536), .ZN(new_n568));
  AOI211_X1 g382(.A(new_n548), .B(new_n545), .C1(new_n568), .C2(new_n531), .ZN(new_n569));
  AOI21_X1  g383(.A(KEYINPUT78), .B1(new_n538), .B2(new_n546), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(new_n564), .A3(new_n561), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n517), .B1(new_n566), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n274), .B1(G234), .B2(new_n264), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n215), .A2(new_n235), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n520), .A2(G128), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT23), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT23), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n520), .B2(G128), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n578), .B(new_n580), .C1(G119), .C2(new_n346), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(G110), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT73), .B1(new_n346), .B2(G119), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT73), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(new_n520), .A3(G128), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n577), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  XOR2_X1   g400(.A(KEYINPUT24), .B(G110), .Z(new_n587));
  NOR2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n576), .B(new_n222), .C1(new_n582), .C2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n581), .A2(G110), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n586), .A2(new_n587), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n590), .B(new_n591), .C1(new_n217), .C2(new_n223), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n320), .A2(G221), .A3(G234), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(KEYINPUT22), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(new_n333), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n596), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(new_n592), .A3(new_n589), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(new_n264), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT25), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n597), .A2(KEYINPUT25), .A3(new_n264), .A4(new_n599), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n575), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n600), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n604), .B1(new_n575), .B2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n329), .A2(new_n515), .A3(new_n573), .A4(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  NAND2_X1  g422(.A1(new_n566), .A2(new_n572), .ZN(new_n609));
  INV_X1    g423(.A(new_n517), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n327), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n514), .ZN(new_n612));
  OAI21_X1  g426(.A(G472), .B1(new_n450), .B2(G902), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n432), .A2(new_n434), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n606), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n611), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n307), .A2(KEYINPUT33), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n300), .A2(new_n619), .A3(new_n306), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n618), .A2(G478), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n316), .A2(new_n310), .ZN(new_n622));
  NAND2_X1  g436(.A1(G478), .A2(G902), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n263), .A2(new_n269), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT86), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n263), .A2(KEYINPUT86), .A3(new_n269), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n624), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n617), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT34), .B(G104), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  NAND3_X1  g446(.A1(new_n259), .A2(KEYINPUT92), .A3(new_n261), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n262), .ZN(new_n634));
  AOI21_X1  g448(.A(KEYINPUT92), .B1(new_n259), .B2(new_n261), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n319), .B(new_n269), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n617), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G107), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  NAND2_X1  g454(.A1(new_n609), .A2(new_n610), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n596), .A2(KEYINPUT36), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n593), .B(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n574), .A2(G902), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n604), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT93), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n641), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n615), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n329), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT94), .B(KEYINPUT37), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G110), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n651), .B(new_n653), .ZN(G12));
  OR2_X1    g468(.A1(new_n326), .A2(G900), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n323), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n636), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n515), .A2(new_n649), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G128), .ZN(G30));
  XNOR2_X1  g474(.A(new_n609), .B(KEYINPUT38), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n319), .B1(new_n270), .B2(new_n271), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n430), .B1(new_n390), .B2(new_n413), .ZN(new_n664));
  OAI21_X1  g478(.A(G472), .B1(new_n664), .B2(G902), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n433), .B1(new_n432), .B2(new_n434), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n450), .A2(KEYINPUT32), .A3(new_n451), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n647), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n517), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n661), .A2(new_n663), .A3(new_n668), .A4(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(KEYINPUT95), .Z(new_n672));
  XOR2_X1   g486(.A(new_n656), .B(KEYINPUT39), .Z(new_n673));
  NOR2_X1   g487(.A1(new_n514), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n672), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(new_n232), .ZN(G45));
  INV_X1    g493(.A(KEYINPUT96), .ZN(new_n680));
  INV_X1    g494(.A(new_n420), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n681), .B1(new_n666), .B2(new_n667), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT93), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n647), .B(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n682), .A2(new_n573), .A3(new_n612), .A4(new_n684), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n686), .B(new_n656), .C1(new_n270), .C2(new_n271), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n680), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n687), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n689), .A2(new_n515), .A3(new_n649), .A4(KEYINPUT96), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  NOR2_X1   g506(.A1(new_n453), .A2(new_n616), .ZN(new_n693));
  INV_X1    g507(.A(new_n611), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n504), .A2(new_n506), .ZN(new_n695));
  INV_X1    g509(.A(new_n482), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n508), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g511(.A(G469), .B1(new_n697), .B2(G902), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n698), .A2(new_n513), .A3(new_n509), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n693), .A2(new_n694), .A3(new_n629), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT41), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G113), .ZN(G15));
  NAND4_X1  g516(.A1(new_n693), .A2(new_n694), .A3(new_n637), .A4(new_n699), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G116), .ZN(G18));
  AOI21_X1  g518(.A(new_n564), .B1(new_n571), .B2(new_n561), .ZN(new_n705));
  NOR4_X1   g519(.A1(new_n569), .A2(new_n570), .A3(new_n565), .A4(new_n560), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n699), .B(new_n610), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT97), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT97), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n609), .A2(new_n709), .A3(new_n610), .A4(new_n699), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n453), .A2(new_n648), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n329), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G119), .ZN(G21));
  NOR2_X1   g528(.A1(new_n662), .A2(new_n641), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n410), .A2(new_n412), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n413), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n717), .B1(new_n429), .B2(new_n431), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n434), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n613), .A2(new_n719), .A3(new_n606), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT98), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n613), .A2(new_n719), .A3(KEYINPUT98), .A4(new_n606), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n699), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n328), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n715), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G122), .ZN(G24));
  NAND3_X1  g542(.A1(new_n613), .A2(new_n719), .A3(new_n669), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n687), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n711), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G125), .ZN(G27));
  INV_X1    g546(.A(KEYINPUT100), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT42), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT99), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n512), .A2(new_n735), .A3(new_n513), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n735), .B1(new_n512), .B2(new_n513), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n705), .A2(new_n706), .A3(new_n517), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n682), .A2(new_n606), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n734), .B1(new_n740), .B2(new_n687), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n566), .A2(new_n572), .A3(new_n610), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n453), .A2(new_n616), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(KEYINPUT100), .B(KEYINPUT42), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n743), .A2(new_n689), .A3(new_n738), .A4(new_n745), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n741), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n189), .ZN(G33));
  NAND3_X1  g562(.A1(new_n743), .A2(new_n658), .A3(new_n738), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G134), .ZN(G36));
  NOR2_X1   g564(.A1(new_n270), .A2(new_n271), .ZN(new_n751));
  AND2_X1   g565(.A1(KEYINPUT101), .A2(KEYINPUT43), .ZN(new_n752));
  NOR2_X1   g566(.A1(KEYINPUT101), .A2(KEYINPUT43), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n751), .B(new_n686), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n627), .A2(new_n628), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n624), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n754), .B1(new_n756), .B2(new_n752), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n647), .B1(new_n613), .B2(new_n614), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT102), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n739), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  XOR2_X1   g576(.A(new_n762), .B(KEYINPUT103), .Z(new_n763));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n493), .A2(new_n501), .ZN(new_n765));
  XOR2_X1   g579(.A(new_n765), .B(KEYINPUT45), .Z(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n503), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n764), .B1(new_n767), .B2(new_n510), .ZN(new_n768));
  OAI211_X1 g582(.A(KEYINPUT46), .B(new_n511), .C1(new_n766), .C2(new_n503), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n509), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n513), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n673), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n760), .A2(new_n761), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n774), .A2(KEYINPUT104), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(KEYINPUT104), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n773), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n763), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT105), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(new_n333), .ZN(G39));
  INV_X1    g594(.A(KEYINPUT47), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n771), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n770), .A2(KEYINPUT47), .A3(new_n513), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n682), .A2(new_n606), .A3(new_n742), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n689), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT106), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(new_n212), .ZN(G42));
  AND2_X1   g602(.A1(new_n698), .A2(new_n509), .ZN(new_n789));
  NOR2_X1   g603(.A1(KEYINPUT107), .A2(KEYINPUT49), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(KEYINPUT107), .A2(KEYINPUT49), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n610), .A2(new_n513), .A3(new_n792), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n661), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n668), .A2(new_n616), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n756), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n656), .B(KEYINPUT111), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n647), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT112), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n715), .A2(new_n612), .A3(new_n668), .A4(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n691), .A2(new_n659), .A3(new_n731), .A4(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n688), .A2(new_n690), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n800), .A2(new_n731), .A3(new_n659), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT108), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n684), .A2(new_n315), .A3(new_n318), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n453), .A2(new_n809), .A3(new_n514), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n633), .A2(new_n262), .ZN(new_n811));
  INV_X1    g625(.A(new_n635), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n811), .A2(new_n812), .B1(G475), .B2(new_n268), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n514), .A2(KEYINPUT99), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n512), .A2(new_n735), .A3(new_n513), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n729), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n810), .A2(new_n813), .B1(new_n817), .B2(new_n629), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n739), .A2(new_n656), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n808), .B(new_n749), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n648), .A2(new_n319), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n813), .A2(new_n682), .A3(new_n612), .A4(new_n821), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n613), .A2(new_n719), .A3(new_n669), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n755), .A2(new_n823), .A3(new_n686), .A4(new_n738), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n819), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n637), .A2(new_n656), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n740), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT108), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n820), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n747), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n627), .A2(new_n319), .A3(new_n628), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n831), .B1(new_n751), .B2(new_n624), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n617), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n727), .A2(new_n833), .A3(new_n607), .A4(new_n703), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n713), .A2(new_n700), .A3(new_n651), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AND4_X1   g650(.A1(KEYINPUT109), .A2(new_n829), .A3(new_n830), .A4(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n747), .B1(new_n820), .B2(new_n828), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT109), .B1(new_n838), .B2(new_n836), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n807), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT53), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n800), .A2(KEYINPUT52), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT110), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n731), .A2(new_n843), .A3(new_n659), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n843), .B1(new_n731), .B2(new_n659), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n691), .B(new_n842), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n806), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT113), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT113), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n846), .A2(new_n849), .A3(new_n806), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n829), .A2(new_n836), .A3(new_n830), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT109), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n838), .A2(KEYINPUT109), .A3(new_n836), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n851), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n841), .A2(new_n858), .A3(KEYINPUT54), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n852), .A2(new_n857), .ZN(new_n860));
  INV_X1    g674(.A(new_n850), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n849), .B1(new_n846), .B2(new_n806), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n854), .A2(new_n855), .B1(new_n806), .B2(new_n803), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n863), .B(new_n864), .C1(new_n865), .C2(KEYINPUT53), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n859), .A2(KEYINPUT114), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT114), .B1(new_n859), .B2(new_n866), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n784), .A2(KEYINPUT116), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n782), .A2(new_n870), .A3(new_n783), .ZN(new_n871));
  INV_X1    g685(.A(new_n789), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n869), .B(new_n871), .C1(new_n513), .C2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT115), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n323), .B1(new_n722), .B2(new_n723), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n757), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n874), .B1(new_n877), .B2(new_n742), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(KEYINPUT115), .A3(new_n739), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n873), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n742), .A2(new_n725), .A3(new_n323), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n757), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n823), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n795), .A2(new_n751), .A3(new_n624), .A4(new_n881), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n661), .A2(new_n610), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n757), .A2(new_n699), .A3(new_n875), .A4(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n888), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n885), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n880), .A2(new_n883), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT51), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n321), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n872), .A2(new_n513), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n878), .B(new_n879), .C1(new_n784), .C2(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n891), .A2(KEYINPUT118), .A3(new_n883), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT118), .B1(new_n891), .B2(new_n883), .ZN(new_n898));
  OAI211_X1 g712(.A(KEYINPUT51), .B(new_n896), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n882), .A2(new_n693), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT48), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n876), .A2(new_n711), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n894), .A2(new_n899), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n795), .A2(new_n629), .A3(new_n881), .ZN(new_n904));
  NOR4_X1   g718(.A1(new_n867), .A2(new_n868), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(G952), .A2(G953), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT119), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n796), .B1(new_n905), .B2(new_n907), .ZN(G75));
  NAND2_X1  g722(.A1(new_n840), .A2(new_n857), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n264), .B1(new_n909), .B2(new_n863), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(G210), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT56), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n538), .B(new_n545), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT55), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n914), .B1(new_n911), .B2(new_n912), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n320), .A2(G952), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(G51));
  NAND2_X1  g732(.A1(new_n910), .A2(new_n767), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT121), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n697), .B(KEYINPUT120), .Z(new_n921));
  OAI21_X1  g735(.A(new_n863), .B1(new_n865), .B2(KEYINPUT53), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT54), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n866), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n510), .B(KEYINPUT57), .Z(new_n926));
  OAI21_X1  g740(.A(new_n921), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n917), .B1(new_n920), .B2(new_n927), .ZN(G54));
  NAND3_X1  g742(.A1(new_n910), .A2(KEYINPUT58), .A3(G475), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n929), .A2(new_n260), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n260), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n930), .A2(new_n931), .A3(new_n917), .ZN(G60));
  XNOR2_X1  g746(.A(new_n623), .B(KEYINPUT59), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(new_n867), .B2(new_n868), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n618), .A2(new_n620), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n917), .ZN(new_n938));
  INV_X1    g752(.A(new_n866), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n864), .B1(new_n909), .B2(new_n863), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n935), .B(new_n933), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT122), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT122), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n924), .A2(new_n943), .A3(new_n935), .A4(new_n933), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n937), .A2(new_n938), .A3(new_n945), .ZN(G63));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g761(.A1(G217), .A2(G902), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT60), .Z(new_n949));
  NAND2_X1  g763(.A1(new_n922), .A2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n597), .A2(new_n599), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n922), .A2(KEYINPUT123), .A3(new_n949), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n938), .ZN(new_n956));
  INV_X1    g770(.A(new_n643), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n952), .B2(new_n954), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n947), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n958), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n960), .A2(KEYINPUT61), .A3(new_n938), .A4(new_n955), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n959), .A2(new_n961), .ZN(G66));
  INV_X1    g776(.A(new_n836), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n320), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n324), .A2(G224), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n964), .B(KEYINPUT124), .C1(new_n320), .C2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(KEYINPUT124), .B2(new_n964), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n568), .B(new_n531), .C1(G898), .C2(new_n320), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n967), .B(new_n968), .Z(G69));
  NAND2_X1  g783(.A1(new_n244), .A2(new_n245), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n444), .B(new_n970), .Z(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT126), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n455), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n320), .B1(new_n974), .B2(G900), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n832), .A2(new_n743), .A3(new_n674), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT125), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n977), .A2(new_n978), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n786), .A2(new_n980), .ZN(new_n981));
  AOI211_X1 g795(.A(new_n979), .B(new_n981), .C1(new_n763), .C2(new_n777), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n691), .B1(new_n844), .B2(new_n845), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n678), .A2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT62), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n982), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n972), .B1(new_n988), .B2(G953), .ZN(new_n989));
  NAND2_X1  g803(.A1(G900), .A2(G953), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n827), .B1(new_n763), .B2(new_n777), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n715), .A2(new_n693), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n747), .B1(new_n772), .B2(new_n992), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n991), .A2(new_n786), .A3(new_n984), .A4(new_n993), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n971), .B(new_n990), .C1(new_n994), .C2(G953), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n989), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n976), .B1(new_n996), .B2(new_n973), .ZN(new_n997));
  AOI211_X1 g811(.A(KEYINPUT126), .B(new_n975), .C1(new_n989), .C2(new_n995), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n997), .A2(new_n998), .ZN(G72));
  NAND3_X1  g813(.A1(new_n982), .A2(new_n987), .A3(new_n836), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT127), .ZN(new_n1001));
  NAND2_X1  g815(.A1(G472), .A2(G902), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT63), .Z(new_n1003));
  AND3_X1   g817(.A1(new_n1000), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1001), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1005));
  NOR4_X1   g819(.A1(new_n1004), .A2(new_n1005), .A3(new_n413), .A4(new_n408), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1003), .B1(new_n994), .B2(new_n963), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1007), .A2(new_n413), .A3(new_n408), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n430), .B1(new_n407), .B2(new_n413), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n841), .A2(new_n858), .A3(new_n1003), .ZN(new_n1010));
  OAI211_X1 g824(.A(new_n1008), .B(new_n938), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1006), .A2(new_n1011), .ZN(G57));
endmodule


