//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n192), .B(KEYINPUT22), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(G137), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT78), .ZN(new_n195));
  XOR2_X1   g009(.A(G119), .B(G128), .Z(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT24), .B(G110), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT23), .B1(new_n199), .B2(G119), .ZN(new_n200));
  AOI21_X1  g014(.A(KEYINPUT74), .B1(new_n199), .B2(G119), .ZN(new_n201));
  XNOR2_X1  g015(.A(new_n200), .B(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n198), .B1(new_n202), .B2(G110), .ZN(new_n203));
  INV_X1    g017(.A(G140), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G125), .ZN(new_n205));
  INV_X1    g019(.A(G125), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G140), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT16), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(new_n204), .A3(G125), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT75), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n205), .A2(new_n207), .A3(KEYINPUT16), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n211), .A2(new_n204), .A3(KEYINPUT75), .A4(G125), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n214), .A2(new_n215), .A3(G146), .A4(new_n216), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n217), .A2(KEYINPUT76), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n217), .A2(KEYINPUT76), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n203), .B(new_n210), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT77), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n214), .A2(new_n216), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT76), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n223), .A2(new_n224), .A3(G146), .A4(new_n215), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n217), .A2(KEYINPUT76), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n209), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT77), .A3(new_n203), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n215), .A2(new_n214), .A3(new_n216), .ZN(new_n230));
  INV_X1    g044(.A(G146), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n217), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n202), .A2(G110), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n196), .A2(new_n197), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n233), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n195), .B1(new_n229), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n237), .ZN(new_n239));
  AOI211_X1 g053(.A(KEYINPUT78), .B(new_n239), .C1(new_n222), .C2(new_n228), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n194), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n239), .B1(new_n222), .B2(new_n228), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n195), .ZN(new_n243));
  INV_X1    g057(.A(new_n194), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n241), .A2(new_n188), .A3(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n247), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n241), .A2(new_n188), .A3(new_n245), .A4(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n190), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n240), .A2(new_n194), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n220), .A2(new_n221), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT77), .B1(new_n227), .B2(new_n203), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n237), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT78), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n243), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n252), .B1(new_n257), .B2(new_n194), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n258), .A2(new_n188), .A3(new_n190), .ZN(new_n259));
  OR2_X1    g073(.A1(new_n251), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G131), .ZN(new_n261));
  INV_X1    g075(.A(G134), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT67), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G134), .ZN(new_n265));
  INV_X1    g079(.A(G137), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n263), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT68), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n268), .B1(new_n262), .B2(G137), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n261), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(KEYINPUT68), .B2(new_n267), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n263), .A2(new_n265), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n266), .A2(KEYINPUT11), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n266), .A2(KEYINPUT11), .A3(G134), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT11), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G137), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n274), .A2(new_n261), .A3(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G143), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(G146), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n231), .A2(G143), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT1), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G128), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n199), .A2(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n231), .A2(G143), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n280), .A2(G146), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n271), .A2(new_n279), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n287), .A2(new_n288), .ZN(new_n292));
  OR3_X1    g106(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n293));
  AND2_X1   g107(.A1(KEYINPUT0), .A2(G128), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n292), .A2(new_n293), .A3(new_n295), .A4(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n287), .A2(new_n288), .A3(new_n294), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT65), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(G143), .B(G146), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(KEYINPUT65), .A3(new_n294), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n297), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n303), .A2(KEYINPUT66), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n263), .A2(new_n265), .B1(KEYINPUT11), .B2(new_n266), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n275), .A2(new_n277), .ZN(new_n306));
  OAI21_X1  g120(.A(G131), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n279), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n297), .A2(new_n300), .A3(new_n302), .A4(KEYINPUT66), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n291), .B1(new_n304), .B2(new_n310), .ZN(new_n311));
  AND2_X1   g125(.A1(KEYINPUT2), .A2(G113), .ZN(new_n312));
  NOR2_X1   g126(.A1(KEYINPUT2), .A2(G113), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(G116), .B(G119), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT69), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n314), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n319), .B1(new_n314), .B2(new_n316), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n318), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n311), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT28), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n271), .A2(new_n279), .A3(new_n290), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT70), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n308), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n279), .A2(new_n307), .A3(KEYINPUT70), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n325), .B1(new_n329), .B2(new_n303), .ZN(new_n330));
  INV_X1    g144(.A(new_n322), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n324), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n279), .A2(new_n307), .A3(KEYINPUT70), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT70), .B1(new_n279), .B2(new_n307), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n303), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AND4_X1   g149(.A1(new_n324), .A2(new_n335), .A3(new_n331), .A4(new_n291), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n323), .B1(new_n332), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n338));
  INV_X1    g152(.A(G237), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n191), .A3(G210), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n338), .B(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT26), .B(G101), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n341), .B(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n337), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT30), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n311), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n335), .A2(KEYINPUT30), .A3(new_n291), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n347), .A3(new_n322), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT31), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n330), .A2(new_n331), .ZN(new_n350));
  INV_X1    g164(.A(new_n343), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n348), .A2(new_n349), .A3(new_n350), .A4(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n348), .A2(new_n350), .A3(new_n351), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT31), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n344), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(G472), .A2(G902), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT32), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n355), .A2(KEYINPUT32), .A3(new_n356), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(KEYINPUT72), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT72), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n357), .A2(new_n362), .A3(new_n358), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  OR2_X1    g178(.A1(new_n332), .A2(new_n336), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n330), .A2(new_n331), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(KEYINPUT29), .A3(new_n351), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT29), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n337), .A2(new_n343), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT73), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n348), .A2(new_n350), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n371), .B1(new_n372), .B2(new_n343), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n369), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n337), .A2(new_n371), .A3(new_n343), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n368), .B(new_n188), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G472), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n260), .B1(new_n364), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT98), .ZN(new_n379));
  XOR2_X1   g193(.A(KEYINPUT9), .B(G234), .Z(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(G221), .B1(new_n381), .B2(G902), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G469), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(new_n188), .ZN(new_n385));
  XOR2_X1   g199(.A(G110), .B(G140), .Z(new_n386));
  INV_X1    g200(.A(G227), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(G953), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n386), .B(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n389), .B(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G104), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT3), .B1(new_n393), .B2(G107), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT3), .ZN(new_n395));
  INV_X1    g209(.A(G107), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n396), .A3(G104), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n393), .A2(G107), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n394), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G101), .ZN(new_n400));
  INV_X1    g214(.A(G101), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n394), .A2(new_n397), .A3(new_n401), .A4(new_n398), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(KEYINPUT4), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT4), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n399), .A2(new_n404), .A3(G101), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n297), .A2(new_n300), .A3(new_n302), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT82), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT82), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n303), .A2(new_n409), .A3(new_n403), .A4(new_n405), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n329), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n289), .A2(KEYINPUT84), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT84), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n301), .A2(new_n414), .A3(new_n286), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n413), .A2(new_n285), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT83), .ZN(new_n417));
  XNOR2_X1  g231(.A(G104), .B(G107), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n417), .B1(new_n418), .B2(new_n401), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n396), .A2(G104), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n393), .A2(G107), .ZN(new_n421));
  OAI211_X1 g235(.A(KEYINPUT83), .B(G101), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n419), .A2(new_n402), .A3(new_n422), .ZN(new_n423));
  OR2_X1    g237(.A1(new_n416), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT10), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n289), .ZN(new_n427));
  OAI22_X1  g241(.A1(new_n286), .A2(new_n288), .B1(new_n287), .B2(G128), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n423), .A2(new_n429), .A3(new_n425), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n411), .A2(new_n412), .A3(new_n426), .A4(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n430), .B1(new_n408), .B2(new_n410), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n412), .B1(new_n434), .B2(new_n426), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n392), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n416), .A2(new_n423), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n423), .A2(new_n429), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT85), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n423), .A2(new_n429), .A3(KEYINPUT85), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n437), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n308), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT12), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n441), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT85), .B1(new_n423), .B2(new_n429), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n424), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT12), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n448), .A3(new_n329), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n432), .A2(new_n444), .A3(new_n449), .A4(new_n391), .ZN(new_n450));
  AOI21_X1  g264(.A(G902), .B1(new_n436), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n385), .B1(new_n451), .B2(new_n384), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n432), .A2(new_n444), .A3(new_n449), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n392), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n411), .A2(new_n426), .A3(new_n431), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n329), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(new_n432), .A3(new_n391), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(G469), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n383), .B1(new_n452), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n339), .A2(new_n191), .A3(G214), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n280), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n339), .A2(new_n191), .A3(G143), .A4(G214), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(KEYINPUT18), .A2(G131), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n208), .B(G146), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n461), .A2(new_n462), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT90), .B1(new_n468), .B2(new_n464), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT90), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n463), .A2(new_n470), .A3(new_n465), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n466), .B(new_n467), .C1(new_n469), .C2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(G113), .B(G122), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(new_n393), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(KEYINPUT92), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n463), .A2(G131), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT17), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n461), .A2(new_n261), .A3(new_n462), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n463), .A2(KEYINPUT17), .A3(G131), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n479), .A2(new_n217), .A3(new_n232), .A4(new_n480), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n472), .A2(new_n475), .A3(new_n481), .ZN(new_n482));
  OR3_X1    g296(.A1(new_n208), .A2(KEYINPUT91), .A3(KEYINPUT19), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n208), .A2(KEYINPUT19), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT91), .B1(new_n208), .B2(KEYINPUT19), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n483), .A2(new_n231), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n476), .A2(new_n478), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n486), .B(new_n487), .C1(new_n218), .C2(new_n219), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n474), .B1(new_n488), .B2(new_n472), .ZN(new_n489));
  OR2_X1    g303(.A1(new_n482), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT20), .ZN(new_n491));
  INV_X1    g305(.A(G475), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n490), .A2(new_n491), .A3(new_n492), .A4(new_n188), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n492), .B(new_n188), .C1(new_n482), .C2(new_n489), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT20), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(KEYINPUT93), .A3(new_n495), .ZN(new_n496));
  OR3_X1    g310(.A1(new_n494), .A2(KEYINPUT93), .A3(KEYINPUT20), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n474), .B1(new_n472), .B2(new_n481), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n188), .B1(new_n482), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(G475), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n496), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G122), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G116), .ZN(new_n503));
  INV_X1    g317(.A(G116), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G122), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(new_n505), .A3(new_n396), .ZN(new_n506));
  XOR2_X1   g320(.A(new_n506), .B(KEYINPUT94), .Z(new_n507));
  OR3_X1    g321(.A1(new_n502), .A2(KEYINPUT14), .A3(G116), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(KEYINPUT14), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n509), .A3(new_n503), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n280), .A2(G128), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n199), .A2(G143), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n272), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n199), .A2(G143), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n280), .A2(G128), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n263), .B(new_n265), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  AOI22_X1  g330(.A1(G107), .A2(new_n510), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n507), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n280), .A2(KEYINPUT13), .A3(G128), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n512), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT13), .B1(new_n280), .B2(G128), .ZN(new_n521));
  OAI21_X1  g335(.A(G134), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n522), .A2(new_n513), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n503), .A2(new_n505), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G107), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n506), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n518), .A2(new_n527), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n381), .A2(new_n187), .A3(G953), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n518), .A2(new_n527), .A3(new_n529), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n188), .ZN(new_n534));
  INV_X1    g348(.A(G478), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n534), .B(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n501), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n459), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(G210), .B1(G237), .B2(G902), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n297), .A2(new_n300), .A3(new_n302), .A4(G125), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n206), .B1(new_n427), .B2(new_n428), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(G224), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT7), .B1(new_n545), .B2(G953), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(G953), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n547), .B1(new_n542), .B2(new_n543), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n544), .A2(new_n546), .B1(new_n548), .B2(KEYINPUT7), .ZN(new_n549));
  INV_X1    g363(.A(G119), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(G116), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n504), .A2(G119), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n552), .A3(KEYINPUT5), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n553), .B(G113), .C1(KEYINPUT5), .C2(new_n551), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n554), .B1(new_n320), .B2(new_n321), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT86), .B1(new_n555), .B2(new_n423), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n314), .A2(new_n316), .A3(new_n319), .ZN(new_n557));
  OR2_X1    g371(.A1(KEYINPUT2), .A2(G113), .ZN(new_n558));
  NAND2_X1  g372(.A1(KEYINPUT2), .A2(G113), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n558), .A2(new_n551), .A3(new_n552), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT69), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n504), .A2(KEYINPUT5), .A3(G119), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n562), .B1(new_n316), .B2(KEYINPUT5), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n557), .A2(new_n561), .B1(new_n563), .B2(G113), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n419), .A2(new_n402), .A3(new_n422), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT86), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n322), .A2(new_n405), .A3(new_n403), .ZN(new_n568));
  XNOR2_X1  g382(.A(G110), .B(G122), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n556), .A2(new_n567), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(KEYINPUT8), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n564), .A2(new_n565), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n555), .A2(new_n423), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n549), .A2(new_n570), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n188), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT88), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n575), .A2(KEYINPUT88), .A3(new_n188), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g394(.A(new_n544), .B(new_n547), .Z(new_n581));
  NAND3_X1  g395(.A1(new_n556), .A2(new_n567), .A3(new_n568), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n569), .A2(KEYINPUT87), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n582), .A2(KEYINPUT6), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT6), .B1(new_n582), .B2(new_n583), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n581), .B1(new_n586), .B2(new_n570), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n541), .B1(new_n580), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT89), .ZN(new_n589));
  INV_X1    g403(.A(new_n585), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n582), .A2(KEYINPUT6), .A3(new_n583), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n570), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n581), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n594), .A2(new_n540), .A3(new_n579), .A4(new_n578), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n588), .A2(new_n589), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT21), .B(G898), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT96), .ZN(new_n598));
  NAND2_X1  g412(.A1(G234), .A2(G237), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n599), .A2(G902), .A3(G953), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT95), .B(G952), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(G953), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n599), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(new_n606), .B(KEYINPUT97), .Z(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(G214), .B1(G237), .B2(G902), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n580), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n612), .A2(KEYINPUT89), .A3(new_n540), .A4(new_n594), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n596), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n379), .B1(new_n539), .B2(new_n614), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n596), .A2(new_n611), .A3(new_n613), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n616), .A2(KEYINPUT98), .A3(new_n538), .A4(new_n459), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n378), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  AND2_X1   g433(.A1(new_n355), .A2(new_n356), .ZN(new_n620));
  INV_X1    g434(.A(G472), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n355), .B2(new_n188), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT99), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT99), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n355), .A2(new_n188), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n624), .B1(new_n625), .B2(new_n621), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n459), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n627), .A2(new_n260), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n610), .B1(new_n588), .B2(new_n595), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n607), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n531), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n533), .A2(new_n633), .A3(KEYINPUT33), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT33), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n531), .B(new_n532), .C1(new_n632), .C2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(G478), .A3(new_n188), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT101), .B(G478), .Z(new_n639));
  NAND2_X1  g453(.A1(new_n534), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n501), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n631), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n629), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT34), .B(G104), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  NAND2_X1  g460(.A1(new_n537), .A2(new_n500), .ZN(new_n647));
  AOI211_X1 g461(.A(new_n647), .B(new_n631), .C1(new_n493), .C2(new_n495), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n629), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(new_n396), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT102), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT35), .ZN(G9));
  INV_X1    g466(.A(new_n627), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n249), .B1(new_n258), .B2(new_n188), .ZN(new_n654));
  INV_X1    g468(.A(new_n250), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n189), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n244), .A2(KEYINPUT36), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n255), .B(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n188), .A3(new_n190), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n656), .A2(KEYINPUT103), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n661));
  INV_X1    g475(.A(new_n659), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n661), .B1(new_n251), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n615), .A2(new_n653), .A3(new_n617), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT37), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n666), .B(G110), .Z(G12));
  AOI22_X1  g481(.A1(new_n364), .A2(new_n377), .B1(new_n660), .B2(new_n663), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n493), .A2(new_n495), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n605), .B1(G900), .B2(new_n600), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n537), .A3(new_n500), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n668), .A2(new_n459), .A3(new_n630), .A4(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT104), .B(G128), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G30));
  NAND2_X1  g490(.A1(new_n596), .A2(new_n613), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(KEYINPUT105), .Z(new_n678));
  INV_X1    g492(.A(KEYINPUT38), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n366), .A2(new_n350), .A3(new_n343), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n188), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n343), .B1(new_n348), .B2(new_n350), .ZN(new_n683));
  OAI21_X1  g497(.A(G472), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n364), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n656), .A2(new_n659), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n670), .B(KEYINPUT39), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n459), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT40), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n680), .A2(new_n688), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n501), .A2(new_n537), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n609), .B(new_n694), .C1(new_n690), .C2(KEYINPUT40), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n280), .ZN(G45));
  NAND3_X1  g511(.A1(new_n501), .A2(new_n641), .A3(new_n670), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT106), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n668), .A2(new_n459), .A3(new_n630), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G146), .ZN(G48));
  XNOR2_X1  g515(.A(new_n451), .B(G469), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n382), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n378), .A2(new_n643), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT41), .B(G113), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT107), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n705), .B(new_n707), .ZN(G15));
  NAND3_X1  g522(.A1(new_n648), .A2(new_n378), .A3(new_n704), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G116), .ZN(G18));
  INV_X1    g524(.A(new_n630), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n703), .A2(new_n608), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n668), .A2(new_n538), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G119), .ZN(G21));
  NOR2_X1   g528(.A1(new_n251), .A2(new_n259), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n352), .B(new_n354), .C1(new_n367), .C2(new_n351), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n622), .B1(new_n356), .B2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n712), .A2(new_n715), .A3(new_n694), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G122), .ZN(G24));
  NAND2_X1  g533(.A1(new_n687), .A2(new_n717), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n698), .B(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n630), .A3(new_n704), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  NAND2_X1  g539(.A1(new_n360), .A2(KEYINPUT72), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT32), .B1(new_n355), .B2(new_n356), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n363), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n377), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n610), .B1(new_n596), .B2(new_n613), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n454), .A2(KEYINPUT108), .A3(new_n457), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n456), .A2(new_n734), .A3(new_n432), .A4(new_n391), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(G469), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n383), .B1(new_n737), .B2(new_n452), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n731), .A2(new_n732), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n732), .B1(new_n731), .B2(new_n738), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n730), .B(new_n715), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(KEYINPUT110), .B1(new_n741), .B2(new_n722), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  INV_X1    g557(.A(new_n740), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n731), .A2(new_n738), .A3(new_n732), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n746), .A2(new_n747), .A3(new_n378), .A4(new_n699), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n742), .A2(new_n743), .A3(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n620), .A2(KEYINPUT111), .A3(KEYINPUT32), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT111), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n360), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n377), .A2(new_n359), .A3(new_n750), .A4(new_n752), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n753), .A2(new_n699), .A3(new_n715), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n754), .A2(KEYINPUT112), .A3(KEYINPUT42), .A4(new_n746), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT42), .B1(new_n739), .B2(new_n740), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n753), .A2(new_n699), .A3(new_n715), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n749), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  NAND3_X1  g576(.A1(new_n746), .A2(new_n378), .A3(new_n673), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G134), .ZN(G36));
  NAND2_X1  g578(.A1(KEYINPUT45), .A2(G469), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n458), .A2(new_n765), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n766), .A2(KEYINPUT113), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n736), .A2(KEYINPUT45), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n766), .A2(KEYINPUT113), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n385), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(KEYINPUT46), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n451), .A2(new_n384), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n772), .A2(KEYINPUT114), .A3(new_n773), .ZN(new_n777));
  INV_X1    g591(.A(new_n770), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n385), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n776), .B(new_n777), .C1(new_n779), .C2(KEYINPUT46), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n780), .A2(new_n382), .A3(new_n689), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n627), .A2(new_n687), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n782), .A2(KEYINPUT115), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n496), .A2(new_n497), .A3(new_n500), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n641), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT43), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n782), .A2(KEYINPUT115), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n783), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n781), .A2(new_n791), .A3(new_n731), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  NAND2_X1  g608(.A1(new_n780), .A2(new_n382), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT47), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n730), .A2(new_n715), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT47), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n780), .A2(new_n798), .A3(new_n382), .ZN(new_n799));
  INV_X1    g613(.A(new_n731), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n722), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n796), .A2(new_n797), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G140), .ZN(G42));
  XNOR2_X1  g617(.A(new_n785), .B(KEYINPUT43), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT119), .B1(new_n804), .B2(new_n605), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n806));
  INV_X1    g620(.A(new_n605), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n787), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n800), .A2(new_n703), .ZN(new_n810));
  AND4_X1   g624(.A1(new_n715), .A2(new_n809), .A3(new_n753), .A4(new_n810), .ZN(new_n811));
  XOR2_X1   g625(.A(new_n811), .B(KEYINPUT48), .Z(new_n812));
  NAND4_X1  g626(.A1(new_n686), .A2(new_n715), .A3(new_n807), .A4(new_n810), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n812), .B(new_n604), .C1(new_n642), .C2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n715), .A2(new_n717), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n816), .B1(new_n805), .B2(new_n808), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(new_n610), .A3(new_n704), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n815), .B1(new_n818), .B2(new_n680), .ZN(new_n819));
  AOI211_X1 g633(.A(new_n703), .B(new_n816), .C1(new_n805), .C2(new_n808), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n678), .B(KEYINPUT38), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(KEYINPUT50), .A3(new_n610), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  OR3_X1    g637(.A1(new_n813), .A2(new_n501), .A3(new_n641), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n796), .A2(new_n799), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n702), .A2(new_n383), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n800), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n825), .B1(new_n828), .B2(new_n817), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT51), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n809), .A2(new_n810), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n832), .A2(new_n720), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n829), .A2(new_n830), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n780), .A2(new_n798), .A3(new_n382), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n798), .B1(new_n780), .B2(new_n382), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n827), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n731), .A3(new_n817), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(new_n833), .A3(new_n823), .A4(new_n824), .ZN(new_n839));
  NAND2_X1  g653(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n830), .A2(new_n831), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n814), .B1(new_n834), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n711), .A2(new_n693), .ZN(new_n844));
  INV_X1    g658(.A(new_n687), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n738), .A2(new_n670), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n685), .A2(new_n844), .A3(new_n845), .A4(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n674), .A2(new_n700), .A3(new_n724), .A4(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n730), .A2(new_n664), .A3(new_n459), .A4(new_n630), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n852), .B1(new_n673), .B2(new_n699), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(KEYINPUT52), .A3(new_n724), .A4(new_n848), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n713), .A2(new_n709), .A3(new_n705), .A4(new_n718), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n749), .B2(new_n760), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n642), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n616), .A2(KEYINPUT116), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n784), .A2(new_n537), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n614), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT116), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n863), .B1(new_n614), .B2(new_n642), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n860), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n629), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n537), .B1(G475), .B2(new_n499), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n731), .A2(new_n671), .A3(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n730), .A2(new_n868), .A3(new_n664), .A4(new_n459), .ZN(new_n869));
  AND4_X1   g683(.A1(new_n618), .A2(new_n866), .A3(new_n665), .A4(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n746), .A2(new_n723), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n870), .A2(new_n871), .A3(new_n763), .A4(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n866), .A2(new_n618), .A3(new_n665), .A4(new_n869), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n763), .A2(new_n872), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT118), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n873), .A2(KEYINPUT53), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n874), .A2(new_n875), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n855), .A2(new_n857), .A3(new_n878), .ZN(new_n879));
  XNOR2_X1  g693(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n858), .A2(new_n877), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n858), .A2(new_n878), .A3(new_n881), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n879), .A2(KEYINPUT53), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n885), .A2(KEYINPUT54), .A3(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n820), .A2(new_n630), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n843), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  OR2_X1    g704(.A1(G952), .A2(G953), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT49), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n702), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n702), .A2(new_n893), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n894), .A2(new_n895), .A3(new_n785), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n685), .A2(new_n260), .A3(new_n383), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n821), .A2(new_n896), .A3(new_n609), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n892), .A2(new_n898), .ZN(G75));
  NOR2_X1   g713(.A1(new_n191), .A2(G952), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n592), .B(new_n581), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT55), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n879), .A2(new_n881), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT53), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n878), .B2(new_n871), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n905), .A2(new_n855), .A3(new_n857), .A4(new_n876), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n907), .A2(G210), .A3(G902), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n902), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n902), .B(KEYINPUT121), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n908), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT122), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n908), .A2(new_n914), .A3(new_n909), .A4(new_n911), .ZN(new_n915));
  AOI211_X1 g729(.A(new_n900), .B(new_n910), .C1(new_n913), .C2(new_n915), .ZN(G51));
  OAI21_X1  g730(.A(KEYINPUT123), .B1(new_n882), .B2(new_n883), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n907), .A2(new_n918), .A3(KEYINPUT54), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n884), .A3(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n385), .B(KEYINPUT57), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n436), .A2(new_n450), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n882), .A2(new_n188), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n778), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n900), .B1(new_n924), .B2(new_n926), .ZN(G54));
  NAND3_X1  g741(.A1(new_n925), .A2(KEYINPUT58), .A3(G475), .ZN(new_n928));
  INV_X1    g742(.A(new_n490), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n930), .A2(new_n931), .A3(new_n900), .ZN(G60));
  INV_X1    g746(.A(new_n900), .ZN(new_n933));
  NAND2_X1  g747(.A1(G478), .A2(G902), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT59), .Z(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n884), .B2(new_n887), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n933), .B1(new_n936), .B2(new_n637), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n634), .B2(new_n636), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n937), .B1(new_n920), .B2(new_n938), .ZN(G63));
  XNOR2_X1  g753(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n187), .A2(new_n188), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n907), .A2(new_n658), .A3(new_n942), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n907), .A2(new_n942), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n933), .B(new_n943), .C1(new_n944), .C2(new_n258), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT61), .B1(new_n943), .B2(KEYINPUT125), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(G66));
  OAI21_X1  g761(.A(G953), .B1(new_n598), .B2(new_n545), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n866), .A2(new_n618), .A3(new_n665), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n856), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n948), .B1(new_n950), .B2(G953), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n586), .B(new_n570), .C1(G898), .C2(new_n191), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(G69));
  AND4_X1   g767(.A1(new_n724), .A2(new_n761), .A3(new_n763), .A4(new_n853), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n781), .A2(new_n715), .A3(new_n753), .A4(new_n844), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n954), .A2(new_n793), .A3(new_n802), .A4(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n346), .A2(new_n347), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(G953), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT62), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n853), .A2(new_n724), .ZN(new_n963));
  OR3_X1    g777(.A1(new_n696), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n962), .B1(new_n696), .B2(new_n963), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n800), .A2(new_n690), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n861), .A2(new_n642), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n378), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(KEYINPUT126), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n969), .A2(KEYINPUT126), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n802), .A2(new_n793), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n966), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n961), .B1(new_n973), .B2(new_n960), .ZN(new_n974));
  OAI21_X1  g788(.A(G900), .B1(new_n960), .B2(G227), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n959), .A2(new_n387), .ZN(new_n976));
  OAI21_X1  g790(.A(G953), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n974), .A2(new_n977), .ZN(G72));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT63), .Z(new_n980));
  INV_X1    g794(.A(new_n950), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n980), .B1(new_n956), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n372), .A2(new_n351), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n980), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n983), .A2(new_n683), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n885), .A2(new_n886), .A3(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n984), .A2(new_n933), .A3(new_n987), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n966), .A2(new_n950), .A3(new_n970), .A4(new_n972), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n980), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT127), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n988), .B1(new_n991), .B2(new_n683), .ZN(G57));
endmodule


