//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1277, new_n1278,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n207), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n202), .A2(G50), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n210), .B1(new_n220), .B2(KEYINPUT1), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n220), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT64), .Z(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G68), .Z(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  NAND2_X1  g0044(.A1(G33), .A2(G41), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n245), .A2(G1), .A3(G13), .ZN(new_n246));
  INV_X1    g0046(.A(G41), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(KEYINPUT5), .ZN(new_n248));
  INV_X1    g0048(.A(G1), .ZN(new_n249));
  OAI211_X1 g0049(.A(new_n249), .B(G45), .C1(new_n247), .C2(KEYINPUT5), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n248), .B1(new_n250), .B2(KEYINPUT83), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT83), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G1), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT5), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G41), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n252), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  OAI211_X1 g0057(.A(G270), .B(new_n246), .C1(new_n251), .C2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT86), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n250), .A2(KEYINPUT83), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n254), .A2(new_n252), .A3(new_n256), .ZN(new_n261));
  INV_X1    g0061(.A(G274), .ZN(new_n262));
  AND2_X1   g0062(.A1(G1), .A2(G13), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n262), .B1(new_n263), .B2(new_n245), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n260), .A2(new_n261), .A3(new_n248), .A4(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n260), .A2(new_n248), .A3(new_n261), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT86), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n266), .A2(new_n267), .A3(G270), .A4(new_n246), .ZN(new_n268));
  AND3_X1   g0068(.A1(new_n259), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G179), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT3), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G33), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n272), .A2(new_n274), .A3(G264), .A4(G1698), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n272), .A2(new_n274), .A3(G257), .A4(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G303), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n275), .B(new_n277), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n246), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n270), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G13), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G1), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G116), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G20), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G283), .ZN(new_n289));
  INV_X1    g0089(.A(G97), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n289), .B(new_n222), .C1(G33), .C2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n221), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n291), .A2(new_n293), .A3(new_n287), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n291), .A2(KEYINPUT20), .A3(new_n293), .A4(new_n287), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n288), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n292), .A2(new_n221), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n284), .A2(G20), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT71), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n283), .A2(new_n222), .A3(G1), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(new_n293), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT71), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n271), .A2(G1), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(new_n286), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n303), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n298), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n269), .A2(new_n282), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n280), .A2(new_n281), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n259), .A2(new_n265), .A3(new_n268), .A4(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G200), .ZN(new_n314));
  INV_X1    g0114(.A(new_n310), .ZN(new_n315));
  INV_X1    g0115(.A(G190), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n314), .B(new_n315), .C1(new_n316), .C2(new_n313), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n318), .B1(new_n298), .B2(new_n309), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT87), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT21), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT21), .ZN(new_n323));
  AOI211_X1 g0123(.A(KEYINPUT87), .B(new_n323), .C1(new_n313), .C2(new_n319), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n311), .B(new_n317), .C1(new_n322), .C2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n279), .A2(G222), .A3(new_n276), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT68), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n279), .A2(G1698), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n272), .A2(new_n274), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n330), .A2(G223), .B1(G77), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n281), .ZN(new_n334));
  INV_X1    g0134(.A(G226), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT66), .ZN(new_n336));
  NOR2_X1   g0136(.A1(G41), .A2(G45), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(G1), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n249), .B(KEYINPUT66), .C1(G41), .C2(G45), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(new_n246), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT67), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n249), .B1(G41), .B2(G45), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n343), .A2(new_n336), .B1(new_n263), .B2(new_n245), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(KEYINPUT67), .A3(new_n339), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n335), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n343), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n264), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n334), .A2(G190), .A3(new_n347), .A4(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT8), .B(G58), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n222), .A2(G33), .ZN(new_n352));
  INV_X1    g0152(.A(G150), .ZN(new_n353));
  NOR2_X1   g0153(.A1(G20), .A2(G33), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n351), .A2(new_n352), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G50), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n222), .B1(new_n201), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n293), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n249), .A2(G20), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n305), .A2(G50), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n304), .A2(new_n357), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT69), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(G50), .ZN(new_n364));
  OAI211_X1 g0164(.A(KEYINPUT69), .B(new_n362), .C1(new_n301), .C2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n359), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT9), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n349), .ZN(new_n370));
  AOI211_X1 g0170(.A(new_n370), .B(new_n346), .C1(new_n333), .C2(new_n281), .ZN(new_n371));
  INV_X1    g0171(.A(G200), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n350), .B(new_n369), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(KEYINPUT9), .B(new_n359), .C1(new_n363), .C2(new_n366), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT72), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n374), .B(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT10), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT10), .B1(new_n367), .B2(new_n368), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n350), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT73), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n371), .B2(new_n372), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n334), .A2(new_n347), .A3(new_n349), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n382), .A2(KEYINPUT73), .A3(G200), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n374), .B(KEYINPUT72), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n379), .A2(new_n381), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n377), .A2(new_n385), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n371), .A2(KEYINPUT70), .A3(new_n270), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT70), .B1(new_n371), .B2(new_n270), .ZN(new_n388));
  OAI221_X1 g0188(.A(new_n367), .B1(G169), .B2(new_n371), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n300), .A2(G68), .B1(KEYINPUT75), .B2(KEYINPUT12), .ZN(new_n391));
  NAND2_X1  g0191(.A1(KEYINPUT75), .A2(KEYINPUT12), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G77), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n352), .A2(new_n394), .B1(new_n222), .B2(G68), .ZN(new_n395));
  OAI22_X1  g0195(.A1(new_n395), .A2(KEYINPUT74), .B1(new_n357), .B2(new_n355), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n395), .A2(KEYINPUT74), .ZN(new_n397));
  OAI211_X1 g0197(.A(KEYINPUT11), .B(new_n293), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n303), .A2(new_n306), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n360), .A2(G68), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n393), .B(new_n398), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  OR2_X1    g0201(.A1(new_n396), .A2(new_n397), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT11), .B1(new_n402), .B2(new_n293), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT14), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT67), .B1(new_n344), .B2(new_n339), .ZN(new_n407));
  AND4_X1   g0207(.A1(KEYINPUT67), .A2(new_n338), .A3(new_n246), .A4(new_n339), .ZN(new_n408));
  OAI21_X1  g0208(.A(G238), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n279), .A2(G232), .A3(G1698), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G97), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n272), .A2(new_n274), .A3(G226), .A4(new_n276), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n370), .B1(new_n413), .B2(new_n281), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT13), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n409), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n415), .B1(new_n409), .B2(new_n414), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n406), .B(G169), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n413), .A2(new_n281), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n349), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n213), .B1(new_n342), .B2(new_n345), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT13), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n409), .A2(new_n414), .A3(new_n415), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(G179), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n422), .A2(new_n423), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n406), .B1(new_n426), .B2(G169), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n405), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n372), .B1(new_n422), .B2(new_n423), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n422), .A2(G190), .A3(new_n423), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n430), .A2(new_n404), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n279), .A2(G232), .A3(new_n276), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n331), .A2(G107), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n433), .B(new_n434), .C1(new_n329), .C2(new_n213), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n370), .B1(new_n435), .B2(new_n281), .ZN(new_n436));
  OAI21_X1  g0236(.A(G244), .B1(new_n407), .B2(new_n408), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(G200), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n436), .A2(new_n437), .A3(G190), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n394), .B1(new_n249), .B2(G20), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n303), .A2(new_n306), .A3(new_n441), .ZN(new_n442));
  OAI22_X1  g0242(.A1(new_n351), .A2(new_n355), .B1(new_n222), .B2(new_n394), .ZN(new_n443));
  XNOR2_X1  g0243(.A(KEYINPUT15), .B(G87), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(new_n352), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n293), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n304), .A2(new_n394), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n442), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n439), .A2(new_n440), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n448), .B1(new_n438), .B2(new_n318), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n436), .A2(new_n437), .A3(new_n270), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n428), .A2(new_n432), .A3(new_n449), .A4(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n390), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n351), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n360), .ZN(new_n456));
  OAI22_X1  g0256(.A1(new_n456), .A2(new_n301), .B1(new_n300), .B2(new_n455), .ZN(new_n457));
  INV_X1    g0257(.A(G58), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(new_n212), .ZN(new_n459));
  OAI21_X1  g0259(.A(G20), .B1(new_n459), .B2(new_n201), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n354), .A2(G159), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT7), .B1(new_n331), .B2(new_n222), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT7), .ZN(new_n464));
  AOI211_X1 g0264(.A(new_n464), .B(G20), .C1(new_n272), .C2(new_n274), .ZN(new_n465));
  OAI21_X1  g0265(.A(G68), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT76), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n464), .B1(new_n279), .B2(G20), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n331), .A2(KEYINPUT7), .A3(new_n222), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n212), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT76), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n462), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n299), .B1(new_n473), .B2(KEYINPUT16), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT16), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(new_n471), .B2(new_n462), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT77), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(KEYINPUT77), .B(new_n475), .C1(new_n471), .C2(new_n462), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n457), .B1(new_n474), .B2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n272), .A2(new_n274), .A3(G226), .A4(G1698), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n272), .A2(new_n274), .A3(G223), .A4(new_n276), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n482), .B(new_n483), .C1(new_n271), .C2(new_n214), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n281), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n338), .A2(G232), .A3(new_n246), .A4(new_n339), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n486), .A2(new_n349), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n318), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n485), .A2(new_n487), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n488), .B1(G179), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT18), .B1(new_n481), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n485), .A2(new_n487), .A3(new_n316), .ZN(new_n492));
  OAI211_X1 g0292(.A(KEYINPUT78), .B(new_n492), .C1(new_n489), .C2(G200), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT78), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n485), .A2(new_n487), .A3(new_n316), .ZN(new_n495));
  AOI21_X1  g0295(.A(G200), .B1(new_n485), .B2(new_n487), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n457), .ZN(new_n499));
  INV_X1    g0299(.A(new_n462), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n471), .A2(KEYINPUT76), .ZN(new_n501));
  AOI211_X1 g0301(.A(new_n467), .B(new_n212), .C1(new_n469), .C2(new_n470), .ZN(new_n502));
  OAI211_X1 g0302(.A(KEYINPUT16), .B(new_n500), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n503), .A2(new_n293), .A3(new_n478), .A4(new_n479), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n498), .A2(new_n499), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT17), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n490), .B1(new_n504), .B2(new_n499), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT18), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n498), .A2(KEYINPUT17), .A3(new_n504), .A4(new_n499), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n491), .A2(new_n507), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT79), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n507), .A2(new_n511), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  XNOR2_X1  g0316(.A(new_n508), .B(KEYINPUT18), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT79), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n454), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n272), .A2(new_n274), .A3(G257), .A4(G1698), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n272), .A2(new_n274), .A3(G250), .A4(new_n276), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G294), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n281), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n265), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT89), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n266), .A2(new_n527), .A3(G264), .A4(new_n246), .ZN(new_n528));
  OAI211_X1 g0328(.A(G264), .B(new_n246), .C1(new_n251), .C2(new_n257), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT89), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n526), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT90), .B1(new_n531), .B2(new_n318), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n528), .ZN(new_n533));
  INV_X1    g0333(.A(new_n526), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT90), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n535), .A2(new_n536), .A3(G169), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n531), .A2(G179), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n532), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n272), .A2(new_n274), .A3(new_n222), .A4(G87), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT22), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT22), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n279), .A2(new_n542), .A3(new_n222), .A4(G87), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g0344(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G116), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n546), .A2(G20), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT23), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n222), .B2(G107), .ZN(new_n549));
  INV_X1    g0349(.A(G107), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n550), .A2(KEYINPUT23), .A3(G20), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n547), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n544), .A2(new_n545), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n545), .B1(new_n544), .B2(new_n552), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n293), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n301), .A2(new_n307), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT25), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n300), .B2(G107), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n304), .A2(KEYINPUT25), .A3(new_n550), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n556), .A2(G107), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n533), .A2(new_n534), .A3(G190), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n562), .A2(new_n555), .A3(new_n560), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n531), .A2(new_n372), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n539), .A2(new_n561), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(G257), .B(new_n246), .C1(new_n251), .C2(new_n257), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n568), .A2(new_n265), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n272), .A2(new_n274), .A3(G244), .A4(new_n276), .ZN(new_n570));
  XOR2_X1   g0370(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n279), .A2(KEYINPUT4), .A3(G244), .A4(new_n276), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n279), .A2(G250), .A3(G1698), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n289), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n281), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n318), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n569), .A2(new_n270), .A3(new_n576), .ZN(new_n579));
  AND2_X1   g0379(.A1(G97), .A2(G107), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT80), .ZN(new_n581));
  OAI22_X1  g0381(.A1(new_n580), .A2(new_n204), .B1(new_n581), .B2(KEYINPUT6), .ZN(new_n582));
  MUX2_X1   g0382(.A(new_n581), .B(G97), .S(KEYINPUT6), .Z(new_n583));
  XNOR2_X1  g0383(.A(G97), .B(G107), .ZN(new_n584));
  OAI211_X1 g0384(.A(G20), .B(new_n582), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n354), .A2(G77), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n469), .A2(new_n470), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n587), .A2(KEYINPUT81), .B1(G107), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT81), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n585), .A2(new_n590), .A3(new_n586), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n299), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n300), .A2(G97), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n556), .B2(G97), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n578), .B(new_n579), .C1(new_n592), .C2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n587), .A2(KEYINPUT81), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n588), .A2(G107), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n591), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n293), .ZN(new_n600));
  INV_X1    g0400(.A(new_n576), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n568), .A2(new_n265), .ZN(new_n602));
  OAI21_X1  g0402(.A(G200), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n569), .A2(G190), .A3(new_n576), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n600), .A2(new_n603), .A3(new_n594), .A4(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n279), .A2(new_n222), .A3(G68), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT19), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n222), .B1(new_n411), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(G87), .B2(new_n205), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n607), .B1(new_n352), .B2(new_n290), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n606), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n611), .A2(new_n293), .B1(new_n304), .B2(new_n444), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n556), .A2(G87), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n272), .A2(new_n274), .A3(G244), .A4(G1698), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n272), .A2(new_n274), .A3(G238), .A4(new_n276), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n616), .A3(new_n546), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n281), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n215), .B1(new_n253), .B2(G1), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n249), .A2(new_n262), .A3(G45), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n246), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT84), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n246), .A2(new_n619), .A3(new_n620), .A4(KEYINPUT84), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n618), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(G200), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n281), .A2(new_n617), .B1(new_n623), .B2(new_n624), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(G190), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n614), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT85), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n618), .A2(G179), .A3(new_n625), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n318), .B1(new_n618), .B2(new_n625), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n626), .A2(G169), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n628), .A2(G179), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n636), .A3(KEYINPUT85), .ZN(new_n637));
  INV_X1    g0437(.A(new_n556), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n612), .B1(new_n638), .B2(new_n444), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n634), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  AND4_X1   g0440(.A1(new_n596), .A2(new_n605), .A3(new_n630), .A4(new_n640), .ZN(new_n641));
  AND4_X1   g0441(.A1(new_n326), .A2(new_n520), .A3(new_n567), .A4(new_n641), .ZN(G372));
  NAND2_X1  g0442(.A1(new_n431), .A2(new_n404), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(new_n429), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n428), .B1(new_n644), .B2(new_n452), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n516), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n491), .A2(new_n510), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n386), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n389), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n596), .A2(KEYINPUT92), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n600), .A2(new_n594), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT92), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n652), .A2(new_n653), .A3(new_n578), .A4(new_n579), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n635), .A2(new_n636), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n639), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n630), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n651), .A2(new_n654), .A3(new_n655), .A4(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n640), .A2(new_n630), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT26), .B1(new_n660), .B2(new_n596), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n659), .A2(new_n657), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n311), .B1(new_n322), .B2(new_n324), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT91), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT91), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n665), .B(new_n311), .C1(new_n322), .C2(new_n324), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n539), .A2(new_n561), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n563), .A2(new_n565), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n630), .A2(new_n657), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n596), .A2(new_n605), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n662), .B1(new_n669), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n650), .B1(new_n519), .B2(new_n676), .ZN(G369));
  OR3_X1    g0477(.A1(new_n285), .A2(KEYINPUT27), .A3(G20), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT27), .B1(new_n285), .B2(G20), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n668), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n682), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n668), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT93), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n684), .B1(new_n555), .B2(new_n560), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n687), .B1(new_n567), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n561), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n318), .B1(new_n533), .B2(new_n534), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n692), .A2(new_n536), .B1(G179), .B2(new_n531), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n691), .B1(new_n693), .B2(new_n532), .ZN(new_n694));
  NOR4_X1   g0494(.A1(new_n694), .A2(KEYINPUT93), .A3(new_n670), .A4(new_n688), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n686), .B1(new_n690), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT94), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n670), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n668), .A2(new_n699), .A3(new_n689), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT93), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n567), .A2(new_n687), .A3(new_n689), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(KEYINPUT94), .A3(new_n686), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n698), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n663), .A2(new_n684), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT95), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n683), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n315), .A2(new_n684), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n664), .A2(new_n666), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n325), .B2(new_n709), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n711), .A2(G330), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n705), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n708), .A2(new_n713), .ZN(G399));
  INV_X1    g0514(.A(new_n208), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G41), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(G1), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT96), .ZN(new_n720));
  OAI22_X1  g0520(.A1(new_n719), .A2(new_n720), .B1(new_n225), .B2(new_n717), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n721), .B1(new_n720), .B2(new_n719), .ZN(new_n722));
  XOR2_X1   g0522(.A(new_n722), .B(KEYINPUT28), .Z(new_n723));
  AND3_X1   g0523(.A1(new_n659), .A2(new_n657), .A3(new_n661), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n694), .B1(new_n664), .B2(new_n666), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n724), .B1(new_n725), .B2(new_n674), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT29), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n726), .A2(new_n727), .A3(new_n684), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n672), .B(new_n673), .C1(new_n663), .C2(new_n694), .ZN(new_n729));
  INV_X1    g0529(.A(new_n657), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n660), .A2(new_n596), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n730), .B1(new_n731), .B2(new_n655), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n651), .A2(new_n658), .A3(new_n654), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT26), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n729), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n684), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(KEYINPUT29), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n728), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n602), .B1(new_n281), .B2(new_n575), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT98), .B1(new_n531), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT98), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n535), .A2(new_n741), .A3(new_n577), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n628), .A2(G179), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n313), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n740), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n628), .A2(new_n282), .A3(new_n525), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n269), .A2(new_n746), .A3(new_n739), .A4(new_n533), .ZN(new_n747));
  XOR2_X1   g0547(.A(KEYINPUT97), .B(KEYINPUT30), .Z(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n533), .A2(new_n576), .A3(new_n569), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n750), .A2(KEYINPUT30), .A3(new_n269), .A4(new_n746), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n745), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n682), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT31), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n326), .A2(new_n567), .A3(new_n641), .A4(new_n684), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT99), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n745), .A2(new_n757), .A3(new_n749), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n751), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n757), .B1(new_n745), .B2(new_n749), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n682), .A2(KEYINPUT31), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n755), .B(new_n756), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G330), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n738), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n723), .B1(new_n767), .B2(G1), .ZN(G364));
  NOR2_X1   g0568(.A1(new_n283), .A2(G20), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n249), .B1(new_n769), .B2(G45), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n716), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n712), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(G330), .B2(new_n711), .ZN(new_n774));
  INV_X1    g0574(.A(new_n772), .ZN(new_n775));
  NAND3_X1  g0575(.A1(G355), .A2(new_n279), .A3(new_n208), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n243), .A2(new_n253), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n715), .A2(new_n279), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(G45), .B2(new_n225), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n776), .B1(G116), .B2(new_n208), .C1(new_n777), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G13), .A2(G33), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n221), .B1(G20), .B2(new_n318), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n775), .B1(new_n780), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT100), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  INV_X1    g0589(.A(new_n784), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n222), .A2(new_n270), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G200), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n316), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n222), .A2(G190), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n795), .A2(new_n270), .A3(new_n372), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G159), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n794), .A2(new_n357), .B1(new_n798), .B2(KEYINPUT32), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n792), .A2(G190), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n799), .B1(G68), .B2(new_n800), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n316), .A2(G179), .A3(G200), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n222), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n798), .A2(KEYINPUT32), .B1(G97), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G190), .A2(G200), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n791), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n279), .B1(new_n807), .B2(new_n394), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n791), .A2(G190), .A3(new_n372), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n808), .B1(G58), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n805), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n270), .A2(G200), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT101), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n814), .A2(new_n222), .A3(new_n316), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G87), .ZN(new_n816));
  NOR3_X1   g0616(.A1(new_n814), .A2(new_n222), .A3(G190), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G107), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n801), .A2(new_n812), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n800), .ZN(new_n820));
  XNOR2_X1  g0620(.A(KEYINPUT33), .B(G317), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT102), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n822), .B2(new_n821), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G283), .A2(new_n817), .B1(new_n815), .B2(G303), .ZN(new_n825));
  INV_X1    g0625(.A(G311), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n807), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G322), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n331), .B1(new_n809), .B2(new_n828), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n827), .B(new_n829), .C1(G329), .C2(new_n797), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G294), .A2(new_n804), .B1(new_n793), .B2(G326), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n824), .A2(new_n825), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n790), .B1(new_n819), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n789), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n783), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n788), .B(new_n834), .C1(new_n711), .C2(new_n835), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n774), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(G396));
  OR2_X1    g0638(.A1(new_n448), .A2(new_n684), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n449), .A2(new_n839), .B1(new_n450), .B2(new_n451), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n450), .A2(new_n451), .A3(new_n684), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(KEYINPUT105), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n449), .A2(new_n839), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n452), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT105), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n845), .A2(new_n846), .A3(new_n841), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n676), .B2(new_n682), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n682), .B1(new_n843), .B2(new_n847), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n850), .B1(new_n676), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n772), .B1(new_n853), .B2(new_n765), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n765), .B2(new_n853), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n784), .A2(new_n781), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n772), .B1(G77), .B2(new_n857), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT103), .ZN(new_n859));
  INV_X1    g0659(.A(new_n807), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n793), .A2(G303), .B1(new_n860), .B2(G116), .ZN(new_n861));
  INV_X1    g0661(.A(G283), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n861), .B1(new_n862), .B2(new_n820), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT104), .Z(new_n864));
  INV_X1    g0664(.A(G294), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n331), .B1(new_n796), .B2(new_n826), .C1(new_n809), .C2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(G97), .B2(new_n804), .ZN(new_n867));
  AOI22_X1  g0667(.A1(G87), .A2(new_n817), .B1(new_n815), .B2(G107), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n864), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n810), .A2(G143), .B1(new_n860), .B2(G159), .ZN(new_n870));
  INV_X1    g0670(.A(G137), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n870), .B1(new_n794), .B2(new_n871), .C1(new_n353), .C2(new_n820), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT34), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n873), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n817), .A2(G68), .ZN(new_n876));
  INV_X1    g0676(.A(G132), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n279), .B1(new_n796), .B2(new_n877), .C1(new_n803), .C2(new_n458), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(G50), .B2(new_n815), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n874), .A2(new_n875), .A3(new_n876), .A4(new_n879), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n869), .A2(new_n880), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n859), .B1(new_n790), .B2(new_n881), .C1(new_n848), .C2(new_n782), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n855), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(G384));
  OAI21_X1  g0684(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n885), .B(KEYINPUT106), .Z(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT35), .ZN(new_n888));
  OAI211_X1 g0688(.A(G116), .B(new_n223), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n888), .B2(new_n887), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n890), .B(KEYINPUT36), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n225), .A2(new_n394), .A3(new_n459), .ZN(new_n892));
  OR2_X1    g0692(.A1(new_n892), .A2(KEYINPUT107), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n892), .A2(KEYINPUT107), .B1(new_n357), .B2(G68), .ZN(new_n894));
  AOI211_X1 g0694(.A(new_n249), .B(G13), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n475), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n457), .B1(new_n474), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n505), .B1(new_n899), .B2(new_n680), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n899), .A2(new_n490), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT37), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n508), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n504), .A2(new_n499), .ZN(new_n904));
  INV_X1    g0704(.A(new_n680), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n903), .A2(new_n906), .A3(new_n907), .A4(new_n505), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n899), .A2(new_n680), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n512), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n909), .A2(new_n911), .A3(KEYINPUT38), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n903), .A2(new_n906), .A3(new_n505), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT37), .ZN(new_n914));
  INV_X1    g0714(.A(new_n906), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n908), .A2(new_n914), .B1(new_n512), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n912), .B1(new_n916), .B2(KEYINPUT38), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT39), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n909), .A2(new_n911), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT38), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(KEYINPUT39), .A3(new_n912), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(G169), .B1(new_n416), .B2(new_n417), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT14), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(new_n424), .A3(new_n418), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(new_n405), .A3(new_n684), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n925), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n842), .B1(new_n726), .B2(new_n851), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n405), .B(new_n682), .C1(new_n928), .C2(new_n644), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n405), .A2(new_n682), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n428), .A2(new_n432), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n909), .A2(new_n911), .A3(KEYINPUT38), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT38), .B1(new_n909), .B2(new_n911), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n933), .B(new_n937), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n647), .A2(new_n680), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n931), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n519), .B1(new_n728), .B2(new_n737), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n943), .A2(new_n649), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n942), .B(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(G330), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n752), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n756), .A2(new_n755), .A3(new_n947), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n934), .A2(new_n936), .B1(new_n847), .B2(new_n843), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n938), .B2(new_n939), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT40), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n948), .A2(new_n949), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT108), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT108), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n948), .A2(new_n949), .A3(new_n956), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n917), .A2(new_n955), .A3(KEYINPUT40), .A4(new_n957), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n520), .A2(new_n948), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n946), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n959), .B2(new_n960), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n945), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n249), .B2(new_n769), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n945), .A2(new_n962), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n896), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT109), .ZN(G367));
  INV_X1    g0767(.A(new_n652), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n673), .B1(new_n968), .B2(new_n684), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n596), .A2(new_n684), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n705), .A2(new_n707), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n596), .B1(new_n969), .B2(new_n668), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n972), .A2(KEYINPUT42), .B1(new_n684), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(KEYINPUT42), .B2(new_n972), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n614), .A2(new_n684), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n730), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n671), .B2(new_n976), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n971), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n713), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(KEYINPUT110), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT110), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n982), .A2(new_n986), .ZN(new_n987));
  AND3_X1   g0787(.A1(new_n984), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n985), .B1(new_n984), .B2(new_n987), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n980), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n984), .A2(new_n987), .ZN(new_n991));
  INV_X1    g0791(.A(new_n985), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n975), .A2(new_n979), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n984), .A2(new_n985), .A3(new_n987), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  AND2_X1   g0796(.A1(new_n990), .A2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n716), .B(KEYINPUT41), .Z(new_n998));
  INV_X1    g0798(.A(KEYINPUT44), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n708), .B2(new_n971), .ZN(new_n1000));
  AOI21_X1  g0800(.A(KEYINPUT94), .B1(new_n703), .B2(new_n686), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n697), .B(new_n685), .C1(new_n701), .C2(new_n702), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n707), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n683), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1005), .A2(KEYINPUT44), .A3(new_n981), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1000), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1003), .A2(new_n1004), .A3(new_n971), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT45), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n708), .A2(KEYINPUT45), .A3(new_n971), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n713), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1007), .A2(new_n1012), .A3(new_n713), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n705), .A2(new_n712), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1017), .A2(new_n713), .A3(new_n707), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n707), .B1(new_n1017), .B2(new_n713), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n1019), .A2(new_n1020), .A3(new_n766), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1015), .A2(new_n1016), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n998), .B1(new_n1022), .B2(new_n767), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n997), .B1(new_n1023), .B2(new_n771), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n785), .B1(new_n208), .B2(new_n444), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n236), .B2(new_n778), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n803), .A2(new_n212), .ZN(new_n1027));
  INV_X1    g0827(.A(G143), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n794), .A2(new_n1028), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1027), .B(new_n1029), .C1(G159), .C2(new_n800), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n815), .A2(G58), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n817), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1032), .A2(new_n394), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n809), .A2(new_n353), .B1(new_n807), .B2(new_n357), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n331), .B(new_n1035), .C1(G137), .C2(new_n797), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1030), .A2(new_n1031), .A3(new_n1034), .A4(new_n1036), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n794), .A2(new_n826), .B1(new_n550), .B2(new_n803), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(G294), .B2(new_n800), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n817), .A2(G97), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n279), .B1(new_n860), .B2(G283), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G303), .A2(new_n810), .B1(new_n797), .B2(G317), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n815), .A2(G116), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT46), .Z(new_n1045));
  OAI21_X1  g0845(.A(new_n1037), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT47), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n775), .B(new_n1026), .C1(new_n1047), .C2(new_n784), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n978), .A2(new_n835), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1024), .A2(new_n1050), .ZN(G387));
  NOR2_X1   g0851(.A1(new_n1021), .A2(new_n717), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1052), .B1(new_n767), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n778), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n233), .A2(G45), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT111), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n351), .A2(G50), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT50), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n718), .ZN(new_n1060));
  AOI211_X1 g0860(.A(G45), .B(new_n1060), .C1(G68), .C2(G77), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1055), .B(new_n1057), .C1(new_n1059), .C2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n279), .A2(new_n208), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n718), .A2(new_n1063), .B1(G107), .B2(new_n208), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n785), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n772), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n705), .A2(new_n835), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n279), .B1(new_n807), .B2(new_n212), .ZN(new_n1068));
  INV_X1    g0868(.A(G159), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n1069), .A2(new_n794), .B1(new_n820), .B2(new_n351), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1068), .B(new_n1070), .C1(G150), .C2(new_n797), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n815), .A2(G77), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n803), .A2(new_n444), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(G50), .B2(new_n810), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT112), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1071), .A2(new_n1040), .A3(new_n1072), .A4(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n279), .B1(new_n797), .B2(G326), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n815), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n1078), .A2(new_n865), .B1(new_n862), .B2(new_n803), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n810), .A2(G317), .B1(new_n860), .B2(G303), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1080), .B1(new_n794), .B2(new_n828), .C1(new_n826), .C2(new_n820), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT48), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n1082), .B2(new_n1081), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT49), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1077), .B1(new_n286), .B2(new_n1032), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1076), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1066), .B(new_n1067), .C1(new_n784), .C2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n1053), .B2(new_n771), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1054), .A2(new_n1090), .ZN(G393));
  INV_X1    g0891(.A(new_n1020), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1092), .A2(new_n1018), .A3(new_n767), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n1007), .A2(new_n1012), .A3(new_n713), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n713), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1096), .A2(new_n1022), .A3(new_n716), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n981), .A2(new_n783), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n785), .B1(new_n290), .B2(new_n208), .C1(new_n240), .C2(new_n1055), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n772), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n820), .A2(new_n357), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n279), .B1(new_n807), .B2(new_n351), .C1(new_n1028), .C2(new_n796), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n803), .A2(new_n394), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1105), .B1(new_n212), .B2(new_n1078), .C1(new_n214), .C2(new_n1032), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G150), .A2(new_n793), .B1(new_n810), .B2(G159), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1107), .B(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n815), .A2(G283), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n331), .B1(new_n807), .B2(new_n865), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(G322), .B2(new_n797), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G116), .A2(new_n804), .B1(new_n800), .B2(G303), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n818), .A2(new_n1110), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G317), .A2(new_n793), .B1(new_n810), .B2(G311), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT52), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n1106), .A2(new_n1109), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1101), .B1(new_n1117), .B2(new_n784), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1098), .A2(new_n771), .B1(new_n1099), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1097), .A2(new_n1119), .ZN(G390));
  INV_X1    g0920(.A(new_n937), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n929), .B1(new_n932), .B2(new_n1121), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n914), .A2(new_n908), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n906), .B1(new_n516), .B2(new_n517), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n921), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(KEYINPUT39), .B1(new_n1125), .B2(new_n912), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n938), .A2(new_n939), .A3(new_n918), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1122), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n930), .B1(new_n1125), .B2(new_n912), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n735), .A2(new_n684), .A3(new_n848), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n841), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n937), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n764), .A2(G330), .A3(new_n848), .A4(new_n937), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1128), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n924), .A2(new_n1122), .B1(new_n1132), .B2(new_n1129), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n948), .A2(G330), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n949), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1135), .B(new_n771), .C1(new_n1136), .C2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n772), .B1(new_n455), .B2(new_n857), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n279), .B1(new_n809), .B2(new_n877), .ZN(new_n1142));
  INV_X1    g0942(.A(G128), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n794), .A2(new_n1143), .B1(new_n1069), .B2(new_n803), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1142), .B(new_n1144), .C1(G125), .C2(new_n797), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT54), .B(G143), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n800), .A2(G137), .B1(new_n860), .B2(new_n1147), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT114), .Z(new_n1149));
  OAI211_X1 g0949(.A(new_n1145), .B(new_n1149), .C1(new_n357), .C2(new_n1032), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n815), .A2(G150), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT53), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1104), .B1(G283), .B2(new_n793), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n550), .B2(new_n820), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n809), .A2(new_n286), .B1(new_n807), .B2(new_n290), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n279), .B(new_n1155), .C1(G294), .C2(new_n797), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1156), .A2(new_n816), .A3(new_n876), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n1150), .A2(new_n1152), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1141), .B1(new_n1158), .B2(new_n784), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n925), .B2(new_n782), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1140), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT115), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1140), .A2(KEYINPUT115), .A3(new_n1160), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1139), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n1136), .B2(new_n1134), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1121), .B1(new_n1137), .B2(new_n849), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1168), .A2(new_n1134), .A3(new_n841), .A4(new_n1130), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n756), .A2(new_n755), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n761), .A2(new_n760), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n763), .B1(new_n1171), .B2(new_n758), .ZN(new_n1172));
  OAI211_X1 g0972(.A(G330), .B(new_n848), .C1(new_n1170), .C2(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n949), .A2(new_n1138), .B1(new_n1173), .B2(new_n1121), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1169), .B1(new_n1174), .B2(new_n932), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n519), .A2(new_n1137), .ZN(new_n1176));
  NOR3_X1   g0976(.A1(new_n943), .A2(new_n649), .A3(new_n1176), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n717), .B1(new_n1167), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1135), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1165), .A2(new_n1183), .ZN(G378));
  AOI21_X1  g0984(.A(new_n954), .B1(new_n922), .B2(new_n912), .ZN(new_n1185));
  OAI21_X1  g0985(.A(G330), .B1(new_n1185), .B2(KEYINPUT40), .ZN(new_n1186));
  AND4_X1   g0986(.A1(KEYINPUT40), .A2(new_n917), .A3(new_n955), .A4(new_n957), .ZN(new_n1187));
  OAI21_X1  g0987(.A(KEYINPUT119), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT119), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n953), .A2(new_n958), .A3(new_n1189), .A4(G330), .ZN(new_n1190));
  XOR2_X1   g0990(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1191));
  XNOR2_X1  g0991(.A(new_n390), .B(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n367), .A2(new_n905), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT118), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1192), .B(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1188), .A2(new_n1190), .A3(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n931), .A2(new_n940), .A3(new_n941), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1195), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1198), .B(KEYINPUT119), .C1(new_n1187), .C2(new_n1186), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1196), .A2(new_n1197), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1197), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n771), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n775), .B1(new_n357), .B2(new_n856), .ZN(new_n1203));
  AOI21_X1  g1003(.A(G50), .B1(new_n271), .B2(new_n247), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n279), .B2(G41), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1027), .B1(G116), .B2(new_n793), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT116), .Z(new_n1207));
  OAI211_X1 g1007(.A(new_n247), .B(new_n331), .C1(new_n796), .C2(new_n862), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n809), .A2(new_n550), .B1(new_n807), .B2(new_n444), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(G97), .C2(new_n800), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n817), .A2(G58), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1207), .A2(new_n1210), .A3(new_n1072), .A4(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1205), .B1(new_n1213), .B2(KEYINPUT58), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n809), .A2(new_n1143), .B1(new_n807), .B2(new_n871), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G132), .B2(new_n800), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(G150), .A2(new_n804), .B1(new_n793), .B2(G125), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(new_n1078), .C2(new_n1146), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT59), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1219), .A2(KEYINPUT117), .ZN(new_n1220));
  AOI211_X1 g1020(.A(G33), .B(G41), .C1(new_n797), .C2(G124), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n1032), .B2(new_n1069), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n1219), .B2(KEYINPUT117), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1220), .A2(new_n1223), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1214), .B(new_n1224), .C1(KEYINPUT58), .C2(new_n1213), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1203), .B1(new_n790), .B2(new_n1225), .C1(new_n1198), .C2(new_n782), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1202), .A2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1177), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT57), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n717), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1190), .A2(new_n1195), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n946), .B1(new_n951), .B2(new_n952), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1189), .B1(new_n1233), .B2(new_n958), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1189), .B(new_n1195), .C1(new_n1233), .C2(new_n958), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n942), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT120), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1196), .A2(new_n1197), .A3(new_n1199), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1201), .A2(KEYINPUT120), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1178), .B(new_n1135), .C1(new_n1136), .C2(new_n1139), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1230), .B1(new_n1242), .B2(new_n1177), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1240), .A2(new_n1241), .A3(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1227), .B1(new_n1231), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(G375));
  NAND2_X1  g1046(.A1(new_n1175), .A2(new_n771), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1121), .A2(new_n781), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT122), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n775), .B1(new_n212), .B2(new_n856), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n820), .A2(new_n1146), .B1(new_n357), .B2(new_n803), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(G137), .A2(new_n810), .B1(new_n797), .B2(G128), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n1252), .B1(new_n353), .B2(new_n807), .C1(new_n1078), .C2(new_n1069), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1251), .B(new_n1253), .C1(G132), .C2(new_n793), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1211), .A2(new_n279), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1255), .B(KEYINPUT123), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n820), .A2(new_n286), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n1073), .B(new_n1258), .C1(G294), .C2(new_n793), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n279), .B1(new_n860), .B2(G107), .ZN(new_n1260));
  OAI221_X1 g1060(.A(new_n1260), .B1(new_n862), .B2(new_n809), .C1(new_n278), .C2(new_n796), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n1261), .B(new_n1033), .C1(G97), .C2(new_n815), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1254), .A2(new_n1257), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1249), .B(new_n1250), .C1(new_n790), .C2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1247), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  OR2_X1    g1066(.A1(new_n1174), .A2(new_n932), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1176), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1268), .B(new_n650), .C1(new_n738), .C2(new_n519), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT121), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1267), .A2(new_n1269), .A3(new_n1270), .A4(new_n1169), .ZN(new_n1271));
  OAI21_X1  g1071(.A(KEYINPUT121), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n998), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1181), .A2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1266), .B1(new_n1273), .B2(new_n1275), .ZN(G381));
  NAND3_X1  g1076(.A1(new_n1054), .A2(new_n837), .A3(new_n1090), .ZN(new_n1277));
  OR4_X1    g1077(.A1(G384), .A2(G390), .A3(new_n1277), .A4(G381), .ZN(new_n1278));
  OR4_X1    g1078(.A1(G387), .A2(new_n1278), .A3(G378), .A4(G375), .ZN(G407));
  AOI22_X1  g1079(.A1(new_n1163), .A2(new_n1164), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n681), .A2(G213), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(KEYINPUT124), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1245), .A2(new_n1280), .A3(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(G407), .A2(G213), .A3(new_n1283), .ZN(G409));
  NAND2_X1  g1084(.A1(new_n1181), .A2(KEYINPUT60), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(new_n1272), .A3(new_n1271), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n717), .B1(new_n1287), .B2(KEYINPUT60), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(G384), .B1(new_n1289), .B2(new_n1266), .ZN(new_n1290));
  AOI211_X1 g1090(.A(new_n1265), .B(new_n883), .C1(new_n1286), .C2(new_n1288), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  AOI211_X1 g1092(.A(new_n1280), .B(new_n1227), .C1(new_n1231), .C2(new_n1244), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1226), .ZN(new_n1294));
  AOI22_X1  g1094(.A1(new_n1237), .A2(new_n1239), .B1(new_n1242), .B2(new_n1177), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1294), .B1(new_n1295), .B2(new_n1274), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1240), .A2(new_n771), .A3(new_n1241), .ZN(new_n1297));
  AOI21_X1  g1097(.A(G378), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1281), .B(new_n1292), .C1(new_n1293), .C2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT62), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1227), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n716), .B1(new_n1295), .B2(KEYINPUT57), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1240), .A2(new_n1241), .A3(new_n1243), .ZN(new_n1303));
  OAI211_X1 g1103(.A(G378), .B(new_n1301), .C1(new_n1302), .C2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1297), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1226), .B1(new_n1229), .B2(new_n998), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1280), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1282), .B1(new_n1304), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1292), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1309), .A2(new_n1300), .ZN(new_n1310));
  AOI22_X1  g1110(.A1(new_n1299), .A2(new_n1300), .B1(new_n1308), .B2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT61), .ZN(new_n1312));
  AND2_X1   g1112(.A1(new_n1282), .A2(G2897), .ZN(new_n1313));
  OAI211_X1 g1113(.A(KEYINPUT125), .B(new_n1313), .C1(new_n1290), .C2(new_n1291), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1281), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(G2897), .ZN(new_n1317));
  AOI21_X1  g1117(.A(KEYINPUT125), .B1(new_n1292), .B2(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1313), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1315), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1312), .B1(new_n1308), .B2(new_n1320), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1024), .A2(new_n1050), .A3(G390), .ZN(new_n1322));
  AOI21_X1  g1122(.A(G390), .B1(new_n1024), .B2(new_n1050), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(G393), .A2(G396), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1277), .ZN(new_n1325));
  NOR3_X1   g1125(.A1(new_n1322), .A2(new_n1323), .A3(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1325), .ZN(new_n1327));
  INV_X1    g1127(.A(G390), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n990), .A2(new_n996), .ZN(new_n1329));
  NOR3_X1   g1129(.A1(new_n1094), .A2(new_n1095), .A3(new_n1093), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1274), .B1(new_n1330), .B2(new_n766), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1329), .B1(new_n1331), .B2(new_n770), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1050), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1328), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1024), .A2(new_n1050), .A3(G390), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1327), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  OAI22_X1  g1136(.A1(new_n1311), .A2(new_n1321), .B1(new_n1326), .B2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT126), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1334), .A2(new_n1327), .A3(new_n1335), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1325), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1316), .B1(new_n1304), .B2(new_n1307), .ZN(new_n1341));
  OAI211_X1 g1141(.A(new_n1339), .B(new_n1340), .C1(new_n1341), .C2(new_n1320), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1282), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT63), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1309), .A2(new_n1344), .ZN(new_n1345));
  OAI211_X1 g1145(.A(new_n1343), .B(new_n1345), .C1(new_n1293), .C2(new_n1298), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(new_n1312), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1342), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1299), .A2(new_n1344), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1338), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1350));
  AOI21_X1  g1150(.A(KEYINPUT61), .B1(new_n1308), .B2(new_n1345), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1326), .A2(new_n1336), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1292), .A2(new_n1317), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT125), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1353), .A2(new_n1354), .A3(new_n1319), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1355), .A2(new_n1314), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1298), .B1(G378), .B2(new_n1245), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1356), .B1(new_n1357), .B2(new_n1316), .ZN(new_n1358));
  NAND4_X1  g1158(.A1(new_n1349), .A2(new_n1351), .A3(new_n1352), .A4(new_n1358), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1359), .A2(KEYINPUT126), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1337), .B1(new_n1350), .B2(new_n1360), .ZN(G405));
  NAND2_X1  g1161(.A1(new_n1309), .A2(KEYINPUT127), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1352), .A2(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(new_n1363), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1352), .A2(new_n1362), .ZN(new_n1365));
  OAI21_X1  g1165(.A(new_n1304), .B1(KEYINPUT127), .B2(new_n1309), .ZN(new_n1366));
  NOR2_X1   g1166(.A1(new_n1245), .A2(G378), .ZN(new_n1367));
  NOR2_X1   g1167(.A1(new_n1366), .A2(new_n1367), .ZN(new_n1368));
  INV_X1    g1168(.A(new_n1368), .ZN(new_n1369));
  NOR3_X1   g1169(.A1(new_n1364), .A2(new_n1365), .A3(new_n1369), .ZN(new_n1370));
  OR2_X1    g1170(.A1(new_n1352), .A2(new_n1362), .ZN(new_n1371));
  AOI21_X1  g1171(.A(new_n1368), .B1(new_n1371), .B2(new_n1363), .ZN(new_n1372));
  NOR2_X1   g1172(.A1(new_n1370), .A2(new_n1372), .ZN(G402));
endmodule


