//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  OR2_X1    g003(.A1(KEYINPUT69), .A2(G116), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT69), .A2(G116), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(G119), .A3(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G116), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT2), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G113), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n195), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT70), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n192), .A2(new_n194), .A3(new_n200), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n195), .A2(KEYINPUT70), .A3(new_n201), .ZN(new_n206));
  INV_X1    g020(.A(G104), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT3), .B1(new_n207), .B2(G107), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G104), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n207), .A2(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n208), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT4), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G101), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(G101), .ZN(new_n216));
  INV_X1    g030(.A(G101), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n208), .A2(new_n211), .A3(new_n217), .A4(new_n212), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(KEYINPUT4), .A3(new_n218), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n205), .A2(new_n206), .A3(new_n215), .A4(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n192), .A2(KEYINPUT5), .A3(new_n194), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n194), .A2(KEYINPUT5), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(new_n196), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT85), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n207), .A2(G107), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n210), .A2(G104), .ZN(new_n228));
  OAI21_X1  g042(.A(G101), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n204), .A2(new_n218), .A3(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n221), .A2(KEYINPUT85), .A3(new_n223), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n226), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(G110), .B(G122), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n220), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G143), .B(G146), .ZN(new_n235));
  AND2_X1   g049(.A1(KEYINPUT0), .A2(G128), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT66), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G146), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G143), .ZN(new_n239));
  INV_X1    g053(.A(G143), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G146), .ZN(new_n241));
  AND4_X1   g055(.A1(KEYINPUT66), .A2(new_n239), .A3(new_n241), .A4(new_n236), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  OR2_X1    g058(.A1(new_n236), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n241), .A2(KEYINPUT65), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n239), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n238), .A2(KEYINPUT65), .A3(G143), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n245), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(G125), .B1(new_n243), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G953), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G224), .ZN(new_n252));
  INV_X1    g066(.A(G125), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n235), .A2(new_n254), .A3(G128), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n238), .A2(KEYINPUT65), .A3(G143), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n256), .B1(new_n246), .B2(new_n239), .ZN(new_n257));
  INV_X1    g071(.A(G128), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n258), .B1(new_n239), .B2(KEYINPUT1), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n253), .B(new_n255), .C1(new_n257), .C2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n250), .A2(KEYINPUT7), .A3(new_n252), .A4(new_n260), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n234), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n233), .B(KEYINPUT8), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n218), .A2(new_n229), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n221), .A2(KEYINPUT85), .A3(new_n223), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT85), .B1(new_n221), .B2(new_n223), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n264), .B1(new_n267), .B2(new_n204), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n224), .A2(new_n264), .A3(new_n204), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT87), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT87), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n230), .A2(new_n271), .A3(new_n224), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n263), .B1(new_n268), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n262), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n260), .A2(KEYINPUT88), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT65), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n277), .B1(new_n240), .B2(G146), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n240), .A2(G146), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n248), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(G128), .B1(new_n279), .B2(new_n254), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT88), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n282), .A2(new_n283), .A3(new_n253), .A4(new_n255), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n276), .A2(new_n250), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n252), .A2(KEYINPUT7), .ZN(new_n286));
  AND3_X1   g100(.A1(new_n285), .A2(KEYINPUT89), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT89), .B1(new_n285), .B2(new_n286), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI211_X1 g103(.A(KEYINPUT90), .B(new_n189), .C1(new_n275), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n220), .A2(new_n232), .ZN(new_n291));
  INV_X1    g105(.A(new_n233), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(KEYINPUT6), .A3(new_n234), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n250), .A2(new_n260), .ZN(new_n295));
  XOR2_X1   g109(.A(new_n252), .B(KEYINPUT86), .Z(new_n296));
  XNOR2_X1  g110(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT6), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n291), .A2(new_n298), .A3(new_n292), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n294), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n290), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n262), .B(new_n274), .C1(new_n288), .C2(new_n287), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT90), .B1(new_n302), .B2(new_n189), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n188), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n189), .B1(new_n275), .B2(new_n289), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT90), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n307), .A2(new_n187), .A3(new_n300), .A4(new_n290), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G469), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n239), .A2(new_n241), .A3(new_n236), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT66), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n235), .A2(KEYINPUT66), .A3(new_n236), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n236), .A2(new_n244), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n313), .A2(new_n314), .B1(new_n280), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n219), .A3(new_n215), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n282), .A2(new_n255), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(KEYINPUT10), .A3(new_n264), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT10), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n259), .A2(new_n235), .ZN(new_n321));
  AND4_X1   g135(.A1(new_n254), .A2(new_n239), .A3(new_n241), .A4(G128), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n218), .A2(new_n229), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n320), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT11), .ZN(new_n326));
  INV_X1    g140(.A(G134), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(G137), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(G137), .ZN(new_n329));
  INV_X1    g143(.A(G137), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(KEYINPUT11), .A3(G134), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G131), .ZN(new_n333));
  INV_X1    g147(.A(G131), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n328), .A2(new_n331), .A3(new_n334), .A4(new_n329), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n317), .A2(new_n319), .A3(new_n325), .A4(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(G110), .B(G140), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n251), .A2(G227), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n339), .B(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n282), .A2(new_n324), .A3(new_n255), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT83), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n322), .B1(new_n281), .B2(new_n280), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT83), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n347), .A3(new_n324), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n264), .B1(new_n322), .B2(new_n321), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n345), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n336), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT12), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n350), .A2(KEYINPUT12), .A3(new_n336), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n343), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n317), .A2(new_n319), .A3(new_n325), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n336), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n342), .B1(new_n357), .B2(new_n338), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n310), .B(new_n189), .C1(new_n355), .C2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n357), .A2(new_n342), .A3(new_n338), .ZN(new_n360));
  INV_X1    g174(.A(new_n338), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(new_n353), .B2(new_n354), .ZN(new_n362));
  OAI211_X1 g176(.A(G469), .B(new_n360), .C1(new_n362), .C2(new_n342), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n310), .A2(new_n189), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n359), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G221), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT9), .B(G234), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n367), .B1(new_n369), .B2(new_n189), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(G214), .B1(G237), .B2(G902), .ZN(new_n373));
  XOR2_X1   g187(.A(new_n373), .B(KEYINPUT84), .Z(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  XOR2_X1   g189(.A(KEYINPUT92), .B(G475), .Z(new_n376));
  NOR2_X1   g190(.A1(G237), .A2(G953), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n377), .A2(G143), .A3(G214), .ZN(new_n378));
  AOI21_X1  g192(.A(G143), .B1(new_n377), .B2(G214), .ZN(new_n379));
  OAI21_X1  g193(.A(G131), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n377), .A2(G214), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n240), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n377), .A2(G143), .A3(G214), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n334), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT17), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n380), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT16), .ZN(new_n387));
  INV_X1    g201(.A(G140), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(G125), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(G125), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n253), .A2(G140), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n389), .B1(new_n392), .B2(new_n387), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n238), .ZN(new_n394));
  XNOR2_X1  g208(.A(G125), .B(G140), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT16), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(G146), .A3(new_n389), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n382), .A2(new_n383), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(KEYINPUT17), .A3(G131), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n386), .A2(new_n394), .A3(new_n397), .A4(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n378), .A2(new_n379), .ZN(new_n401));
  NAND2_X1  g215(.A1(KEYINPUT18), .A2(G131), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n392), .A2(G146), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n395), .A2(new_n238), .ZN(new_n404));
  AOI22_X1  g218(.A1(new_n401), .A2(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT91), .ZN(new_n406));
  INV_X1    g220(.A(new_n402), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n406), .B1(new_n398), .B2(new_n407), .ZN(new_n408));
  AOI211_X1 g222(.A(KEYINPUT91), .B(new_n402), .C1(new_n382), .C2(new_n383), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n405), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G113), .B(G122), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(new_n207), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n400), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n412), .B1(new_n400), .B2(new_n410), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n376), .B1(new_n415), .B2(new_n189), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n251), .A2(G952), .ZN(new_n418));
  NAND2_X1  g232(.A1(G234), .A2(G237), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(G902), .A3(G953), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT21), .B(G898), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n421), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(G475), .A2(G902), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n395), .A2(KEYINPUT19), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n395), .A2(KEYINPUT19), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n238), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n380), .A2(new_n384), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(new_n431), .A3(new_n397), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n412), .B1(new_n410), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n427), .B1(new_n413), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT20), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n410), .A2(new_n432), .ZN(new_n436));
  INV_X1    g250(.A(new_n412), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n400), .A2(new_n410), .A3(new_n412), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(new_n427), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n435), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n417), .A2(new_n426), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n369), .A2(G217), .A3(new_n251), .ZN(new_n445));
  XNOR2_X1  g259(.A(G128), .B(G143), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(new_n327), .ZN(new_n447));
  XNOR2_X1  g261(.A(KEYINPUT93), .B(G122), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G116), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n190), .A2(G122), .A3(new_n191), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n210), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  AND2_X1   g266(.A1(KEYINPUT69), .A2(G116), .ZN(new_n453));
  NOR2_X1   g267(.A1(KEYINPUT69), .A2(G116), .ZN(new_n454));
  INV_X1    g268(.A(G122), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT14), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n456), .A2(KEYINPUT95), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT95), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n459), .B1(new_n450), .B2(KEYINPUT14), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n449), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT96), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT96), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n463), .B(new_n449), .C1(new_n458), .C2(new_n460), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n456), .A2(new_n457), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n452), .B1(new_n466), .B2(G107), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n449), .A2(new_n450), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G107), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n469), .A2(new_n451), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n446), .A2(KEYINPUT13), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n258), .A2(KEYINPUT13), .A3(G143), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(new_n327), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n446), .A2(new_n327), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n471), .A2(new_n473), .B1(new_n474), .B2(KEYINPUT94), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n475), .B1(KEYINPUT94), .B2(new_n474), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n445), .B1(new_n467), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n477), .ZN(new_n479));
  INV_X1    g293(.A(new_n445), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n461), .A2(KEYINPUT96), .B1(new_n457), .B2(new_n456), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n210), .B1(new_n481), .B2(new_n464), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n479), .B(new_n480), .C1(new_n482), .C2(new_n452), .ZN(new_n483));
  AOI21_X1  g297(.A(G902), .B1(new_n478), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G478), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n485), .A2(KEYINPUT15), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  AOI211_X1 g302(.A(G902), .B(new_n486), .C1(new_n478), .C2(new_n483), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n444), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  AND4_X1   g304(.A1(new_n309), .A2(new_n372), .A3(new_n375), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n258), .A2(G119), .ZN(new_n493));
  NOR2_X1   g307(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(G119), .B(G128), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n495), .B1(new_n496), .B2(new_n492), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT80), .B(G110), .ZN(new_n498));
  XOR2_X1   g312(.A(KEYINPUT24), .B(G110), .Z(new_n499));
  OAI22_X1  g313(.A1(new_n497), .A2(new_n498), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(new_n397), .A3(new_n404), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n394), .A2(new_n397), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n497), .A2(G110), .B1(new_n496), .B2(new_n499), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT79), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT79), .B1(new_n502), .B2(new_n503), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT81), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT81), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n508), .B(new_n501), .C1(new_n504), .C2(new_n505), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT22), .B(G137), .ZN(new_n510));
  INV_X1    g324(.A(G234), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n367), .A2(new_n511), .A3(G953), .ZN(new_n512));
  XOR2_X1   g326(.A(new_n510), .B(new_n512), .Z(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n507), .A2(new_n509), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n506), .A2(KEYINPUT81), .A3(new_n513), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(G217), .B1(new_n511), .B2(G902), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT77), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(G902), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT25), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n509), .A2(new_n514), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n497), .A2(G110), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n499), .A2(new_n496), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n253), .A2(KEYINPUT16), .A3(G140), .ZN(new_n527));
  AOI211_X1 g341(.A(new_n238), .B(new_n527), .C1(KEYINPUT16), .C2(new_n395), .ZN(new_n528));
  AOI21_X1  g342(.A(G146), .B1(new_n396), .B2(new_n389), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n525), .B(new_n526), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT79), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT79), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n508), .B1(new_n534), .B2(new_n501), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n524), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n516), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n523), .B(new_n189), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n520), .ZN(new_n539));
  AOI21_X1  g353(.A(G902), .B1(new_n515), .B2(new_n516), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n540), .A2(new_n523), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n522), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT82), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT82), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n544), .B(new_n522), .C1(new_n539), .C2(new_n541), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(G472), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n316), .A2(new_n336), .ZN(new_n548));
  INV_X1    g362(.A(new_n329), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n327), .A2(G137), .ZN(new_n550));
  OAI21_X1  g364(.A(G131), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n335), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n318), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n206), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n204), .A2(new_n203), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n200), .B1(new_n192), .B2(new_n194), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n548), .B(new_n554), .C1(new_n555), .C2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n560), .A2(KEYINPUT28), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n548), .A2(new_n554), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n558), .A2(new_n555), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n559), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n561), .B1(new_n565), .B2(KEYINPUT28), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n377), .A2(G210), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT27), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT26), .B(G101), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n568), .B(new_n569), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n570), .A2(KEYINPUT29), .ZN(new_n571));
  AOI21_X1  g385(.A(G902), .B1(new_n566), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n561), .ZN(new_n574));
  XOR2_X1   g388(.A(new_n570), .B(KEYINPUT72), .Z(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT74), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n280), .A2(new_n315), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n313), .A2(new_n314), .ZN(new_n579));
  AND4_X1   g393(.A1(KEYINPUT67), .A2(new_n336), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT67), .B1(new_n316), .B2(new_n336), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT68), .B1(new_n346), .B2(new_n552), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT68), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n318), .A2(new_n584), .A3(new_n553), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n577), .B(new_n563), .C1(new_n582), .C2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(KEYINPUT73), .B(KEYINPUT28), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n559), .A2(KEYINPUT74), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n583), .B(new_n585), .C1(new_n580), .C2(new_n581), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n590), .B1(new_n563), .B2(new_n591), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n574), .B(new_n576), .C1(new_n589), .C2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT75), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n591), .A2(new_n563), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n587), .B(new_n588), .C1(new_n595), .C2(new_n590), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT75), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n596), .A2(new_n597), .A3(new_n574), .A4(new_n576), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n591), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n548), .A2(new_n554), .A3(KEYINPUT30), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n563), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n559), .ZN(new_n603));
  INV_X1    g417(.A(new_n570), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT29), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n594), .A2(new_n598), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT76), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n573), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n594), .A2(new_n598), .A3(new_n605), .A4(KEYINPUT76), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n547), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n574), .B1(new_n589), .B2(new_n592), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n575), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n602), .A2(new_n559), .A3(new_n570), .ZN(new_n613));
  NOR2_X1   g427(.A1(KEYINPUT71), .A2(KEYINPUT31), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT71), .B(KEYINPUT31), .Z(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n602), .A2(new_n559), .A3(new_n570), .A4(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n612), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT32), .ZN(new_n621));
  NOR2_X1   g435(.A1(G472), .A2(G902), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n621), .B1(new_n620), .B2(new_n622), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n491), .B(new_n546), .C1(new_n610), .C2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G101), .ZN(G3));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n309), .A2(new_n373), .A3(new_n426), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n417), .A2(new_n443), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT98), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT95), .B1(new_n456), .B2(new_n457), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n450), .A2(new_n459), .A3(KEYINPUT14), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n632), .A2(new_n633), .B1(G116), .B2(new_n448), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n465), .B1(new_n634), .B2(new_n463), .ZN(new_n635));
  INV_X1    g449(.A(new_n464), .ZN(new_n636));
  OAI21_X1  g450(.A(G107), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n452), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n480), .B1(new_n639), .B2(new_n479), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n467), .A2(new_n477), .A3(new_n445), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n189), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n631), .B1(new_n642), .B2(new_n485), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n484), .A2(KEYINPUT98), .A3(G478), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n485), .A2(G902), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(KEYINPUT97), .B1(new_n640), .B2(new_n641), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT33), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT97), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n478), .B2(new_n483), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT33), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n647), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n630), .B1(new_n645), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n628), .B1(new_n629), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n630), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n652), .A2(KEYINPUT33), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n652), .A2(KEYINPUT33), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n646), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n642), .A2(new_n631), .A3(new_n485), .ZN(new_n661));
  OAI21_X1  g475(.A(KEYINPUT98), .B1(new_n484), .B2(G478), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n657), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n373), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n304), .B2(new_n308), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n664), .A2(new_n666), .A3(KEYINPUT99), .A4(new_n426), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n656), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n543), .A2(new_n545), .A3(new_n372), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n620), .A2(new_n189), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(G472), .ZN(new_n671));
  INV_X1    g485(.A(new_n601), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n591), .B2(new_n599), .ZN(new_n673));
  AOI211_X1 g487(.A(new_n560), .B(new_n604), .C1(new_n673), .C2(new_n563), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n619), .B1(new_n674), .B2(new_n614), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n576), .B1(new_n596), .B2(new_n574), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n622), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n669), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n668), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT34), .B(G104), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G6));
  INV_X1    g496(.A(new_n427), .ZN(new_n683));
  AOI211_X1 g497(.A(KEYINPUT20), .B(new_n683), .C1(new_n438), .C2(new_n439), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(KEYINPUT100), .B2(new_n435), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT100), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n434), .A2(new_n686), .A3(KEYINPUT20), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n417), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n642), .A2(new_n486), .ZN(new_n689));
  INV_X1    g503(.A(new_n489), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n309), .A2(new_n691), .A3(new_n373), .A4(new_n426), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT101), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT101), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n666), .A2(new_n694), .A3(new_n426), .A4(new_n691), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n679), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT35), .B(G107), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G9));
  AOI21_X1  g513(.A(new_n547), .B1(new_n620), .B2(new_n189), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n620), .B2(new_n622), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n514), .A2(KEYINPUT36), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n506), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n521), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n704), .B1(new_n539), .B2(new_n541), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n491), .A2(new_n701), .A3(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT37), .B(G110), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT102), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n706), .B(new_n708), .ZN(G12));
  AND4_X1   g523(.A1(new_n309), .A2(new_n372), .A3(new_n373), .A4(new_n705), .ZN(new_n710));
  XOR2_X1   g524(.A(new_n420), .B(KEYINPUT104), .Z(new_n711));
  OR2_X1    g525(.A1(KEYINPUT103), .A2(G900), .ZN(new_n712));
  NAND2_X1  g526(.A1(KEYINPUT103), .A2(G900), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n423), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n691), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n710), .B(new_n717), .C1(new_n610), .C2(new_n625), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G128), .ZN(G30));
  OAI211_X1 g533(.A(new_n373), .B(new_n630), .C1(new_n488), .C2(new_n489), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n540), .A2(new_n523), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n519), .B1(new_n540), .B2(new_n523), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n722), .A2(new_n723), .B1(new_n521), .B2(new_n703), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n677), .A2(KEYINPUT32), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n565), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n576), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n189), .B1(new_n674), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(G472), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n725), .B1(new_n728), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n715), .B(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n372), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT40), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n309), .B(KEYINPUT38), .ZN(new_n739));
  OR2_X1    g553(.A1(new_n737), .A2(KEYINPUT40), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n733), .A2(new_n738), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G143), .ZN(G45));
  OAI211_X1 g556(.A(new_n630), .B(new_n715), .C1(new_n645), .C2(new_n654), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n744), .B(new_n710), .C1(new_n610), .C2(new_n625), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G146), .ZN(G48));
  NAND2_X1  g560(.A1(new_n543), .A2(new_n545), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n606), .A2(new_n607), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n609), .A3(new_n572), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(G472), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n747), .B1(new_n750), .B2(new_n728), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n355), .A2(new_n358), .ZN(new_n752));
  OAI21_X1  g566(.A(G469), .B1(new_n752), .B2(G902), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n371), .A3(new_n359), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n668), .A2(new_n751), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(KEYINPUT41), .B(G113), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(G15));
  NAND3_X1  g572(.A1(new_n696), .A2(new_n751), .A3(new_n755), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G116), .ZN(G18));
  AOI22_X1  g574(.A1(new_n749), .A2(G472), .B1(new_n726), .B2(new_n727), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n666), .A2(new_n490), .A3(new_n705), .A4(new_n755), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n193), .ZN(G21));
  AOI21_X1  g578(.A(new_n720), .B1(new_n304), .B2(new_n308), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n616), .B(new_n619), .C1(new_n576), .C2(new_n566), .ZN(new_n766));
  AOI22_X1  g580(.A1(new_n670), .A2(G472), .B1(new_n622), .B2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n542), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n754), .A2(new_n425), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n765), .A2(new_n767), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G122), .ZN(G24));
  NAND2_X1  g585(.A1(new_n766), .A2(new_n622), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n671), .A2(new_n705), .A3(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n309), .A2(new_n373), .A3(new_n755), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n773), .A2(new_n743), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n253), .ZN(G27));
  INV_X1    g590(.A(KEYINPUT107), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n366), .A2(KEYINPUT106), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT106), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n359), .A2(new_n363), .A3(new_n779), .A4(new_n365), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n778), .A2(new_n371), .A3(new_n780), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n304), .A2(new_n308), .A3(new_n373), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n777), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n778), .A2(new_n371), .A3(new_n780), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n304), .A2(new_n308), .A3(new_n373), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n784), .A2(new_n785), .A3(KEYINPUT107), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n744), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n768), .B1(new_n610), .B2(new_n625), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT42), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n781), .A2(new_n782), .A3(new_n777), .ZN(new_n790));
  OAI21_X1  g604(.A(KEYINPUT107), .B1(new_n784), .B2(new_n785), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n743), .A2(KEYINPUT42), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n751), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n789), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(new_n334), .ZN(G33));
  NAND3_X1  g610(.A1(new_n751), .A2(new_n717), .A3(new_n792), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT108), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n751), .A2(new_n792), .A3(KEYINPUT108), .A4(new_n717), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G134), .ZN(G36));
  OAI21_X1  g616(.A(new_n360), .B1(new_n362), .B2(new_n342), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT45), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(G469), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n803), .A2(new_n804), .ZN(new_n807));
  OR3_X1    g621(.A1(new_n806), .A2(KEYINPUT109), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(KEYINPUT109), .B1(new_n806), .B2(new_n807), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n364), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n810), .A2(KEYINPUT46), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n359), .B1(new_n810), .B2(KEYINPUT46), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n371), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n813), .A2(new_n735), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n678), .A2(new_n705), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT110), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n645), .A2(new_n654), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n630), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT43), .ZN(new_n821));
  OR3_X1    g635(.A1(new_n818), .A2(KEYINPUT43), .A3(new_n630), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n817), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT44), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n785), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n815), .B(new_n825), .C1(new_n824), .C2(new_n823), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G137), .ZN(G39));
  INV_X1    g641(.A(KEYINPUT47), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n813), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(KEYINPUT47), .B(new_n371), .C1(new_n811), .C2(new_n812), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n546), .A2(new_n743), .A3(new_n785), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(new_n761), .A3(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(G140), .ZN(G42));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n835));
  INV_X1    g649(.A(new_n711), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n821), .A2(new_n836), .A3(new_n822), .ZN(new_n837));
  INV_X1    g651(.A(new_n772), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n838), .A2(new_n700), .A3(new_n542), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n739), .A2(new_n373), .A3(new_n754), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n837), .A2(KEYINPUT50), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT50), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n821), .A2(new_n839), .A3(new_n836), .A4(new_n822), .ZN(new_n843));
  INV_X1    g657(.A(new_n840), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n838), .A2(new_n700), .A3(new_n724), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n785), .A2(new_n754), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n837), .A2(new_n847), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n821), .A2(new_n836), .A3(new_n822), .A4(new_n849), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT117), .B1(new_n851), .B2(new_n773), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n726), .A2(new_n727), .B1(G472), .B2(new_n731), .ZN(new_n854));
  AND4_X1   g668(.A1(new_n546), .A2(new_n854), .A3(new_n421), .A4(new_n849), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(new_n657), .A3(new_n818), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n846), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n753), .A2(new_n359), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n370), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n829), .A2(new_n830), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n843), .A2(new_n785), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(KEYINPUT116), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n860), .A2(new_n861), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT116), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n857), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT51), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n835), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n855), .A2(new_n664), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n418), .B(new_n869), .C1(new_n843), .C2(new_n774), .ZN(new_n870));
  OR3_X1    g684(.A1(new_n851), .A2(KEYINPUT48), .A3(new_n788), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT48), .B1(new_n851), .B2(new_n788), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n857), .A2(KEYINPUT51), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n861), .B1(new_n860), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(new_n875), .B2(new_n860), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n873), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n868), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n866), .A2(new_n835), .A3(new_n867), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT52), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n370), .B1(new_n366), .B2(KEYINPUT106), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n309), .A2(new_n715), .A3(new_n883), .A4(new_n780), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT114), .B1(new_n733), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT114), .ZN(new_n887));
  NOR4_X1   g701(.A1(new_n854), .A2(new_n884), .A3(new_n725), .A4(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n848), .A2(new_n744), .A3(new_n666), .A4(new_n755), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n745), .A2(new_n890), .A3(new_n718), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n882), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n732), .B1(new_n623), .B2(new_n624), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n705), .A2(new_n720), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n887), .B1(new_n895), .B2(new_n884), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n733), .A2(KEYINPUT114), .A3(new_n885), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n666), .A2(new_n372), .A3(new_n705), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n750), .B2(new_n728), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n775), .B1(new_n900), .B2(new_n717), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n898), .A2(new_n901), .A3(KEYINPUT52), .A4(new_n745), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n892), .A2(KEYINPUT115), .A3(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n891), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT115), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n904), .A2(new_n905), .A3(KEYINPUT52), .A4(new_n898), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT53), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n770), .B1(new_n761), .B2(new_n762), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n756), .A2(new_n759), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT112), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n546), .B(new_n755), .C1(new_n610), .C2(new_n625), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n909), .B1(new_n915), .B2(new_n668), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n916), .A2(KEYINPUT112), .A3(new_n759), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT113), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n309), .A2(new_n375), .A3(new_n426), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n919), .B1(new_n920), .B2(new_n655), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n374), .B1(new_n304), .B2(new_n308), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n664), .A2(new_n922), .A3(KEYINPUT113), .A4(new_n426), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n679), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n543), .A2(new_n545), .A3(new_n372), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n630), .B1(new_n690), .B2(new_n689), .ZN(new_n926));
  AND4_X1   g740(.A1(new_n309), .A2(new_n375), .A3(new_n426), .A4(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n925), .A2(new_n701), .A3(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n924), .A2(new_n626), .A3(new_n706), .A4(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n792), .A2(new_n744), .A3(new_n848), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n750), .A2(new_n728), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n372), .A2(new_n705), .ZN(new_n932));
  INV_X1    g746(.A(new_n715), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n688), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n488), .A2(new_n489), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NOR4_X1   g750(.A1(new_n932), .A2(new_n785), .A3(new_n934), .A4(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n931), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n930), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n929), .A2(new_n939), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n751), .A2(new_n792), .A3(new_n793), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT42), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n743), .B1(new_n790), .B2(new_n791), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n542), .B1(new_n750), .B2(new_n728), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n940), .A2(new_n801), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n918), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n907), .A2(new_n908), .A3(new_n948), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n940), .A2(new_n801), .A3(new_n946), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT112), .B1(new_n916), .B2(new_n759), .ZN(new_n951));
  AND4_X1   g765(.A1(KEYINPUT112), .A2(new_n756), .A3(new_n759), .A4(new_n910), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n892), .A2(new_n902), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n950), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(KEYINPUT53), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n949), .A2(new_n956), .A3(KEYINPUT54), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n626), .A2(new_n706), .A3(new_n928), .ZN(new_n958));
  AOI22_X1  g772(.A1(new_n943), .A2(new_n848), .B1(new_n931), .B2(new_n937), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n958), .A2(new_n959), .A3(new_n924), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n960), .A2(new_n795), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n961), .A2(new_n801), .A3(new_n913), .A4(new_n917), .ZN(new_n962));
  INV_X1    g776(.A(new_n954), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n908), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n916), .A2(KEYINPUT53), .A3(new_n759), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n947), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n966), .A2(new_n906), .A3(new_n903), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n957), .B1(KEYINPUT54), .B2(new_n968), .ZN(new_n969));
  OAI22_X1  g783(.A1(new_n881), .A2(new_n969), .B1(G952), .B2(G953), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n858), .B(KEYINPUT49), .Z(new_n971));
  NOR3_X1   g785(.A1(new_n820), .A2(new_n971), .A3(new_n893), .ZN(new_n972));
  INV_X1    g786(.A(new_n739), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n768), .A2(new_n375), .A3(new_n371), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT111), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n972), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n970), .A2(new_n976), .ZN(G75));
  NOR2_X1   g791(.A1(new_n251), .A2(G952), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n189), .B1(new_n964), .B2(new_n967), .ZN(new_n980));
  AOI21_X1  g794(.A(KEYINPUT56), .B1(new_n980), .B2(G210), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n294), .A2(new_n299), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(new_n297), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT55), .Z(new_n984));
  OAI21_X1  g798(.A(new_n979), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  AOI22_X1  g799(.A1(new_n908), .A2(new_n955), .B1(new_n907), .B2(new_n966), .ZN(new_n986));
  OAI21_X1  g800(.A(KEYINPUT120), .B1(new_n986), .B2(new_n189), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT120), .ZN(new_n988));
  AOI21_X1  g802(.A(KEYINPUT53), .B1(new_n948), .B2(new_n954), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n903), .A2(new_n906), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n911), .A2(new_n908), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n991), .A2(new_n946), .A3(new_n801), .A4(new_n940), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n988), .B(G902), .C1(new_n989), .C2(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n987), .A2(new_n188), .A3(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT56), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n984), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n985), .B1(new_n995), .B2(new_n997), .ZN(G51));
  AND2_X1   g812(.A1(new_n808), .A2(new_n809), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n987), .A2(new_n999), .A3(new_n994), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT121), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n364), .B(KEYINPUT57), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n989), .A2(KEYINPUT54), .A3(new_n993), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT54), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1004), .B1(new_n964), .B2(new_n967), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1002), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n752), .ZN(new_n1007));
  AOI22_X1  g821(.A1(new_n1000), .A2(new_n1001), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n987), .A2(KEYINPUT121), .A3(new_n999), .A4(new_n994), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n978), .B1(new_n1008), .B2(new_n1009), .ZN(G54));
  NAND2_X1  g824(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT122), .Z(new_n1012));
  NAND3_X1  g826(.A1(new_n987), .A2(new_n994), .A3(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1013), .A2(new_n438), .A3(new_n439), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n987), .A2(new_n440), .A3(new_n994), .A4(new_n1012), .ZN(new_n1015));
  AND3_X1   g829(.A1(new_n1014), .A2(new_n979), .A3(new_n1015), .ZN(G60));
  NAND2_X1  g830(.A1(new_n650), .A2(new_n653), .ZN(new_n1017));
  NAND2_X1  g831(.A1(G478), .A2(G902), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1018), .B(KEYINPUT59), .ZN(new_n1019));
  OAI211_X1 g833(.A(new_n1017), .B(new_n1019), .C1(new_n1003), .C2(new_n1005), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(new_n979), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1017), .B1(new_n969), .B2(new_n1019), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1021), .A2(new_n1022), .ZN(G63));
  NAND2_X1  g837(.A1(G217), .A2(G902), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1024), .B(KEYINPUT60), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1025), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n968), .A2(new_n703), .A3(new_n1026), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n986), .A2(new_n1025), .ZN(new_n1028));
  OAI211_X1 g842(.A(new_n1027), .B(new_n979), .C1(new_n1028), .C2(new_n517), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT61), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1029), .B(new_n1030), .ZN(G66));
  INV_X1    g845(.A(new_n424), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n251), .B1(new_n1032), .B2(G224), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n953), .A2(new_n924), .A3(new_n958), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1033), .B1(new_n1034), .B2(new_n251), .ZN(new_n1035));
  INV_X1    g849(.A(G898), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n982), .B1(new_n1036), .B2(G953), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n1035), .B(new_n1037), .ZN(G69));
  NOR2_X1   g852(.A1(new_n428), .A2(new_n429), .ZN(new_n1039));
  XNOR2_X1  g853(.A(new_n673), .B(new_n1039), .ZN(new_n1040));
  XOR2_X1   g854(.A(KEYINPUT123), .B(KEYINPUT124), .Z(new_n1041));
  XNOR2_X1  g855(.A(new_n1040), .B(new_n1041), .ZN(new_n1042));
  NAND2_X1  g856(.A1(G900), .A2(G953), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n944), .A2(new_n765), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n904), .B1(new_n814), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n1045), .A2(new_n795), .ZN(new_n1046));
  NAND4_X1  g860(.A1(new_n1046), .A2(new_n801), .A3(new_n826), .A4(new_n833), .ZN(new_n1047));
  OAI211_X1 g861(.A(new_n1042), .B(new_n1043), .C1(new_n1047), .C2(G953), .ZN(new_n1048));
  INV_X1    g862(.A(KEYINPUT126), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g864(.A(new_n1042), .B(KEYINPUT125), .ZN(new_n1051));
  INV_X1    g865(.A(new_n1051), .ZN(new_n1052));
  NOR2_X1   g866(.A1(new_n737), .A2(new_n785), .ZN(new_n1053));
  OAI211_X1 g867(.A(new_n751), .B(new_n1053), .C1(new_n664), .C2(new_n926), .ZN(new_n1054));
  NAND3_X1  g868(.A1(new_n826), .A2(new_n833), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n904), .A2(new_n741), .ZN(new_n1056));
  XNOR2_X1  g870(.A(new_n1056), .B(KEYINPUT62), .ZN(new_n1057));
  OR2_X1    g871(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n1052), .B1(new_n1058), .B2(new_n251), .ZN(new_n1059));
  AOI21_X1  g873(.A(new_n251), .B1(G227), .B2(G900), .ZN(new_n1060));
  OR3_X1    g874(.A1(new_n1050), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  OAI21_X1  g875(.A(new_n1060), .B1(new_n1050), .B2(new_n1059), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1061), .A2(new_n1062), .ZN(G72));
  NAND2_X1  g877(.A1(new_n603), .A2(new_n570), .ZN(new_n1064));
  NAND2_X1  g878(.A1(G472), .A2(G902), .ZN(new_n1065));
  XOR2_X1   g879(.A(new_n1065), .B(KEYINPUT63), .Z(new_n1066));
  OAI211_X1 g880(.A(KEYINPUT127), .B(new_n1066), .C1(new_n1058), .C2(new_n1034), .ZN(new_n1067));
  INV_X1    g881(.A(KEYINPUT127), .ZN(new_n1068));
  NOR3_X1   g882(.A1(new_n1055), .A2(new_n1034), .A3(new_n1057), .ZN(new_n1069));
  INV_X1    g883(.A(new_n1066), .ZN(new_n1070));
  OAI21_X1  g884(.A(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g885(.A(new_n1064), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g886(.A(new_n1066), .B1(new_n1047), .B2(new_n1034), .ZN(new_n1073));
  NAND4_X1  g887(.A1(new_n1073), .A2(new_n559), .A3(new_n604), .A4(new_n602), .ZN(new_n1074));
  NAND2_X1  g888(.A1(new_n603), .A2(new_n604), .ZN(new_n1075));
  AOI21_X1  g889(.A(new_n1070), .B1(new_n1075), .B2(new_n613), .ZN(new_n1076));
  NAND3_X1  g890(.A1(new_n949), .A2(new_n956), .A3(new_n1076), .ZN(new_n1077));
  NAND3_X1  g891(.A1(new_n1074), .A2(new_n979), .A3(new_n1077), .ZN(new_n1078));
  NOR2_X1   g892(.A1(new_n1072), .A2(new_n1078), .ZN(G57));
endmodule


