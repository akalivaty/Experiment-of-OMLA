//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n581,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n624, new_n627, new_n628, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1214,
    new_n1215;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT66), .ZN(G261));
  NAND2_X1  g031(.A1(new_n454), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n452), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n460), .B1(new_n459), .B2(new_n458), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT68), .Z(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT69), .B1(new_n463), .B2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n463), .A2(G2104), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n464), .A2(new_n467), .A3(G137), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G101), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(new_n468), .A3(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n471), .A2(new_n476), .ZN(G160));
  NAND3_X1  g052(.A1(new_n464), .A2(new_n467), .A3(new_n468), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT70), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n478), .B(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n472), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n480), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND4_X1  g064(.A1(new_n473), .A2(new_n468), .A3(G138), .A4(new_n472), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(G126), .A2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(KEYINPUT4), .A2(G138), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n495), .A2(new_n468), .A3(new_n464), .A4(new_n467), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(G2104), .C1(G114), .C2(new_n472), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n492), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT73), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT72), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n504), .A2(new_n506), .B1(new_n503), .B2(G543), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n501), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n503), .A2(G543), .ZN(new_n511));
  AND3_X1   g086(.A1(new_n505), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n512));
  AOI21_X1  g087(.A(KEYINPUT72), .B1(new_n505), .B2(KEYINPUT5), .ZN(new_n513));
  OAI211_X1 g088(.A(G62), .B(new_n511), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n509), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n509), .A2(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT71), .B1(new_n519), .B2(G651), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(new_n509), .A3(KEYINPUT6), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n518), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n507), .A2(new_n523), .A3(G88), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(G50), .A3(G543), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n510), .A2(new_n517), .A3(new_n524), .A4(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND2_X1  g102(.A1(new_n507), .A2(new_n523), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G89), .ZN(new_n530));
  AOI211_X1 g105(.A(new_n505), .B(new_n518), .C1(new_n520), .C2(new_n522), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G51), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n507), .A2(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND3_X1   g112(.A1(new_n530), .A2(new_n532), .A3(new_n537), .ZN(G168));
  AOI22_X1  g113(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n509), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n523), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n528), .A2(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(KEYINPUT74), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n545), .A2(KEYINPUT74), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(G171));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n528), .A2(new_n550), .B1(new_n542), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT76), .ZN(new_n553));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n509), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n559), .B1(new_n558), .B2(new_n557), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n553), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  INV_X1    g142(.A(G53), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT9), .B1(new_n542), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n531), .A2(new_n570), .A3(G53), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n569), .A2(new_n571), .B1(G91), .B2(new_n529), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n555), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g152(.A(KEYINPUT77), .B(new_n573), .C1(new_n555), .C2(new_n574), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n577), .A2(G651), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n572), .A2(new_n579), .ZN(G299));
  INV_X1    g155(.A(new_n548), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n546), .ZN(G301));
  NAND3_X1  g157(.A1(new_n530), .A2(new_n532), .A3(new_n537), .ZN(G286));
  INV_X1    g158(.A(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(KEYINPUT78), .B1(new_n528), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n507), .A2(new_n523), .A3(new_n586), .A4(G87), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n523), .A2(G49), .A3(G543), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n588), .A2(new_n592), .ZN(G288));
  NAND3_X1  g168(.A1(new_n507), .A2(new_n523), .A3(G86), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n507), .A2(new_n523), .A3(KEYINPUT79), .A4(G86), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g173(.A(G61), .B(new_n511), .C1(new_n512), .C2(new_n513), .ZN(new_n599));
  NAND2_X1  g174(.A1(G73), .A2(G543), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(new_n531), .B2(G48), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n598), .A2(new_n602), .ZN(G305));
  AOI22_X1  g178(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(new_n509), .ZN(new_n605));
  INV_X1    g180(.A(G85), .ZN(new_n606));
  INV_X1    g181(.A(G47), .ZN(new_n607));
  OAI22_X1  g182(.A1(new_n528), .A2(new_n606), .B1(new_n542), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(new_n529), .A2(G92), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  XOR2_X1   g189(.A(KEYINPUT80), .B(G66), .Z(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n555), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n616), .A2(G651), .B1(G54), .B2(new_n531), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g195(.A(new_n619), .B1(G171), .B2(G868), .ZN(G321));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NOR2_X1   g197(.A1(G286), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(G299), .B(KEYINPUT81), .Z(new_n624));
  AOI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(new_n622), .ZN(G297));
  XNOR2_X1  g200(.A(G297), .B(KEYINPUT82), .ZN(G280));
  INV_X1    g201(.A(new_n618), .ZN(new_n627));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n561), .A2(new_n622), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n618), .A2(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(new_n622), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n482), .A2(G135), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n484), .A2(G123), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n637));
  INV_X1    g212(.A(G111), .ZN(new_n638));
  AOI22_X1  g213(.A1(new_n636), .A2(new_n637), .B1(new_n638), .B2(G2105), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n637), .B2(new_n636), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n634), .A2(new_n635), .A3(new_n640), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(G2096), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(G2096), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n472), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT12), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2100), .Z(new_n647));
  NAND3_X1  g222(.A1(new_n642), .A2(new_n643), .A3(new_n647), .ZN(G156));
  XOR2_X1   g223(.A(KEYINPUT15), .B(G2435), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2438), .ZN(new_n650));
  XOR2_X1   g225(.A(G2427), .B(G2430), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT84), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(KEYINPUT14), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2451), .B(G2454), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n655), .B(new_n659), .Z(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(G14), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n663), .B2(new_n661), .ZN(G401));
  XNOR2_X1  g240(.A(G2084), .B(G2090), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT85), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2072), .B(G2078), .Z(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n667), .A2(new_n668), .ZN(new_n674));
  INV_X1    g249(.A(new_n670), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT88), .B(KEYINPUT17), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n674), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n670), .B(KEYINPUT87), .Z(new_n680));
  OAI211_X1 g255(.A(new_n679), .B(new_n669), .C1(new_n674), .C2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n673), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G2096), .B(G2100), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G227));
  XOR2_X1   g259(.A(G1971), .B(G1976), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  XOR2_X1   g262(.A(G1961), .B(G1966), .Z(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT20), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n687), .A2(new_n688), .ZN(new_n692));
  NOR3_X1   g267(.A1(new_n686), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(new_n686), .B2(new_n692), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1981), .B(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(G229));
  INV_X1    g276(.A(G1961), .ZN(new_n702));
  NAND2_X1  g277(.A1(G171), .A2(G16), .ZN(new_n703));
  NOR2_X1   g278(.A1(G5), .A2(G16), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(KEYINPUT99), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT99), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n703), .A2(new_n708), .A3(new_n705), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n702), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT100), .Z(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G33), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT25), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n473), .A2(new_n468), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n717), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n716), .B1(new_n718), .B2(new_n472), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n482), .B2(G139), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT94), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n713), .B1(new_n722), .B2(new_n712), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(G2072), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n712), .A2(G32), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n482), .A2(G141), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n484), .A2(G129), .ZN(new_n727));
  NAND3_X1  g302(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT26), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  AND2_X1   g306(.A1(G105), .A2(G2104), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n730), .A2(new_n731), .B1(new_n472), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n726), .A2(new_n727), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n725), .B1(new_n734), .B2(G29), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT27), .B(G1996), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT24), .ZN(new_n738));
  INV_X1    g313(.A(G34), .ZN(new_n739));
  AOI21_X1  g314(.A(G29), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n738), .B2(new_n739), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G160), .B2(new_n712), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n742), .A2(G2084), .ZN(new_n743));
  NOR3_X1   g318(.A1(new_n724), .A2(new_n737), .A3(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT95), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n723), .B2(G2072), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n723), .A2(new_n745), .A3(G2072), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n744), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(KEYINPUT96), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n712), .A2(G35), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G162), .B2(new_n712), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(KEYINPUT29), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(KEYINPUT29), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G2090), .ZN(new_n756));
  INV_X1    g331(.A(G2090), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n753), .A2(new_n757), .A3(new_n754), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n712), .A2(G26), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT28), .Z(new_n760));
  OAI21_X1  g335(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n761));
  INV_X1    g336(.A(G116), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(G2105), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n484), .B2(G128), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT93), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n482), .B2(G140), .ZN(new_n766));
  INV_X1    g341(.A(G140), .ZN(new_n767));
  NOR3_X1   g342(.A1(new_n481), .A2(KEYINPUT93), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n764), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n760), .B1(new_n769), .B2(G29), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2067), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n756), .A2(new_n758), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G16), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G21), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G168), .B2(new_n773), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n775), .A2(G1966), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT97), .Z(new_n777));
  INV_X1    g352(.A(G1956), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n773), .A2(G20), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT23), .Z(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G299), .B2(G16), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n777), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n562), .A2(G16), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G16), .B2(G19), .ZN(new_n784));
  INV_X1    g359(.A(G1341), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n742), .A2(G2084), .ZN(new_n787));
  OAI221_X1 g362(.A(new_n787), .B1(new_n775), .B2(G1966), .C1(new_n641), .C2(new_n712), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n773), .A2(G4), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n627), .B2(new_n773), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n791), .A2(G1348), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n791), .A2(G1348), .ZN(new_n793));
  NOR2_X1   g368(.A1(G27), .A2(G29), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G164), .B2(G29), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n795), .A2(G2078), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n795), .A2(G2078), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT31), .B(G11), .ZN(new_n798));
  INV_X1    g373(.A(G28), .ZN(new_n799));
  AOI21_X1  g374(.A(G29), .B1(new_n799), .B2(KEYINPUT30), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  OAI22_X1  g376(.A1(new_n801), .A2(KEYINPUT98), .B1(KEYINPUT30), .B2(new_n799), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n801), .A2(KEYINPUT98), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n798), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OR3_X1    g379(.A1(new_n796), .A2(new_n797), .A3(new_n804), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n792), .A2(new_n793), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n782), .A2(new_n789), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n707), .A2(new_n702), .A3(new_n709), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n781), .A2(new_n778), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n784), .B2(new_n785), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n808), .B(new_n810), .C1(new_n735), .C2(new_n736), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n772), .A2(new_n807), .A3(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT96), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n744), .B(new_n813), .C1(new_n746), .C2(new_n748), .ZN(new_n814));
  AND4_X1   g389(.A1(new_n711), .A2(new_n750), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n773), .A2(G22), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G166), .B2(new_n773), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(KEYINPUT92), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(KEYINPUT92), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(G1971), .ZN(new_n821));
  INV_X1    g396(.A(G1971), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n818), .A2(new_n822), .A3(new_n819), .ZN(new_n823));
  NOR2_X1   g398(.A1(G16), .A2(G23), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n591), .B1(new_n585), .B2(new_n587), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n824), .B1(new_n825), .B2(G16), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT33), .B(G1976), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n826), .B(new_n829), .ZN(new_n830));
  MUX2_X1   g405(.A(G6), .B(G305), .S(G16), .Z(new_n831));
  XOR2_X1   g406(.A(KEYINPUT32), .B(G1981), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT89), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n831), .B(new_n833), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n821), .A2(new_n823), .A3(new_n830), .A4(new_n834), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n835), .A2(KEYINPUT34), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(KEYINPUT34), .ZN(new_n837));
  OR2_X1    g412(.A1(G25), .A2(G29), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n482), .A2(G131), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n484), .A2(G119), .ZN(new_n840));
  OR2_X1    g415(.A1(G95), .A2(G2105), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n841), .B(G2104), .C1(G107), .C2(new_n472), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n838), .B1(new_n843), .B2(new_n712), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT35), .B(G1991), .Z(new_n845));
  AND2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n773), .A2(G24), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n609), .B2(new_n773), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G1986), .ZN(new_n850));
  NOR3_X1   g425(.A1(new_n846), .A2(new_n847), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n836), .A2(new_n837), .A3(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT36), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n815), .A2(new_n853), .ZN(G311));
  AND3_X1   g429(.A1(new_n815), .A2(new_n853), .A3(KEYINPUT101), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT101), .B1(new_n815), .B2(new_n853), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(G150));
  NAND2_X1  g432(.A1(new_n627), .A2(G559), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT38), .ZN(new_n859));
  AOI22_X1  g434(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(new_n509), .ZN(new_n861));
  INV_X1    g436(.A(G93), .ZN(new_n862));
  INV_X1    g437(.A(G55), .ZN(new_n863));
  OAI22_X1  g438(.A1(new_n528), .A2(new_n862), .B1(new_n542), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n561), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n553), .A2(new_n560), .A3(new_n865), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n859), .B(new_n869), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n870), .A2(KEYINPUT39), .ZN(new_n871));
  INV_X1    g446(.A(G860), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(KEYINPUT39), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n865), .A2(new_n872), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT37), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(G145));
  XOR2_X1   g452(.A(new_n641), .B(G160), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n488), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n769), .B(new_n499), .ZN(new_n880));
  INV_X1    g455(.A(new_n734), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n880), .A2(new_n881), .ZN(new_n883));
  OR3_X1    g458(.A1(new_n882), .A2(new_n883), .A3(new_n720), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n843), .B(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n645), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n843), .B(KEYINPUT102), .ZN(new_n888));
  INV_X1    g463(.A(new_n645), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n482), .A2(G142), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n484), .A2(G130), .ZN(new_n893));
  OR2_X1    g468(.A1(G106), .A2(G2105), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n894), .B(G2104), .C1(G118), .C2(new_n472), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n896), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n887), .A2(new_n890), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n722), .B1(new_n882), .B2(new_n883), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n884), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n900), .B1(new_n884), .B2(new_n901), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n879), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n904), .ZN(new_n906));
  INV_X1    g481(.A(new_n879), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n907), .A3(new_n902), .ZN(new_n908));
  INV_X1    g483(.A(G37), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g486(.A1(new_n867), .A2(new_n868), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT103), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n912), .A2(KEYINPUT103), .ZN(new_n915));
  INV_X1    g490(.A(new_n631), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n912), .A2(KEYINPUT103), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n631), .B1(new_n918), .B2(new_n913), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n618), .B(G299), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT41), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n921), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n917), .A2(new_n919), .A3(new_n924), .ZN(new_n925));
  OR3_X1    g500(.A1(new_n923), .A2(KEYINPUT42), .A3(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(G303), .B(G305), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n609), .B(new_n825), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT104), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  XOR2_X1   g506(.A(new_n930), .B(new_n931), .Z(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT42), .B1(new_n923), .B2(new_n925), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n926), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n933), .B1(new_n926), .B2(new_n934), .ZN(new_n936));
  OAI21_X1  g511(.A(G868), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n866), .A2(new_n622), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(G295));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n938), .ZN(G331));
  AOI21_X1  g515(.A(G171), .B1(new_n867), .B2(new_n868), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n867), .A2(G171), .A3(new_n868), .ZN(new_n943));
  AOI21_X1  g518(.A(G168), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n943), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n945), .A2(new_n941), .A3(G286), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n922), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT105), .ZN(new_n948));
  INV_X1    g523(.A(new_n944), .ZN(new_n949));
  INV_X1    g524(.A(new_n946), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(new_n950), .A3(new_n924), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n922), .B(new_n952), .C1(new_n944), .C2(new_n946), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n948), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(G37), .B1(new_n954), .B2(new_n933), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n948), .A2(new_n932), .A3(new_n951), .A4(new_n953), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT43), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n921), .A2(new_n958), .A3(KEYINPUT41), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(new_n922), .B2(new_n958), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n944), .A2(new_n946), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n951), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(G37), .B1(new_n962), .B2(new_n933), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n963), .A2(KEYINPUT43), .A3(new_n956), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT44), .B1(new_n957), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(new_n955), .B2(new_n956), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n963), .A2(new_n967), .A3(new_n956), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n965), .A2(new_n970), .ZN(G397));
  INV_X1    g546(.A(G1384), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n499), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n476), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n469), .A2(new_n470), .ZN(new_n977));
  OAI211_X1 g552(.A(G40), .B(new_n976), .C1(new_n977), .C2(G2105), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G2067), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n769), .B(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G1996), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n734), .B(new_n982), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n843), .B(new_n845), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OR2_X1    g561(.A1(G290), .A2(G1986), .ZN(new_n987));
  NAND2_X1  g562(.A1(G290), .A2(G1986), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n979), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G8), .ZN(new_n991));
  INV_X1    g566(.A(G40), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n471), .A2(new_n992), .A3(new_n476), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n972), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n975), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT107), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT107), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n975), .A2(new_n997), .A3(new_n993), .A4(new_n994), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n822), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n499), .A2(new_n1000), .A3(new_n972), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT108), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n499), .A2(KEYINPUT108), .A3(new_n1000), .A4(new_n972), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1000), .B1(new_n499), .B2(new_n972), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(new_n978), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n757), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n991), .B1(new_n999), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT111), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n524), .B(new_n525), .C1(new_n516), .C2(KEYINPUT73), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n508), .A2(new_n501), .A3(new_n509), .ZN(new_n1012));
  OAI211_X1 g587(.A(KEYINPUT55), .B(G8), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT109), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(G303), .A2(KEYINPUT109), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT110), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT110), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1015), .A2(new_n1019), .A3(new_n1016), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  AND4_X1   g597(.A1(new_n1010), .A2(new_n1018), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1021), .B1(new_n1017), .B2(KEYINPUT110), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1010), .B1(new_n1024), .B2(new_n1020), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1009), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1976), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT52), .B1(G288), .B2(new_n1027), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n499), .A2(new_n972), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n991), .B1(new_n1029), .B2(new_n993), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n588), .A2(new_n592), .A3(G1976), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1028), .A2(KEYINPUT112), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n825), .B2(G1976), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1033), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1032), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1035), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1029), .A2(new_n993), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(G8), .ZN(new_n1041));
  INV_X1    g616(.A(G1981), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n598), .A2(new_n602), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n523), .A2(G48), .A3(G543), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT113), .B(G86), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n507), .A2(new_n523), .A3(new_n1045), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n507), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1044), .B(new_n1046), .C1(new_n1047), .C2(new_n509), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G1981), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1043), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT49), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1041), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1043), .A2(KEYINPUT49), .A3(new_n1049), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1039), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1038), .A2(new_n1054), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1018), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1007), .A2(new_n757), .A3(new_n1001), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n991), .B1(new_n999), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1055), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1026), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n702), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n975), .A2(new_n994), .ZN(new_n1064));
  NAND2_X1  g639(.A1(KEYINPUT53), .A2(G40), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n471), .A2(G2078), .A3(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1064), .A2(new_n976), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(G2078), .B1(new_n996), .B2(new_n998), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1063), .B(new_n1067), .C1(new_n1068), .C2(KEYINPUT53), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1061), .A2(G301), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n1072));
  INV_X1    g647(.A(G2084), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1005), .A2(new_n1073), .A3(new_n1007), .ZN(new_n1074));
  INV_X1    g649(.A(G1966), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n995), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G8), .ZN(new_n1078));
  NAND2_X1  g653(.A1(G286), .A2(G8), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT123), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1080), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1078), .A2(new_n1079), .A3(new_n1083), .ZN(new_n1084));
  OAI211_X1 g659(.A(G8), .B(new_n1082), .C1(new_n1077), .C2(G286), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1079), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1072), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  AOI211_X1 g664(.A(KEYINPUT124), .B(new_n1087), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT62), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OR3_X1    g666(.A1(new_n1089), .A2(new_n1090), .A3(KEYINPUT62), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1071), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1055), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1009), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1024), .A2(new_n1020), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT111), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1024), .A2(new_n1010), .A3(new_n1020), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1095), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  AOI211_X1 g674(.A(new_n991), .B(G286), .C1(new_n1074), .C2(new_n1076), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT63), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1094), .B1(new_n1099), .B2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1094), .B(new_n1100), .C1(new_n1009), .C2(new_n1096), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1106), .A2(new_n1027), .A3(new_n825), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n1043), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1105), .A2(KEYINPUT63), .B1(new_n1030), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1104), .A2(new_n1109), .A3(KEYINPUT114), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1101), .B(new_n1100), .C1(new_n1096), .C2(new_n1058), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1055), .B1(new_n1026), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1108), .A2(new_n1030), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1038), .A2(new_n1100), .A3(new_n1054), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1115), .B1(new_n1056), .B2(new_n1095), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1114), .B1(new_n1116), .B2(new_n1101), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1111), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1068), .A2(KEYINPUT53), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n702), .B2(new_n1062), .ZN(new_n1120));
  NAND2_X1  g695(.A1(G301), .A2(KEYINPUT54), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n1122));
  NAND2_X1  g697(.A1(G171), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n474), .A2(new_n475), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n472), .B1(new_n1124), .B2(KEYINPUT125), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(KEYINPUT125), .B2(new_n1124), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1064), .A2(new_n1066), .A3(new_n1126), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1121), .A2(new_n1123), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1120), .A2(new_n1128), .B1(new_n1069), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(new_n1061), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1133), .A2(KEYINPUT116), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(KEYINPUT116), .ZN(new_n1136));
  NAND3_X1  g711(.A1(G299), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n572), .A2(new_n579), .A3(KEYINPUT116), .A4(new_n1133), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  XOR2_X1   g714(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(G2072), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1064), .A2(new_n993), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT115), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n973), .A2(KEYINPUT50), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1144), .A2(new_n993), .A3(new_n1001), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1143), .B1(new_n1145), .B2(new_n778), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1145), .A2(new_n1143), .A3(new_n778), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1139), .B(new_n1142), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1040), .A2(G2067), .ZN(new_n1149));
  INV_X1    g724(.A(G1348), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1149), .B1(new_n1062), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT118), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(G1348), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT118), .B1(new_n1154), .B2(new_n1149), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1153), .A2(new_n627), .A3(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1142), .B1(new_n1147), .B2(new_n1146), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1148), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(KEYINPUT119), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT119), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1162), .B(new_n1148), .C1(new_n1156), .C2(new_n1159), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT60), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1153), .A2(new_n1164), .A3(new_n1155), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1164), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n618), .A2(KEYINPUT122), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n613), .A2(new_n1169), .A3(new_n617), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  AOI211_X1 g746(.A(new_n1164), .B(new_n1171), .C1(new_n1153), .C2(new_n1155), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1174), .B1(new_n1159), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1148), .A2(new_n1177), .A3(KEYINPUT61), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1040), .ZN(new_n1179));
  XNOR2_X1  g754(.A(KEYINPUT58), .B(G1341), .ZN(new_n1180));
  XNOR2_X1  g755(.A(KEYINPUT120), .B(G1996), .ZN(new_n1181));
  OAI22_X1  g756(.A1(new_n1179), .A2(new_n1180), .B1(new_n995), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT121), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n562), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT59), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1176), .A2(new_n1178), .A3(new_n1185), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1161), .B(new_n1163), .C1(new_n1173), .C2(new_n1186), .ZN(new_n1187));
  AOI22_X1  g762(.A1(new_n1110), .A2(new_n1118), .B1(new_n1132), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1093), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1110), .A2(new_n1118), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1132), .A2(new_n1187), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1191), .A2(new_n1192), .A3(new_n1189), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n990), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n979), .A2(new_n982), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n1195), .B(KEYINPUT46), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n981), .A2(new_n881), .ZN(new_n1197));
  INV_X1    g772(.A(new_n979), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1196), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  XOR2_X1   g774(.A(new_n1199), .B(KEYINPUT127), .Z(new_n1200));
  AND2_X1   g775(.A1(new_n1200), .A2(KEYINPUT47), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1200), .A2(KEYINPUT47), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n987), .A2(new_n1198), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1203), .B(KEYINPUT48), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1204), .B1(new_n986), .B2(new_n979), .ZN(new_n1205));
  INV_X1    g780(.A(new_n845), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n843), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n984), .A2(new_n1207), .ZN(new_n1208));
  OR2_X1    g783(.A1(new_n769), .A2(G2067), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1198), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NOR4_X1   g785(.A1(new_n1201), .A2(new_n1202), .A3(new_n1205), .A4(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1194), .A2(new_n1211), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g787(.A(G319), .ZN(new_n1214));
  NOR4_X1   g788(.A1(G229), .A2(new_n1214), .A3(G401), .A4(G227), .ZN(new_n1215));
  OAI211_X1 g789(.A(new_n910), .B(new_n1215), .C1(new_n968), .C2(new_n969), .ZN(G225));
  INV_X1    g790(.A(G225), .ZN(G308));
endmodule


