//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202));
  OR2_X1    g001(.A1(G71gat), .A2(G78gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G71gat), .A2(G78gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT9), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n202), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G57gat), .B(G64gat), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n204), .B(new_n203), .C1(new_n209), .C2(new_n206), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT21), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XOR2_X1   g012(.A(G127gat), .B(G155gat), .Z(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(G211gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G15gat), .B(G22gat), .ZN(new_n218));
  INV_X1    g017(.A(G1gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT16), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G1gat), .B2(new_n218), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n222), .A2(G8gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(G8gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n211), .A2(new_n212), .ZN(new_n226));
  NOR3_X1   g025(.A1(new_n225), .A2(G183gat), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(G183gat), .B1(new_n225), .B2(new_n226), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n230));
  NAND2_X1  g029(.A1(G231gat), .A2(G233gat), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n230), .B(new_n231), .Z(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n228), .A2(new_n229), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n233), .B1(new_n228), .B2(new_n229), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n217), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n236), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(new_n216), .A3(new_n234), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  AND2_X1   g039(.A1(G232gat), .A2(G233gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n241), .A2(KEYINPUT41), .ZN(new_n242));
  XNOR2_X1  g041(.A(G190gat), .B(G218gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G99gat), .A2(G106gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT8), .ZN(new_n247));
  NAND2_X1  g046(.A1(G85gat), .A2(G92gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT7), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G85gat), .ZN(new_n251));
  INV_X1    g050(.A(G92gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n247), .A2(new_n250), .A3(new_n253), .A4(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G99gat), .B(G106gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT87), .ZN(new_n259));
  AOI22_X1  g058(.A1(KEYINPUT8), .A2(new_n246), .B1(new_n251), .B2(new_n252), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n260), .A2(new_n256), .A3(new_n250), .A4(new_n254), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n255), .A2(KEYINPUT87), .A3(new_n257), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT88), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n262), .A2(KEYINPUT88), .A3(new_n263), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G43gat), .B(G50gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT15), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT14), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n272), .B(KEYINPUT84), .C1(G29gat), .C2(G36gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(G29gat), .A2(G36gat), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n273), .B(new_n274), .C1(new_n269), .C2(KEYINPUT15), .ZN(new_n275));
  OR3_X1    g074(.A1(KEYINPUT84), .A2(G29gat), .A3(G36gat), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT84), .B1(G29gat), .B2(G36gat), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n276), .A2(KEYINPUT14), .A3(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n271), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g078(.A1(G43gat), .A2(G50gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(G43gat), .A2(G50gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT15), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n282), .A2(new_n283), .B1(G29gat), .B2(G36gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n276), .A2(KEYINPUT14), .A3(new_n277), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n284), .A2(new_n270), .A3(new_n285), .A4(new_n273), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n279), .A2(new_n286), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n268), .A2(new_n287), .B1(KEYINPUT41), .B2(new_n241), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n269), .A2(KEYINPUT15), .A3(KEYINPUT17), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT17), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT85), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n292), .B1(new_n287), .B2(new_n293), .ZN(new_n294));
  AOI211_X1 g093(.A(KEYINPUT85), .B(new_n291), .C1(new_n279), .C2(new_n286), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n267), .B(new_n266), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G134gat), .B(G162gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n288), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n298), .B1(new_n288), .B2(new_n296), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n245), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n301), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n303), .A2(new_n299), .A3(new_n244), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n240), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT89), .ZN(new_n306));
  XNOR2_X1  g105(.A(G176gat), .B(G204gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT92), .ZN(new_n308));
  XNOR2_X1  g107(.A(G120gat), .B(G148gat), .ZN(new_n309));
  XOR2_X1   g108(.A(new_n308), .B(new_n309), .Z(new_n310));
  INV_X1    g109(.A(KEYINPUT10), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n211), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n268), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n262), .A2(new_n211), .A3(new_n263), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT90), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT90), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n262), .A2(new_n316), .A3(new_n211), .A4(new_n263), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n208), .A2(new_n210), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n319), .A2(new_n258), .A3(new_n261), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  AND4_X1   g120(.A1(KEYINPUT91), .A2(new_n318), .A3(new_n311), .A4(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n320), .B1(new_n315), .B2(new_n317), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT91), .B1(new_n323), .B2(new_n311), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n313), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G230gat), .A2(G233gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n323), .A2(new_n326), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n310), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n310), .ZN(new_n331));
  AOI211_X1 g130(.A(new_n328), .B(new_n331), .C1(new_n325), .C2(new_n326), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT89), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n240), .A2(new_n302), .A3(new_n334), .A4(new_n304), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n306), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT93), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n306), .A2(new_n333), .A3(KEYINPUT93), .A4(new_n335), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G1gat), .B(G29gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT0), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n343), .B(G57gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(new_n251), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(G155gat), .B(G162gat), .Z(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G155gat), .ZN(new_n349));
  INV_X1    g148(.A(G162gat), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT2), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(G141gat), .B(G148gat), .Z(new_n352));
  NAND3_X1  g151(.A1(new_n348), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n351), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n347), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G113gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(G120gat), .ZN(new_n359));
  INV_X1    g158(.A(G120gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(G113gat), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n359), .B1(KEYINPUT71), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT71), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n363), .B1(new_n360), .B2(G113gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  XOR2_X1   g164(.A(G127gat), .B(G134gat), .Z(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(KEYINPUT1), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT1), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n368), .B1(new_n359), .B2(new_n361), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n365), .A2(new_n367), .B1(new_n369), .B2(new_n366), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n357), .A2(KEYINPUT4), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT4), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n365), .A2(new_n367), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n369), .A2(new_n366), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n372), .B1(new_n375), .B2(new_n356), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT80), .B1(new_n371), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n356), .A2(KEYINPUT3), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n353), .A2(new_n355), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n378), .A2(new_n375), .A3(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(KEYINPUT80), .B(KEYINPUT4), .C1(new_n375), .C2(new_n356), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n377), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G225gat), .A2(G233gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(KEYINPUT79), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT39), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n357), .A2(new_n370), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n356), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n387), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n389), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n346), .B1(new_n388), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n385), .A2(new_n389), .A3(new_n387), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(KEYINPUT40), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n371), .A2(new_n376), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n390), .A2(new_n387), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n381), .ZN(new_n401));
  OAI221_X1 g200(.A(KEYINPUT5), .B1(new_n393), .B2(new_n394), .C1(new_n399), .C2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n387), .A2(KEYINPUT5), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n403), .B1(new_n384), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n404), .ZN(new_n406));
  NOR4_X1   g205(.A1(new_n377), .A2(new_n383), .A3(KEYINPUT81), .A4(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n402), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n346), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n398), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT40), .B1(new_n396), .B2(new_n397), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT22), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT75), .B(G211gat), .ZN(new_n414));
  INV_X1    g213(.A(G218gat), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OR2_X1    g215(.A1(KEYINPUT74), .A2(G204gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(KEYINPUT74), .A2(G204gat), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(G197gat), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n418), .ZN(new_n420));
  INV_X1    g219(.A(G197gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n416), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G211gat), .B(G218gat), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT76), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n416), .A2(new_n424), .A3(new_n419), .A4(new_n422), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n423), .A2(KEYINPUT76), .A3(new_n425), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(KEYINPUT27), .B(G183gat), .ZN(new_n432));
  INV_X1    g231(.A(G190gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n434), .A2(new_n435), .B1(G183gat), .B2(G190gat), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(G169gat), .ZN(new_n438));
  INV_X1    g237(.A(G176gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT26), .ZN(new_n441));
  NAND2_X1  g240(.A1(G169gat), .A2(G176gat), .ZN(new_n442));
  NOR2_X1   g241(.A1(G169gat), .A2(G176gat), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT26), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n434), .B2(new_n435), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n437), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT25), .B1(new_n443), .B2(KEYINPUT23), .ZN(new_n449));
  NAND2_X1  g248(.A1(G183gat), .A2(G190gat), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT66), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT24), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n452), .B1(new_n451), .B2(new_n450), .ZN(new_n453));
  AND3_X1   g252(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n454));
  INV_X1    g253(.A(G183gat), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n454), .B1(new_n455), .B2(new_n433), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n449), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT23), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n442), .B1(new_n440), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT65), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT65), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n461), .B(new_n442), .C1(new_n440), .C2(new_n458), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT67), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n457), .A2(new_n463), .A3(KEYINPUT67), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n459), .B1(new_n458), .B2(new_n440), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT64), .ZN(new_n471));
  OR2_X1    g270(.A1(new_n470), .A2(KEYINPUT64), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT25), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n448), .B1(new_n468), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(G226gat), .A2(G233gat), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n478), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n457), .A2(new_n463), .A3(KEYINPUT67), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT67), .B1(new_n457), .B2(new_n463), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n476), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT68), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g284(.A(KEYINPUT68), .B(new_n476), .C1(new_n481), .C2(new_n482), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT70), .B1(new_n437), .B2(new_n447), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n434), .A2(new_n435), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT70), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n488), .A2(new_n436), .A3(new_n489), .A4(new_n446), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n485), .A2(new_n486), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT29), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n480), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n479), .B1(new_n494), .B2(KEYINPUT77), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n486), .A2(new_n491), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT29), .B1(new_n496), .B2(new_n485), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT77), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n497), .A2(new_n498), .A3(new_n480), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n431), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n478), .B1(new_n477), .B2(KEYINPUT29), .ZN(new_n501));
  INV_X1    g300(.A(new_n492), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n501), .B1(new_n502), .B2(new_n478), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n503), .A2(new_n431), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G8gat), .B(G36gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(G64gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(new_n252), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n500), .A2(new_n505), .A3(KEYINPUT30), .A4(new_n509), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(KEYINPUT78), .B(KEYINPUT30), .Z(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n498), .B1(new_n497), .B2(new_n480), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n494), .A2(KEYINPUT77), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(new_n479), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n504), .B1(new_n518), .B2(new_n431), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n515), .B1(new_n519), .B2(new_n509), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n412), .B1(new_n513), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT29), .B1(new_n426), .B2(new_n428), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n356), .B1(new_n522), .B2(KEYINPUT3), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n429), .A2(new_n430), .B1(new_n493), .B2(new_n380), .ZN(new_n525));
  INV_X1    g324(.A(G228gat), .ZN(new_n526));
  INV_X1    g325(.A(G233gat), .ZN(new_n527));
  OAI22_X1  g326(.A1(new_n524), .A2(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G22gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n429), .A2(new_n493), .A3(new_n430), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n357), .B1(new_n530), .B2(new_n379), .ZN(new_n531));
  INV_X1    g330(.A(new_n525), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n526), .A2(new_n527), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n528), .B(new_n529), .C1(new_n531), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT82), .ZN(new_n536));
  XNOR2_X1  g335(.A(G78gat), .B(G106gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT31), .B(G50gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n534), .A2(new_n531), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n533), .B1(new_n532), .B2(new_n523), .ZN(new_n541));
  OAI21_X1  g340(.A(G22gat), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n536), .A2(new_n539), .B1(new_n542), .B2(new_n535), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT82), .ZN(new_n544));
  AND4_X1   g343(.A1(new_n544), .A2(new_n542), .A3(new_n535), .A4(new_n539), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT38), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT37), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n506), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n519), .A2(KEYINPUT37), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n547), .B1(new_n551), .B2(new_n510), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n509), .A2(KEYINPUT38), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT37), .B1(new_n500), .B2(new_n505), .ZN(new_n554));
  INV_X1    g353(.A(new_n431), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n516), .A2(new_n517), .A3(new_n555), .A4(new_n479), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n548), .B1(new_n503), .B2(new_n431), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n553), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT6), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n402), .B(new_n345), .C1(new_n405), .C2(new_n407), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n409), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n408), .A2(KEYINPUT6), .A3(new_n346), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n519), .A2(new_n509), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n559), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n521), .B(new_n546), .C1(new_n552), .C2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n543), .A2(new_n545), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n514), .B1(new_n506), .B2(new_n510), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n570), .A2(new_n564), .A3(new_n511), .A4(new_n512), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n486), .A2(new_n491), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT68), .B1(new_n468), .B2(new_n476), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n370), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G227gat), .A2(G233gat), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n485), .A2(new_n375), .A3(new_n486), .A4(new_n491), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT32), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT33), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G15gat), .B(G43gat), .Z(new_n582));
  XNOR2_X1  g381(.A(G71gat), .B(G99gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n579), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n584), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n578), .B(KEYINPUT32), .C1(new_n580), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n574), .A2(new_n577), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n575), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT34), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n590), .A2(KEYINPUT73), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n576), .B1(new_n574), .B2(new_n577), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT73), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT34), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT72), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n592), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n588), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n588), .A2(new_n597), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT36), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n592), .A2(new_n595), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n588), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT36), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n585), .A2(new_n595), .A3(new_n592), .A4(new_n587), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AOI22_X1  g404(.A1(new_n569), .A2(new_n571), .B1(new_n600), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n568), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n513), .A2(new_n520), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT35), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n569), .B1(new_n604), .B2(new_n602), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n564), .A4(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n546), .B1(new_n598), .B2(new_n599), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT35), .B1(new_n571), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n607), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT86), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n223), .A2(new_n224), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n617), .B1(new_n294), .B2(new_n295), .ZN(new_n618));
  NAND2_X1  g417(.A1(G229gat), .A2(G233gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n225), .A2(new_n287), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT18), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n225), .B(new_n287), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n619), .B(KEYINPUT13), .Z(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n618), .A2(KEYINPUT18), .A3(new_n619), .A4(new_n620), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n623), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT83), .ZN(new_n629));
  XNOR2_X1  g428(.A(G113gat), .B(G141gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT11), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(new_n438), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G197gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n634), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n636), .A2(new_n628), .A3(KEYINPUT83), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n615), .A2(new_n616), .A3(new_n638), .ZN(new_n639));
  AOI22_X1  g438(.A1(new_n568), .A2(new_n606), .B1(new_n611), .B2(new_n613), .ZN(new_n640));
  INV_X1    g439(.A(new_n638), .ZN(new_n641));
  OAI21_X1  g440(.A(KEYINPUT86), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n341), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n565), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g444(.A1(new_n639), .A2(new_n642), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n570), .A2(new_n511), .A3(new_n512), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT16), .B(G8gat), .Z(new_n648));
  NAND4_X1  g447(.A1(new_n646), .A2(new_n647), .A3(new_n340), .A4(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT42), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n643), .A2(KEYINPUT42), .A3(new_n647), .A4(new_n648), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n646), .A2(new_n647), .A3(new_n340), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(G8gat), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n651), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT94), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n651), .A2(new_n654), .A3(new_n652), .A4(KEYINPUT94), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(G1325gat));
  INV_X1    g458(.A(G15gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n602), .A2(new_n604), .ZN(new_n661));
  AND4_X1   g460(.A1(new_n660), .A2(new_n646), .A3(new_n661), .A4(new_n340), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n600), .A2(new_n605), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n660), .B1(new_n643), .B2(new_n664), .ZN(new_n665));
  OR3_X1    g464(.A1(new_n662), .A2(new_n665), .A3(KEYINPUT95), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT95), .B1(new_n662), .B2(new_n665), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(G1326gat));
  NAND2_X1  g467(.A1(new_n643), .A2(new_n569), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT43), .B(G22gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT96), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n669), .B(new_n671), .ZN(G1327gat));
  INV_X1    g471(.A(new_n240), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n333), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n304), .A2(new_n302), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n646), .A2(new_n677), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n678), .A2(G29gat), .A3(new_n564), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n679), .A2(KEYINPUT45), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n674), .A2(new_n641), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n615), .A2(new_n683), .A3(new_n675), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT44), .B1(new_n640), .B2(new_n676), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n682), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(G29gat), .B1(new_n687), .B2(new_n564), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n679), .A2(KEYINPUT45), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n680), .A2(new_n688), .A3(new_n689), .ZN(G1328gat));
  NOR2_X1   g489(.A1(new_n608), .A2(G36gat), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n646), .A2(new_n677), .A3(new_n691), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n692), .A2(KEYINPUT46), .ZN(new_n693));
  OAI21_X1  g492(.A(G36gat), .B1(new_n687), .B2(new_n608), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(KEYINPUT46), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(G1329gat));
  INV_X1    g495(.A(KEYINPUT97), .ZN(new_n697));
  INV_X1    g496(.A(G43gat), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n661), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n697), .B1(new_n678), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT47), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n678), .A2(new_n699), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n698), .B1(new_n686), .B2(new_n664), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n700), .B(new_n701), .C1(new_n703), .C2(new_n704), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(G1330gat));
  INV_X1    g507(.A(G50gat), .ZN(new_n709));
  AND4_X1   g508(.A1(new_n709), .A2(new_n646), .A3(new_n569), .A4(new_n677), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n709), .B1(new_n686), .B2(new_n569), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT98), .B(KEYINPUT48), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  OR3_X1    g512(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n710), .B2(new_n711), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(G1331gat));
  INV_X1    g515(.A(new_n333), .ZN(new_n717));
  AND4_X1   g516(.A1(new_n641), .A2(new_n717), .A3(new_n306), .A4(new_n335), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n615), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n565), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g521(.A(new_n608), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(new_n728), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(G1333gat));
  INV_X1    g530(.A(G71gat), .ZN(new_n732));
  INV_X1    g531(.A(new_n661), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n719), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT101), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n663), .A2(new_n732), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n735), .B1(new_n720), .B2(new_n736), .ZN(new_n737));
  NOR4_X1   g536(.A1(new_n719), .A2(KEYINPUT101), .A3(new_n732), .A4(new_n663), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n734), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g539(.A1(new_n719), .A2(new_n546), .ZN(new_n741));
  XNOR2_X1  g540(.A(KEYINPUT102), .B(G78gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1335gat));
  NOR2_X1   g542(.A1(new_n638), .A2(new_n240), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n615), .A2(new_n675), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n333), .B1(new_n745), .B2(KEYINPUT51), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n615), .A2(new_n747), .A3(new_n675), .A4(new_n744), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n749), .A2(new_n251), .A3(new_n565), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n744), .A2(new_n717), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT103), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n683), .B1(new_n615), .B2(new_n675), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n640), .A2(KEYINPUT44), .A3(new_n676), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(G85gat), .B1(new_n755), .B2(new_n564), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n750), .A2(new_n756), .ZN(G1336gat));
  INV_X1    g556(.A(KEYINPUT104), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n758), .A2(KEYINPUT52), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(KEYINPUT52), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n608), .A2(G92gat), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n748), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n752), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n764), .B1(new_n684), .B2(new_n685), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n252), .B1(new_n765), .B2(new_n647), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n759), .B(new_n760), .C1(new_n763), .C2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G92gat), .B1(new_n755), .B2(new_n608), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n768), .A2(new_n758), .A3(KEYINPUT52), .A4(new_n762), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n767), .A2(new_n769), .ZN(G1337gat));
  INV_X1    g569(.A(G99gat), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n755), .A2(new_n771), .A3(new_n663), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n749), .A2(new_n661), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n772), .B1(new_n773), .B2(new_n771), .ZN(G1338gat));
  OAI211_X1 g573(.A(new_n569), .B(new_n752), .C1(new_n753), .C2(new_n754), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT105), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n775), .A2(new_n776), .A3(G106gat), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n546), .A2(G106gat), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n746), .A2(KEYINPUT106), .A3(new_n748), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n776), .B1(new_n775), .B2(G106gat), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT53), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n749), .A2(new_n778), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n775), .A2(new_n784), .A3(G106gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(KEYINPUT106), .A2(KEYINPUT53), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n783), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n782), .A2(new_n787), .ZN(G1339gat));
  NOR2_X1   g587(.A1(new_n336), .A2(new_n638), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n636), .A2(new_n628), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n619), .B1(new_n618), .B2(new_n620), .ZN(new_n792));
  OAI22_X1  g591(.A1(new_n792), .A2(KEYINPUT107), .B1(new_n624), .B2(new_n625), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n792), .A2(KEYINPUT107), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n633), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n318), .A2(new_n311), .A3(new_n321), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT91), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n323), .A2(KEYINPUT91), .A3(new_n311), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n326), .B1(new_n268), .B2(new_n312), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n798), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n797), .B1(new_n805), .B2(new_n327), .ZN(new_n806));
  INV_X1    g605(.A(new_n326), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n807), .B1(new_n803), .B2(new_n313), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n310), .B1(new_n808), .B2(new_n798), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n332), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n804), .B1(new_n322), .B2(new_n324), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT54), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n325), .A2(new_n798), .A3(new_n326), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n331), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n797), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n796), .A2(new_n810), .A3(new_n675), .A4(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n810), .A2(new_n816), .A3(new_n638), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n791), .B(new_n795), .C1(new_n330), .C2(new_n332), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT108), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n675), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n819), .A2(KEYINPUT108), .A3(new_n820), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n818), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n790), .B1(new_n825), .B2(new_n240), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n826), .A2(new_n610), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n647), .A2(new_n564), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n829), .A2(new_n358), .A3(new_n641), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n819), .A2(KEYINPUT108), .A3(new_n820), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT108), .B1(new_n819), .B2(new_n820), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n831), .A2(new_n832), .A3(new_n675), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n673), .B1(new_n833), .B2(new_n818), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n564), .B1(new_n834), .B2(new_n790), .ZN(new_n835));
  INV_X1    g634(.A(new_n612), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(new_n608), .A3(new_n638), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n830), .B1(new_n839), .B2(new_n358), .ZN(G1340gat));
  NOR3_X1   g639(.A1(new_n829), .A2(new_n360), .A3(new_n333), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n838), .A2(new_n608), .A3(new_n717), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(new_n842), .B2(new_n360), .ZN(G1341gat));
  NAND4_X1  g642(.A1(new_n827), .A2(G127gat), .A3(new_n240), .A4(new_n828), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT109), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n838), .A2(new_n608), .A3(new_n240), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n847), .A2(KEYINPUT110), .ZN(new_n848));
  AOI21_X1  g647(.A(G127gat), .B1(new_n847), .B2(KEYINPUT110), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(G1342gat));
  NAND2_X1  g649(.A1(new_n608), .A2(new_n675), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT111), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n852), .A2(G134gat), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT56), .B1(new_n837), .B2(new_n853), .ZN(new_n854));
  OR3_X1    g653(.A1(new_n837), .A2(KEYINPUT56), .A3(new_n853), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n827), .A2(new_n675), .A3(new_n828), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n856), .A2(KEYINPUT112), .A3(G134gat), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT112), .B1(new_n856), .B2(G134gat), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n854), .B(new_n855), .C1(new_n857), .C2(new_n858), .ZN(G1343gat));
  NAND4_X1  g658(.A1(new_n826), .A2(new_n565), .A3(new_n569), .A4(new_n663), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n860), .A2(new_n647), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n641), .A2(G141gat), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT113), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n861), .A2(KEYINPUT113), .A3(new_n862), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n826), .A2(new_n867), .A3(new_n569), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n828), .A2(new_n663), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n821), .A2(new_n676), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n817), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n673), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n546), .B1(new_n873), .B2(new_n790), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n868), .B(new_n870), .C1(new_n867), .C2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(G141gat), .B1(new_n875), .B2(new_n641), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n865), .A2(new_n866), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT58), .ZN(new_n878));
  XNOR2_X1  g677(.A(KEYINPUT114), .B(KEYINPUT58), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n876), .A2(new_n863), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(G1344gat));
  INV_X1    g680(.A(G148gat), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n861), .A2(new_n882), .A3(new_n717), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n875), .A2(new_n333), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n884), .A2(KEYINPUT59), .A3(new_n882), .ZN(new_n885));
  XNOR2_X1  g684(.A(KEYINPUT115), .B(KEYINPUT59), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n826), .A2(new_n569), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT57), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n638), .B1(new_n338), .B2(new_n339), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT116), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n873), .A3(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n546), .A2(KEYINPUT57), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n888), .A2(new_n717), .A3(new_n870), .A4(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n886), .B1(new_n896), .B2(G148gat), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n883), .B1(new_n885), .B2(new_n897), .ZN(G1345gat));
  OAI21_X1  g697(.A(G155gat), .B1(new_n875), .B2(new_n673), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n861), .A2(new_n349), .A3(new_n240), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(G1346gat));
  OAI21_X1  g700(.A(G162gat), .B1(new_n875), .B2(new_n676), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n852), .A2(G162gat), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n860), .B2(new_n903), .ZN(G1347gat));
  NOR2_X1   g703(.A1(new_n608), .A2(new_n565), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n827), .A2(new_n638), .A3(new_n905), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n906), .A2(KEYINPUT117), .A3(G169gat), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT117), .B1(new_n906), .B2(G169gat), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n565), .B1(new_n834), .B2(new_n790), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n647), .A3(new_n836), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n638), .A2(new_n438), .ZN(new_n911));
  OAI22_X1  g710(.A1(new_n907), .A2(new_n908), .B1(new_n910), .B2(new_n911), .ZN(G1348gat));
  NAND2_X1  g711(.A1(new_n827), .A2(new_n905), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n333), .A2(new_n439), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT118), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n439), .B1(new_n910), .B2(new_n333), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n913), .A2(KEYINPUT118), .A3(new_n915), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(G1349gat));
  NOR2_X1   g719(.A1(KEYINPUT119), .A2(KEYINPUT60), .ZN(new_n921));
  AND2_X1   g720(.A1(KEYINPUT119), .A2(KEYINPUT60), .ZN(new_n922));
  INV_X1    g721(.A(new_n910), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n432), .A3(new_n240), .ZN(new_n924));
  OAI21_X1  g723(.A(G183gat), .B1(new_n913), .B2(new_n673), .ZN(new_n925));
  AOI211_X1 g724(.A(new_n921), .B(new_n922), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  AND4_X1   g725(.A1(KEYINPUT119), .A2(new_n924), .A3(KEYINPUT60), .A4(new_n925), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(G1350gat));
  NOR3_X1   g727(.A1(new_n910), .A2(G190gat), .A3(new_n676), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT120), .ZN(new_n930));
  OAI21_X1  g729(.A(G190gat), .B1(new_n913), .B2(new_n676), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n930), .A2(new_n933), .A3(new_n934), .ZN(G1351gat));
  AND2_X1   g734(.A1(new_n592), .A2(new_n595), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n936), .A2(new_n596), .A3(new_n587), .A4(new_n585), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n588), .A2(new_n597), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n603), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n647), .B(new_n569), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT121), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n826), .A2(new_n942), .A3(new_n564), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT122), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n909), .A2(new_n945), .A3(new_n942), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n638), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT123), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n867), .B1(new_n826), .B2(new_n569), .ZN(new_n950));
  INV_X1    g749(.A(new_n894), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n889), .B(KEYINPUT116), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n951), .B1(new_n952), .B2(new_n873), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n949), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n546), .B1(new_n834), .B2(new_n790), .ZN(new_n955));
  OAI211_X1 g754(.A(KEYINPUT123), .B(new_n895), .C1(new_n955), .C2(new_n867), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n905), .A2(new_n663), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n958), .A2(new_n421), .A3(new_n641), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n948), .B1(new_n957), .B2(new_n959), .ZN(G1352gat));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n961));
  OR2_X1    g760(.A1(new_n961), .A2(KEYINPUT124), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(KEYINPUT124), .ZN(new_n963));
  INV_X1    g762(.A(G204gat), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n717), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n962), .B(new_n963), .C1(new_n943), .C2(new_n965), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n943), .A2(new_n965), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n967), .B2(new_n962), .ZN(new_n968));
  INV_X1    g767(.A(new_n958), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(new_n717), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n970), .B1(new_n954), .B2(new_n956), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n968), .B1(new_n971), .B2(new_n964), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(KEYINPUT125), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT125), .ZN(new_n974));
  OAI211_X1 g773(.A(new_n968), .B(new_n974), .C1(new_n971), .C2(new_n964), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n975), .ZN(G1353gat));
  NAND3_X1  g775(.A1(new_n947), .A2(new_n414), .A3(new_n240), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n958), .A2(new_n673), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n888), .A2(new_n895), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(KEYINPUT126), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT126), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n888), .A2(new_n981), .A3(new_n895), .A4(new_n978), .ZN(new_n982));
  AND4_X1   g781(.A1(KEYINPUT63), .A2(new_n980), .A3(G211gat), .A4(new_n982), .ZN(new_n983));
  INV_X1    g782(.A(G211gat), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n984), .B1(new_n979), .B2(KEYINPUT126), .ZN(new_n985));
  AOI21_X1  g784(.A(KEYINPUT63), .B1(new_n985), .B2(new_n982), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n977), .B1(new_n983), .B2(new_n986), .ZN(G1354gat));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n944), .A2(new_n946), .A3(new_n675), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(new_n415), .ZN(new_n990));
  INV_X1    g789(.A(new_n990), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n676), .A2(new_n415), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n969), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n993), .B1(new_n954), .B2(new_n956), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n988), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  INV_X1    g794(.A(new_n994), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n996), .A2(KEYINPUT127), .A3(new_n990), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n995), .A2(new_n997), .ZN(G1355gat));
endmodule


