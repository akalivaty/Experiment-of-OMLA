//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958;
  XNOR2_X1  g000(.A(KEYINPUT69), .B(G113gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G120gat), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  INV_X1    g003(.A(G120gat), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT1), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G127gat), .B(G134gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n203), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT70), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n203), .A2(KEYINPUT70), .A3(new_n206), .A4(new_n207), .ZN(new_n211));
  NAND2_X1  g010(.A1(G113gat), .A2(G120gat), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n207), .B1(new_n212), .B2(new_n206), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT68), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT68), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n206), .A2(new_n212), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(new_n207), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n210), .A2(new_n211), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G169gat), .ZN(new_n219));
  INV_X1    g018(.A(G176gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  NOR3_X1   g021(.A1(new_n221), .A2(KEYINPUT26), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G183gat), .ZN(new_n224));
  INV_X1    g023(.A(G190gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n222), .A2(KEYINPUT26), .ZN(new_n227));
  NOR3_X1   g026(.A1(new_n223), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT27), .B(G183gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(KEYINPUT28), .A3(new_n225), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT28), .ZN(new_n233));
  NOR2_X1   g032(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT65), .B(G183gat), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n234), .B1(new_n235), .B2(KEYINPUT27), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n233), .B1(new_n236), .B2(G190gat), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n232), .B1(new_n237), .B2(KEYINPUT67), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n239), .B(new_n233), .C1(new_n236), .C2(G190gat), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n229), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT24), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(G183gat), .A3(G190gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n243), .B1(new_n226), .B2(new_n242), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(G190gat), .B2(new_n235), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n235), .A2(G190gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n248), .A2(KEYINPUT66), .A3(new_n244), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  OR2_X1    g049(.A1(new_n222), .A2(KEYINPUT23), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n222), .A2(KEYINPUT23), .ZN(new_n252));
  INV_X1    g051(.A(new_n221), .ZN(new_n253));
  AND4_X1   g052(.A1(KEYINPUT25), .A2(new_n251), .A3(new_n252), .A4(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT25), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT64), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n256), .B1(G183gat), .B2(G190gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT64), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n244), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n259), .A2(new_n252), .A3(new_n253), .A4(new_n251), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n250), .A2(new_n254), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n218), .B1(new_n241), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n237), .A2(KEYINPUT67), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n263), .A2(new_n240), .A3(new_n231), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(new_n228), .ZN(new_n265));
  INV_X1    g064(.A(new_n218), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n245), .A2(new_n246), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT66), .B1(new_n248), .B2(new_n244), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n254), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n260), .A2(new_n255), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n265), .A2(new_n266), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G227gat), .ZN(new_n273));
  INV_X1    g072(.A(G233gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n262), .A2(new_n272), .A3(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(KEYINPUT71), .B(KEYINPUT33), .Z(new_n277));
  XNOR2_X1  g076(.A(G15gat), .B(G43gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(G71gat), .B(G99gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n276), .B(KEYINPUT32), .C1(new_n277), .C2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n280), .B1(new_n276), .B2(KEYINPUT32), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n276), .A2(new_n277), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n283), .B1(new_n282), .B2(new_n284), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n281), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT34), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n262), .A2(new_n272), .ZN(new_n289));
  INV_X1    g088(.A(new_n275), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI211_X1 g090(.A(KEYINPUT34), .B(new_n275), .C1(new_n262), .C2(new_n272), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n287), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n293), .B(new_n281), .C1(new_n285), .C2(new_n286), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  OR3_X1    g097(.A1(new_n287), .A2(new_n297), .A3(new_n294), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT36), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT74), .A4(new_n300), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n295), .A2(new_n296), .A3(KEYINPUT36), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G155gat), .B(G162gat), .ZN(new_n307));
  XOR2_X1   g106(.A(G141gat), .B(G148gat), .Z(new_n308));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT2), .ZN(new_n311));
  INV_X1    g110(.A(G155gat), .ZN(new_n312));
  INV_X1    g111(.A(G162gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n308), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  OAI221_X1 g115(.A(new_n308), .B1(new_n311), .B2(new_n314), .C1(new_n309), .C2(new_n307), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT77), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n316), .A2(KEYINPUT77), .A3(new_n317), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(KEYINPUT4), .A3(new_n218), .ZN(new_n323));
  NAND2_X1  g122(.A1(G225gat), .A2(G233gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n210), .A2(new_n211), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n214), .A2(new_n217), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n325), .A2(new_n326), .B1(new_n318), .B2(KEYINPUT3), .ZN(new_n327));
  INV_X1    g126(.A(new_n318), .ZN(new_n328));
  XOR2_X1   g127(.A(KEYINPUT76), .B(KEYINPUT3), .Z(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n218), .A2(new_n328), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT4), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n323), .A2(new_n324), .A3(new_n331), .A4(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT78), .B(KEYINPUT5), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n218), .B(new_n328), .ZN(new_n337));
  INV_X1    g136(.A(new_n324), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n336), .ZN(new_n341));
  AOI211_X1 g140(.A(new_n338), .B(new_n341), .C1(new_n327), .C2(new_n330), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n332), .A2(KEYINPUT4), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n320), .A2(new_n218), .A3(new_n333), .A4(new_n321), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n342), .A2(KEYINPUT79), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT79), .B1(new_n342), .B2(new_n345), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n340), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G1gat), .B(G29gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(KEYINPUT0), .ZN(new_n350));
  XNOR2_X1  g149(.A(G57gat), .B(G85gat), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n350), .B(new_n351), .Z(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n340), .B(new_n352), .C1(new_n346), .C2(new_n347), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n356), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n348), .A2(new_n353), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G226gat), .A2(G233gat), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n264), .A2(new_n228), .B1(new_n269), .B2(new_n270), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n360), .B1(new_n361), .B2(KEYINPUT29), .ZN(new_n362));
  OAI211_X1 g161(.A(G226gat), .B(G233gat), .C1(new_n241), .C2(new_n261), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G197gat), .B(G204gat), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT22), .ZN(new_n366));
  INV_X1    g165(.A(G211gat), .ZN(new_n367));
  INV_X1    g166(.A(G218gat), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  XOR2_X1   g169(.A(G211gat), .B(G218gat), .Z(new_n371));
  XOR2_X1   g170(.A(new_n370), .B(new_n371), .Z(new_n372));
  NAND2_X1  g171(.A1(new_n364), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n372), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n362), .A2(new_n374), .A3(new_n363), .ZN(new_n375));
  XNOR2_X1  g174(.A(G8gat), .B(G36gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(G64gat), .B(G92gat), .ZN(new_n377));
  XOR2_X1   g176(.A(new_n376), .B(new_n377), .Z(new_n378));
  NAND3_X1  g177(.A1(new_n373), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n357), .A2(new_n359), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n373), .A2(new_n375), .ZN(new_n382));
  XOR2_X1   g181(.A(KEYINPUT87), .B(KEYINPUT37), .Z(new_n383));
  OAI21_X1  g182(.A(KEYINPUT88), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT88), .ZN(new_n385));
  INV_X1    g184(.A(new_n383), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n373), .A2(new_n385), .A3(new_n375), .A4(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n378), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n375), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n374), .B1(new_n362), .B2(new_n363), .ZN(new_n390));
  OR3_X1    g189(.A1(new_n389), .A2(KEYINPUT86), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT37), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n392), .B1(new_n389), .B2(KEYINPUT86), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT38), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n388), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n382), .A2(KEYINPUT37), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n388), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT38), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n381), .B(new_n395), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT29), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT3), .B1(new_n374), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n401), .A2(new_n328), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n330), .A2(new_n400), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n403), .A2(KEYINPUT82), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n374), .B1(new_n403), .B2(KEYINPUT82), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n402), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(G228gat), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n406), .A2(new_n407), .A3(new_n274), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n274), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n372), .A2(KEYINPUT81), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n370), .A2(new_n371), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n410), .B(new_n400), .C1(KEYINPUT81), .C2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n322), .B1(new_n412), .B2(new_n329), .ZN(new_n413));
  AOI211_X1 g212(.A(new_n409), .B(new_n413), .C1(new_n372), .C2(new_n403), .ZN(new_n414));
  XNOR2_X1  g213(.A(G78gat), .B(G106gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT31), .B(G50gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n417), .A2(G22gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(KEYINPUT83), .A2(G22gat), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n418), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  OR3_X1    g220(.A1(new_n408), .A2(new_n414), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n421), .B1(new_n408), .B2(new_n414), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT39), .B1(new_n337), .B2(new_n338), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT84), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(KEYINPUT84), .B(KEYINPUT39), .C1(new_n337), .C2(new_n338), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n345), .A2(new_n331), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n427), .B(new_n428), .C1(new_n429), .C2(new_n324), .ZN(new_n430));
  OR2_X1    g229(.A1(KEYINPUT85), .A2(KEYINPUT40), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n324), .B1(new_n345), .B2(new_n331), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT39), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n353), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n430), .A2(new_n431), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n354), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n431), .B1(new_n430), .B2(new_n434), .ZN(new_n437));
  NOR3_X1   g236(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n378), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n439), .B1(new_n389), .B2(new_n390), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n440), .A2(KEYINPUT30), .A3(new_n379), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT30), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n373), .A2(new_n442), .A3(new_n375), .A4(new_n378), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n424), .B1(new_n438), .B2(new_n445), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n357), .A2(new_n359), .B1(new_n441), .B2(new_n443), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n399), .A2(new_n446), .B1(new_n448), .B2(new_n424), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n306), .A2(new_n449), .ZN(new_n450));
  NOR3_X1   g249(.A1(new_n448), .A2(KEYINPUT35), .A3(new_n424), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n298), .A2(new_n299), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n422), .A2(new_n423), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n447), .A2(new_n454), .A3(new_n295), .A4(new_n296), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n455), .A2(KEYINPUT89), .A3(KEYINPUT35), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT89), .B1(new_n455), .B2(KEYINPUT35), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n453), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n450), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G134gat), .B(G162gat), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n462), .B(KEYINPUT101), .Z(new_n463));
  INV_X1    g262(.A(G29gat), .ZN(new_n464));
  INV_X1    g263(.A(G36gat), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT14), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT14), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n467), .B1(G29gat), .B2(G36gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(G29gat), .A2(G36gat), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT15), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT15), .A4(new_n469), .ZN(new_n473));
  XNOR2_X1  g272(.A(G43gat), .B(G50gat), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n473), .A2(new_n474), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT17), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT91), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n475), .A2(KEYINPUT91), .A3(new_n476), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT17), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n479), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT97), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT96), .ZN(new_n488));
  AND2_X1   g287(.A1(KEYINPUT95), .A2(G85gat), .ZN(new_n489));
  NOR2_X1   g288(.A1(KEYINPUT95), .A2(G85gat), .ZN(new_n490));
  NOR3_X1   g289(.A1(new_n489), .A2(new_n490), .A3(G92gat), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT8), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n492), .B1(G99gat), .B2(G106gat), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n488), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  OR2_X1    g293(.A1(KEYINPUT95), .A2(G85gat), .ZN(new_n495));
  INV_X1    g294(.A(G92gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(KEYINPUT95), .A2(G85gat), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(G99gat), .ZN(new_n499));
  INV_X1    g298(.A(G106gat), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT8), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n498), .A2(KEYINPUT96), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n494), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G85gat), .A2(G92gat), .ZN(new_n504));
  XOR2_X1   g303(.A(new_n504), .B(KEYINPUT7), .Z(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n487), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  AOI211_X1 g306(.A(KEYINPUT97), .B(new_n505), .C1(new_n494), .C2(new_n502), .ZN(new_n508));
  XOR2_X1   g307(.A(G99gat), .B(G106gat), .Z(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NOR3_X1   g309(.A1(new_n507), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n498), .A2(KEYINPUT96), .A3(new_n501), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT96), .B1(new_n498), .B2(new_n501), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n506), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT97), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n503), .A2(new_n487), .A3(new_n506), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n509), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT98), .B1(new_n511), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n510), .B1(new_n507), .B2(new_n508), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT98), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n515), .A2(new_n509), .A3(new_n516), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n486), .A2(new_n518), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n482), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT91), .B1(new_n475), .B2(new_n476), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n519), .A2(new_n526), .A3(new_n521), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT99), .ZN(new_n528));
  NAND3_X1  g327(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n528), .B1(new_n527), .B2(new_n529), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n523), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT100), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT100), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n523), .B(new_n534), .C1(new_n530), .C2(new_n531), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n533), .A2(new_n225), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n225), .B1(new_n533), .B2(new_n535), .ZN(new_n537));
  NOR3_X1   g336(.A1(new_n536), .A2(new_n537), .A3(G218gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n531), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n534), .B1(new_n541), .B2(new_n523), .ZN(new_n542));
  INV_X1    g341(.A(new_n535), .ZN(new_n543));
  OAI21_X1  g342(.A(G190gat), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n533), .A2(new_n225), .A3(new_n535), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n368), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n463), .B1(new_n538), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(G218gat), .B1(new_n536), .B2(new_n537), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n544), .A2(new_n368), .A3(new_n545), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n462), .A2(KEYINPUT101), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(G57gat), .B(G64gat), .Z(new_n553));
  INV_X1    g352(.A(KEYINPUT9), .ZN(new_n554));
  INV_X1    g353(.A(G71gat), .ZN(new_n555));
  INV_X1    g354(.A(G78gat), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G71gat), .B(G78gat), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n553), .A2(new_n559), .A3(new_n557), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT21), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G127gat), .ZN(new_n568));
  INV_X1    g367(.A(G8gat), .ZN(new_n569));
  INV_X1    g368(.A(G1gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(G15gat), .B(G22gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT92), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n571), .A2(new_n572), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n570), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n575), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n570), .A2(KEYINPUT16), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(new_n578), .A3(new_n573), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n569), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n576), .A2(new_n579), .A3(new_n569), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT94), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n563), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n561), .A2(KEYINPUT94), .A3(new_n562), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n584), .B1(new_n588), .B2(new_n564), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n568), .B(new_n589), .Z(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(G155gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(G183gat), .B(G211gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n590), .B(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G120gat), .B(G148gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT103), .ZN(new_n597));
  XOR2_X1   g396(.A(G176gat), .B(G204gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G230gat), .A2(G233gat), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n601), .B(KEYINPUT104), .Z(new_n602));
  INV_X1    g401(.A(KEYINPUT10), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n603), .B1(new_n586), .B2(new_n587), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n519), .A2(new_n521), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT102), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT102), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n519), .A2(new_n604), .A3(new_n521), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n563), .B1(new_n511), .B2(new_n517), .ZN(new_n610));
  INV_X1    g409(.A(new_n563), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n519), .A2(new_n611), .A3(new_n521), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n603), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n602), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n601), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n519), .A2(new_n611), .A3(new_n521), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n611), .B1(new_n519), .B2(new_n521), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n600), .B1(new_n615), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n600), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n609), .A2(new_n613), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n621), .B1(new_n601), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n552), .A2(new_n595), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n583), .A2(new_n526), .ZN(new_n626));
  NAND2_X1  g425(.A1(G229gat), .A2(G233gat), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n626), .B(new_n627), .C1(new_n485), .C2(new_n583), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT93), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT18), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT18), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n628), .A2(KEYINPUT93), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n584), .A2(new_n483), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n626), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n627), .B(KEYINPUT13), .Z(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n630), .A2(new_n632), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G113gat), .B(G141gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT90), .B(G197gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT11), .B(G169gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n642), .B(KEYINPUT12), .Z(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n637), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n630), .A2(new_n632), .A3(new_n636), .A4(new_n643), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n625), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n459), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n357), .A2(new_n359), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g454(.A1(new_n651), .A2(new_n445), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT105), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(G8gat), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT16), .B(G8gat), .Z(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT42), .ZN(new_n660));
  INV_X1    g459(.A(new_n659), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  OAI221_X1 g461(.A(new_n658), .B1(new_n656), .B2(new_n660), .C1(new_n662), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g462(.A(G15gat), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n651), .A2(new_n664), .A3(new_n452), .ZN(new_n665));
  INV_X1    g464(.A(new_n305), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n666), .B1(new_n301), .B2(new_n302), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n667), .A2(KEYINPUT106), .A3(new_n304), .ZN(new_n668));
  AOI21_X1  g467(.A(KEYINPUT106), .B1(new_n667), .B2(new_n304), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(G15gat), .B1(new_n650), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n665), .A2(new_n671), .ZN(G1326gat));
  NAND2_X1  g471(.A1(new_n651), .A2(new_n424), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT107), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT43), .B(G22gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1327gat));
  OR2_X1    g475(.A1(new_n620), .A2(new_n623), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n595), .A2(new_n648), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n552), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n306), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n667), .A2(KEYINPUT106), .A3(new_n304), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n381), .A2(new_n395), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n398), .B1(new_n388), .B2(new_n396), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n446), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OR3_X1    g486(.A1(new_n447), .A2(new_n454), .A3(KEYINPUT108), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT108), .B1(new_n447), .B2(new_n454), .ZN(new_n689));
  AND3_X1   g488(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n683), .A2(new_n684), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n681), .B1(new_n691), .B2(new_n458), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n680), .B1(new_n459), .B2(new_n679), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n653), .B(new_n678), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n464), .B1(new_n694), .B2(KEYINPUT109), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n692), .A2(new_n693), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n696), .A2(new_n697), .A3(new_n653), .A4(new_n678), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n552), .B1(new_n450), .B2(new_n458), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n678), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n653), .A2(new_n464), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(KEYINPUT45), .Z(new_n704));
  NAND2_X1  g503(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT110), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT110), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n699), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(G1328gat));
  AND2_X1   g508(.A1(new_n696), .A2(new_n678), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n465), .B1(new_n710), .B2(new_n445), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n701), .A2(G36gat), .A3(new_n444), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT46), .Z(new_n713));
  OR2_X1    g512(.A1(new_n711), .A2(new_n713), .ZN(G1329gat));
  NAND2_X1  g513(.A1(new_n683), .A2(new_n684), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n696), .A2(new_n715), .A3(new_n678), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G43gat), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT47), .ZN(new_n718));
  INV_X1    g517(.A(G43gat), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n700), .A2(new_n719), .A3(new_n452), .A4(new_n678), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n718), .B1(new_n717), .B2(new_n720), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(G1330gat));
  INV_X1    g522(.A(KEYINPUT48), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n424), .B(new_n678), .C1(new_n692), .C2(new_n693), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(G50gat), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n724), .B1(new_n726), .B2(KEYINPUT111), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n701), .A2(G50gat), .A3(new_n454), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n728), .B1(new_n725), .B2(G50gat), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n727), .B(new_n729), .ZN(G1331gat));
  NAND4_X1  g529(.A1(new_n552), .A2(new_n648), .A3(new_n595), .A4(new_n677), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n731), .B1(new_n691), .B2(new_n458), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n653), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n445), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n735), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT49), .B(G64gat), .Z(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(new_n735), .B2(new_n737), .ZN(G1333gat));
  NAND3_X1  g537(.A1(new_n732), .A2(new_n555), .A3(new_n452), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n732), .A2(new_n715), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n740), .B2(new_n555), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g541(.A1(new_n732), .A2(new_n424), .ZN(new_n743));
  XNOR2_X1  g542(.A(KEYINPUT112), .B(G78gat), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1335gat));
  NOR2_X1   g544(.A1(new_n692), .A2(new_n693), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n595), .A2(new_n647), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n624), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n653), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n490), .B2(new_n489), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n691), .A2(new_n458), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n552), .A2(new_n748), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n754), .A2(KEYINPUT51), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT51), .B1(new_n754), .B2(new_n755), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n677), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n653), .A2(new_n495), .A3(new_n497), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n753), .B1(new_n758), .B2(new_n759), .ZN(G1336gat));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(KEYINPUT52), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n624), .A2(new_n444), .A3(G92gat), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT113), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n756), .B2(new_n757), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n445), .B(new_n749), .C1(new_n692), .C2(new_n693), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(G92gat), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n762), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n761), .A2(KEYINPUT52), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(G1337gat));
  NAND2_X1  g569(.A1(new_n751), .A2(new_n715), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT115), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G99gat), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n771), .A2(KEYINPUT115), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n452), .A2(new_n499), .ZN(new_n775));
  OAI22_X1  g574(.A1(new_n773), .A2(new_n774), .B1(new_n758), .B2(new_n775), .ZN(G1338gat));
  NAND3_X1  g575(.A1(new_n696), .A2(new_n424), .A3(new_n749), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G106gat), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n454), .A2(G106gat), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n677), .B(new_n779), .C1(new_n756), .C2(new_n757), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT53), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n778), .A2(new_n783), .A3(new_n780), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(G1339gat));
  NOR2_X1   g584(.A1(new_n625), .A2(new_n647), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n609), .A2(new_n613), .A3(new_n602), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n617), .A2(new_n618), .ZN(new_n788));
  AOI22_X1  g587(.A1(new_n788), .A2(new_n603), .B1(new_n606), .B2(new_n608), .ZN(new_n789));
  OAI211_X1 g588(.A(KEYINPUT54), .B(new_n787), .C1(new_n789), .C2(new_n616), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n600), .B1(new_n614), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(new_n792), .A3(KEYINPUT55), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n790), .A2(new_n792), .A3(KEYINPUT116), .A4(KEYINPUT55), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n623), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n642), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n486), .A2(new_n584), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n627), .B1(new_n799), .B2(new_n626), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n634), .A2(new_n635), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n798), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n646), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n790), .A2(new_n792), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n547), .A2(new_n551), .A3(new_n797), .A4(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n624), .A2(new_n803), .ZN(new_n808));
  AOI22_X1  g607(.A1(new_n804), .A2(new_n805), .B1(new_n645), .B2(new_n646), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n808), .B1(new_n797), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n552), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI211_X1 g611(.A(KEYINPUT117), .B(new_n808), .C1(new_n797), .C2(new_n809), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n807), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n595), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n786), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n652), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n454), .A2(new_n295), .A3(new_n296), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n819), .A2(new_n445), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n648), .A2(new_n202), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n816), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n445), .A2(new_n652), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n823), .A2(new_n454), .A3(new_n452), .A4(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(G113gat), .B1(new_n825), .B2(new_n648), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n822), .A2(new_n826), .ZN(G1340gat));
  NOR3_X1   g626(.A1(new_n825), .A2(new_n205), .A3(new_n624), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n820), .A2(new_n677), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n829), .B2(new_n205), .ZN(G1341gat));
  INV_X1    g629(.A(G127gat), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n820), .A2(new_n831), .A3(new_n595), .ZN(new_n832));
  OAI21_X1  g631(.A(G127gat), .B1(new_n825), .B2(new_n815), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(G1342gat));
  INV_X1    g633(.A(G134gat), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n552), .A2(new_n445), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n817), .A2(new_n835), .A3(new_n818), .A4(new_n836), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n837), .A2(KEYINPUT56), .ZN(new_n838));
  OAI21_X1  g637(.A(G134gat), .B1(new_n825), .B2(new_n552), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(KEYINPUT56), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(G1343gat));
  INV_X1    g640(.A(KEYINPUT121), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n842), .A2(KEYINPUT58), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n683), .A2(new_n684), .A3(new_n824), .ZN(new_n845));
  XOR2_X1   g644(.A(new_n845), .B(KEYINPUT118), .Z(new_n846));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n847), .B(new_n848), .C1(new_n816), .C2(new_n454), .ZN(new_n849));
  INV_X1    g648(.A(new_n786), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n851));
  INV_X1    g650(.A(new_n803), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n677), .B2(new_n852), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n624), .A2(new_n803), .A3(KEYINPUT120), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n795), .A2(new_n796), .ZN(new_n856));
  INV_X1    g655(.A(new_n623), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n856), .A2(new_n857), .A3(new_n809), .ZN(new_n858));
  AOI22_X1  g657(.A1(new_n855), .A2(new_n858), .B1(new_n547), .B2(new_n551), .ZN(new_n859));
  INV_X1    g658(.A(new_n807), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n815), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n850), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(KEYINPUT57), .A3(new_n424), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n849), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n808), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n858), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT117), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n810), .A2(new_n811), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n552), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n595), .B1(new_n869), .B2(new_n807), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n424), .B1(new_n870), .B2(new_n786), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n847), .B1(new_n871), .B2(new_n848), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n647), .B(new_n846), .C1(new_n864), .C2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(G141gat), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n842), .A2(KEYINPUT58), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n715), .A2(new_n454), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n823), .A2(new_n876), .A3(new_n653), .A4(new_n444), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n648), .A2(G141gat), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n875), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n844), .B1(new_n874), .B2(new_n881), .ZN(new_n882));
  AOI211_X1 g681(.A(new_n843), .B(new_n880), .C1(new_n873), .C2(G141gat), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(G1344gat));
  AOI21_X1  g683(.A(new_n454), .B1(new_n850), .B2(new_n861), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n424), .A2(KEYINPUT57), .ZN(new_n886));
  OAI22_X1  g685(.A1(new_n885), .A2(KEYINPUT57), .B1(new_n816), .B2(new_n886), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n846), .A2(new_n677), .A3(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(G148gat), .ZN(new_n889));
  OAI21_X1  g688(.A(KEYINPUT59), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n889), .A2(KEYINPUT59), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n846), .B1(new_n864), .B2(new_n872), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(new_n624), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n877), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n889), .A3(new_n677), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(G1345gat));
  OAI21_X1  g696(.A(G155gat), .B1(new_n892), .B2(new_n815), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n895), .A2(new_n312), .A3(new_n595), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1346gat));
  OAI21_X1  g699(.A(G162gat), .B1(new_n892), .B2(new_n552), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n817), .A2(new_n876), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n836), .A2(new_n313), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(G1347gat));
  NOR2_X1   g703(.A1(new_n653), .A2(new_n444), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n818), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n816), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(G169gat), .B1(new_n907), .B2(new_n647), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n823), .A2(new_n454), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n452), .A2(new_n905), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n648), .A2(new_n219), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n908), .B1(new_n911), .B2(new_n912), .ZN(G1348gat));
  AOI21_X1  g712(.A(G176gat), .B1(new_n907), .B2(new_n677), .ZN(new_n914));
  XOR2_X1   g713(.A(new_n914), .B(KEYINPUT122), .Z(new_n915));
  OR2_X1    g714(.A1(new_n909), .A2(new_n910), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n916), .A2(new_n220), .A3(new_n624), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n915), .A2(new_n917), .ZN(G1349gat));
  NAND3_X1  g717(.A1(new_n907), .A2(new_n230), .A3(new_n595), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT123), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n235), .B1(new_n916), .B2(new_n815), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT60), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT60), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n920), .A2(new_n921), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1350gat));
  OAI211_X1 g725(.A(KEYINPUT124), .B(G190gat), .C1(new_n916), .C2(new_n552), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n909), .A2(new_n552), .A3(new_n910), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n929), .B2(new_n225), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n927), .A2(KEYINPUT61), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n907), .A2(new_n225), .A3(new_n679), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n931), .B(new_n932), .C1(KEYINPUT61), .C2(new_n930), .ZN(G1351gat));
  NAND2_X1  g732(.A1(new_n670), .A2(new_n905), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n871), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(G197gat), .B1(new_n935), .B2(new_n647), .ZN(new_n936));
  INV_X1    g735(.A(new_n934), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n887), .A2(new_n937), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n647), .A2(G197gat), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(G1352gat));
  XOR2_X1   g739(.A(KEYINPUT125), .B(G204gat), .Z(new_n941));
  NAND3_X1  g740(.A1(new_n935), .A2(new_n677), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n941), .B1(new_n938), .B2(new_n677), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n943), .B2(KEYINPUT62), .ZN(new_n944));
  OAI21_X1  g743(.A(KEYINPUT126), .B1(new_n942), .B2(KEYINPUT62), .ZN(new_n945));
  OR3_X1    g744(.A1(new_n942), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(G1353gat));
  NAND3_X1  g746(.A1(new_n935), .A2(new_n367), .A3(new_n595), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n887), .A2(KEYINPUT127), .A3(new_n595), .A4(new_n937), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n949), .A2(G211gat), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n887), .A2(new_n595), .A3(new_n937), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT63), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  AND4_X1   g753(.A1(KEYINPUT63), .A2(new_n953), .A3(G211gat), .A4(new_n949), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n948), .B1(new_n954), .B2(new_n955), .ZN(G1354gat));
  NAND3_X1  g755(.A1(new_n935), .A2(new_n368), .A3(new_n679), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n938), .A2(new_n679), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n957), .B1(new_n958), .B2(new_n368), .ZN(G1355gat));
endmodule


