//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT91), .Z(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G104), .ZN(new_n190));
  OR2_X1    g004(.A1(KEYINPUT84), .A2(G107), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT84), .A2(G107), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n190), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G104), .ZN(new_n194));
  OAI21_X1  g008(.A(G107), .B1(new_n194), .B2(KEYINPUT3), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(KEYINPUT3), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT85), .B1(new_n193), .B2(new_n197), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT84), .A2(G107), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT84), .A2(G107), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n189), .B(G104), .C1(new_n199), .C2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT85), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n201), .A2(new_n202), .A3(new_n196), .A4(new_n195), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n198), .A2(new_n203), .A3(G101), .ZN(new_n204));
  INV_X1    g018(.A(G101), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n201), .A2(new_n205), .A3(new_n196), .A4(new_n195), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT4), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT86), .B1(new_n204), .B2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n198), .A2(new_n203), .A3(G101), .ZN(new_n209));
  OR2_X1    g023(.A1(new_n209), .A2(KEYINPUT4), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT70), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT69), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n213));
  INV_X1    g027(.A(G113), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT69), .B1(KEYINPUT2), .B2(G113), .ZN(new_n216));
  AOI22_X1  g030(.A1(new_n215), .A2(new_n216), .B1(KEYINPUT2), .B2(G113), .ZN(new_n217));
  XNOR2_X1  g031(.A(G116), .B(G119), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n211), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n215), .A2(new_n216), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT2), .A2(G113), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n218), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(new_n211), .A3(new_n223), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT86), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n209), .A2(new_n228), .A3(KEYINPUT4), .A4(new_n206), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n208), .A2(new_n210), .A3(new_n227), .A4(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT5), .ZN(new_n231));
  INV_X1    g045(.A(G119), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n232), .A3(G116), .ZN(new_n233));
  XOR2_X1   g047(.A(new_n233), .B(KEYINPUT92), .Z(new_n234));
  OAI21_X1  g048(.A(G113), .B1(new_n223), .B2(new_n231), .ZN(new_n235));
  OAI22_X1  g049(.A1(new_n234), .A2(new_n235), .B1(new_n222), .B2(new_n223), .ZN(new_n236));
  NOR3_X1   g050(.A1(new_n199), .A2(new_n200), .A3(G104), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT87), .B1(new_n194), .B2(G107), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT87), .ZN(new_n239));
  INV_X1    g053(.A(G107), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n240), .A3(G104), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(G101), .B1(new_n237), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n206), .ZN(new_n244));
  OR2_X1    g058(.A1(new_n236), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n230), .A2(new_n245), .ZN(new_n246));
  XOR2_X1   g060(.A(G110), .B(G122), .Z(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n247), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n230), .A2(new_n245), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(KEYINPUT6), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G146), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(G143), .ZN(new_n253));
  INV_X1    g067(.A(G143), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT64), .B1(new_n254), .B2(G146), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT64), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(new_n252), .A3(G143), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n253), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n254), .A2(G146), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n252), .A2(G143), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OR2_X1    g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n258), .A2(new_n259), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G125), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n255), .A2(new_n257), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n266), .A2(new_n267), .A3(G128), .A4(new_n260), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n260), .A2(new_n261), .ZN(new_n269));
  INV_X1    g083(.A(G128), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT67), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT67), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G128), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n267), .B1(G143), .B2(new_n252), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n269), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n268), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n265), .B1(new_n277), .B2(G125), .ZN(new_n278));
  INV_X1    g092(.A(G953), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G224), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n280), .B(KEYINPUT93), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n278), .B(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n246), .A2(new_n283), .A3(new_n247), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n251), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G902), .ZN(new_n286));
  NAND2_X1  g100(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n278), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n281), .A2(KEYINPUT7), .ZN(new_n289));
  XOR2_X1   g103(.A(new_n288), .B(new_n289), .Z(new_n290));
  INV_X1    g104(.A(new_n244), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n236), .B(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n247), .B(KEYINPUT8), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n290), .B(new_n250), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n285), .A2(new_n286), .A3(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G210), .B1(G237), .B2(G902), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n296), .A2(KEYINPUT95), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n297), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n285), .A2(new_n286), .A3(new_n299), .A4(new_n294), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n188), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  XOR2_X1   g115(.A(KEYINPUT9), .B(G234), .Z(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(G221), .B1(new_n303), .B2(G902), .ZN(new_n304));
  XOR2_X1   g118(.A(new_n304), .B(KEYINPUT82), .Z(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(G110), .B(G140), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n279), .A2(G227), .ZN(new_n308));
  XOR2_X1   g122(.A(new_n307), .B(new_n308), .Z(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n208), .A2(new_n210), .A3(new_n264), .A4(new_n229), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT10), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n277), .A2(new_n244), .A3(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n275), .A2(new_n270), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n268), .B1(new_n258), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n291), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n313), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT11), .ZN(new_n318));
  INV_X1    g132(.A(G134), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n318), .B1(new_n319), .B2(G137), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(G137), .ZN(new_n321));
  INV_X1    g135(.A(G137), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(KEYINPUT11), .A3(G134), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n320), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G131), .ZN(new_n325));
  INV_X1    g139(.A(G131), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n320), .A2(new_n323), .A3(new_n326), .A4(new_n321), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n311), .A2(new_n317), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n328), .B1(new_n311), .B2(new_n317), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n310), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n311), .A2(new_n317), .A3(new_n328), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n277), .A2(new_n244), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT88), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n328), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT12), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT89), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n337), .B1(new_n328), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n316), .A2(new_n333), .A3(KEYINPUT88), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n336), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n339), .B1(new_n336), .B2(new_n340), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n332), .B(new_n309), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(G902), .B1(new_n331), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n306), .B1(new_n344), .B2(G469), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT90), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(new_n329), .B2(new_n310), .ZN(new_n347));
  INV_X1    g161(.A(new_n330), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n332), .A2(KEYINPUT90), .A3(new_n309), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n332), .B1(new_n341), .B2(new_n342), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n309), .B(KEYINPUT83), .Z(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(G902), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n345), .B1(G469), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G234), .ZN(new_n356));
  OAI21_X1  g170(.A(G217), .B1(new_n356), .B2(G902), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(KEYINPUT76), .ZN(new_n358));
  INV_X1    g172(.A(G140), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G125), .ZN(new_n360));
  INV_X1    g174(.A(G125), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G140), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n360), .A2(new_n362), .A3(KEYINPUT78), .A4(KEYINPUT16), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n360), .A2(new_n362), .A3(KEYINPUT16), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT78), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n365), .B1(new_n360), .B2(KEYINPUT16), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n363), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G146), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n252), .B(new_n363), .C1(new_n364), .C2(new_n366), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n270), .A2(G119), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n370), .B1(new_n274), .B2(G119), .ZN(new_n371));
  XOR2_X1   g185(.A(KEYINPUT24), .B(G110), .Z(new_n372));
  AOI22_X1  g186(.A1(new_n368), .A2(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G110), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n274), .A2(KEYINPUT23), .A3(G119), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT77), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT23), .B1(new_n270), .B2(G119), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(new_n370), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n274), .A2(KEYINPUT77), .A3(KEYINPUT23), .A4(G119), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n377), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n373), .B1(new_n374), .B2(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n377), .A2(new_n380), .A3(new_n374), .A4(new_n379), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n383), .B1(new_n371), .B2(new_n372), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n360), .A2(new_n362), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(KEYINPUT79), .A3(new_n252), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT79), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n360), .A2(new_n362), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n387), .B1(new_n388), .B2(G146), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n368), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n384), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT22), .B(G137), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(KEYINPUT80), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n279), .A2(G221), .A3(G234), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n394), .B(new_n396), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n382), .A2(new_n392), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n397), .B1(new_n382), .B2(new_n392), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT25), .B1(new_n400), .B2(new_n286), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n382), .A2(new_n392), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n394), .B(new_n395), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n382), .A2(new_n392), .A3(new_n397), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n404), .A2(KEYINPUT25), .A3(new_n286), .A4(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n358), .B1(new_n401), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT81), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n404), .A2(new_n286), .A3(new_n405), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(new_n358), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n408), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n358), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT25), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n414), .B1(new_n416), .B2(new_n406), .ZN(new_n417));
  OAI21_X1  g231(.A(KEYINPUT81), .B1(new_n417), .B2(new_n411), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n301), .A2(new_n355), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT28), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n256), .B1(G143), .B2(new_n252), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n254), .A2(KEYINPUT64), .A3(G146), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n260), .B(new_n259), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n259), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n269), .A2(new_n425), .A3(new_n263), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n424), .A2(KEYINPUT65), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT65), .B1(new_n424), .B2(new_n426), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n427), .A2(new_n328), .A3(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n322), .A2(G134), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n319), .A2(G137), .ZN(new_n431));
  OAI21_X1  g245(.A(G131), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n327), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT66), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n268), .A2(new_n276), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n327), .A2(new_n432), .A3(KEYINPUT66), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n227), .B1(new_n429), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n325), .A2(new_n327), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n264), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT71), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n225), .A2(new_n226), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT71), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n440), .A2(new_n264), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n436), .A2(new_n327), .A3(new_n432), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n442), .A2(new_n443), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n421), .B1(new_n439), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n443), .A2(new_n441), .A3(new_n446), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n421), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(G101), .ZN(new_n454));
  INV_X1    g268(.A(G237), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n455), .A2(new_n279), .A3(G210), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n454), .B(new_n456), .Z(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT30), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n429), .B2(new_n438), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT68), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n442), .A2(KEYINPUT30), .A3(new_n445), .A4(new_n446), .ZN(new_n464));
  OAI211_X1 g278(.A(KEYINPUT68), .B(new_n460), .C1(new_n429), .C2(new_n438), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n463), .A2(new_n227), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n447), .A2(new_n457), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT72), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n447), .A2(KEYINPUT72), .A3(new_n457), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n466), .A2(new_n471), .A3(KEYINPUT31), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT31), .B1(new_n466), .B2(new_n471), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n459), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(G472), .A2(G902), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT73), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT32), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT32), .ZN(new_n479));
  AOI211_X1 g293(.A(KEYINPUT73), .B(new_n479), .C1(new_n474), .C2(new_n475), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n466), .A2(new_n447), .ZN(new_n481));
  AOI21_X1  g295(.A(KEYINPUT29), .B1(new_n481), .B2(new_n458), .ZN(new_n482));
  INV_X1    g296(.A(new_n451), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n448), .A2(new_n483), .A3(new_n458), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT74), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n457), .B1(new_n466), .B2(new_n447), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT74), .ZN(new_n488));
  NOR4_X1   g302(.A1(new_n487), .A2(new_n484), .A3(new_n488), .A4(KEYINPUT29), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n442), .A2(new_n445), .A3(new_n446), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n227), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n447), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT28), .ZN(new_n493));
  OR2_X1    g307(.A1(new_n451), .A2(KEYINPUT75), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n451), .A2(KEYINPUT75), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n457), .A2(KEYINPUT29), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n286), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n486), .A2(new_n489), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G472), .ZN(new_n501));
  OAI22_X1  g315(.A1(new_n478), .A2(new_n480), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(G475), .ZN(new_n503));
  INV_X1    g317(.A(G122), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n214), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(G113), .A2(G122), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT98), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT98), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n505), .A2(new_n509), .A3(new_n506), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(G104), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(G104), .B1(new_n508), .B2(new_n510), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT99), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT99), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n508), .A2(new_n510), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n194), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n515), .B1(new_n517), .B2(new_n511), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n455), .A2(new_n279), .A3(G214), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n254), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n455), .A2(new_n279), .A3(G143), .A4(G214), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT96), .ZN(new_n524));
  NAND2_X1  g338(.A1(KEYINPUT18), .A2(G131), .ZN(new_n525));
  OR3_X1    g339(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n525), .B1(new_n523), .B2(new_n524), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n390), .B1(new_n252), .B2(new_n385), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n523), .A2(G131), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n521), .A2(new_n326), .A3(new_n522), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n523), .A2(KEYINPUT17), .A3(G131), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n534), .A2(new_n368), .A3(new_n369), .A4(new_n535), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n519), .A2(new_n530), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n517), .A2(new_n511), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n531), .A2(new_n533), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT19), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n385), .B1(KEYINPUT97), .B2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n541), .B1(new_n385), .B2(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n368), .B(new_n539), .C1(new_n543), .C2(G146), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n538), .B1(new_n530), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n503), .B(new_n286), .C1(new_n537), .C2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT20), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n545), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n519), .A2(new_n530), .A3(new_n536), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n551), .A2(KEYINPUT20), .A3(new_n503), .A4(new_n286), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n538), .B1(new_n530), .B2(new_n536), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n286), .B1(new_n537), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(G475), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n548), .A2(new_n552), .A3(new_n555), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n504), .A2(G116), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n504), .A2(KEYINPUT100), .A3(G116), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT100), .B1(new_n504), .B2(G116), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n199), .A2(new_n200), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n254), .B1(new_n271), .B2(new_n273), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n270), .A2(G143), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT101), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT101), .ZN(new_n566));
  INV_X1    g380(.A(new_n564), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT67), .B(G128), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n566), .B(new_n567), .C1(new_n568), .C2(new_n254), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n565), .A2(new_n319), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n563), .B1(KEYINPUT13), .B2(new_n564), .ZN(new_n571));
  OR2_X1    g385(.A1(new_n564), .A2(KEYINPUT13), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n562), .B(new_n570), .C1(new_n573), .C2(new_n319), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n560), .A2(new_n561), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n557), .B(KEYINPUT14), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n558), .A2(new_n559), .ZN(new_n577));
  OAI21_X1  g391(.A(G107), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n565), .A2(new_n319), .A3(new_n569), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n319), .B1(new_n565), .B2(new_n569), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n575), .B(new_n578), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n302), .A2(G217), .A3(new_n279), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n574), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n583), .B1(new_n574), .B2(new_n581), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n286), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G478), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(KEYINPUT15), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n588), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n286), .B(new_n590), .C1(new_n584), .C2(new_n585), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(G234), .A2(G237), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(G952), .A3(new_n279), .ZN(new_n595));
  XOR2_X1   g409(.A(KEYINPUT21), .B(G898), .Z(new_n596));
  NAND3_X1  g410(.A1(new_n594), .A2(G902), .A3(G953), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(KEYINPUT102), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n556), .A2(new_n593), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(KEYINPUT103), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n420), .A2(new_n502), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  NAND2_X1  g417(.A1(new_n295), .A2(new_n296), .ZN(new_n604));
  INV_X1    g418(.A(new_n188), .ZN(new_n605));
  INV_X1    g419(.A(new_n296), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n285), .A2(new_n286), .A3(new_n606), .A4(new_n294), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n604), .A2(new_n599), .A3(new_n605), .A4(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n548), .A2(new_n552), .A3(new_n555), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT104), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(KEYINPUT104), .A2(KEYINPUT33), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n612), .B(new_n613), .C1(new_n584), .C2(new_n585), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n574), .A2(new_n581), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n582), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n574), .A2(new_n581), .A3(new_n583), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n616), .A2(new_n610), .A3(new_n611), .A4(new_n617), .ZN(new_n618));
  AOI211_X1 g432(.A(new_n587), .B(G902), .C1(new_n614), .C2(new_n618), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n586), .A2(new_n587), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n609), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n608), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n413), .A2(new_n418), .ZN(new_n623));
  INV_X1    g437(.A(new_n476), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n501), .B1(new_n474), .B2(new_n286), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n622), .A2(new_n626), .A3(new_n355), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT34), .B(G104), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G6));
  NAND2_X1  g443(.A1(new_n556), .A2(new_n592), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n608), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n631), .A2(new_n626), .A3(new_n355), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  OAI21_X1  g448(.A(KEYINPUT105), .B1(new_n403), .B2(KEYINPUT36), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT105), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT36), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n397), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n402), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n635), .A2(new_n638), .A3(new_n382), .A4(new_n392), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n640), .A2(new_n286), .A3(new_n414), .A4(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT106), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n417), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n624), .A2(new_n625), .A3(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n601), .A2(new_n646), .A3(new_n301), .A4(new_n355), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT107), .B(KEYINPUT37), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(new_n374), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n647), .B(new_n649), .ZN(G12));
  NAND2_X1  g464(.A1(new_n354), .A2(G469), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n331), .A2(new_n343), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n286), .ZN(new_n653));
  INV_X1    g467(.A(G469), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n305), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(new_n645), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n595), .B(KEYINPUT108), .ZN(new_n658));
  INV_X1    g472(.A(G900), .ZN(new_n659));
  INV_X1    g473(.A(new_n597), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n593), .A2(new_n609), .A3(new_n661), .ZN(new_n662));
  AND4_X1   g476(.A1(new_n605), .A2(new_n662), .A3(new_n604), .A4(new_n607), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n502), .A2(new_n657), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G128), .ZN(G30));
  NAND2_X1  g479(.A1(new_n476), .A2(new_n477), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n479), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT32), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI22_X1  g483(.A1(new_n466), .A2(new_n471), .B1(new_n458), .B2(new_n492), .ZN(new_n670));
  OAI21_X1  g484(.A(G472), .B1(new_n670), .B2(G902), .ZN(new_n671));
  AOI21_X1  g485(.A(KEYINPUT109), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  OAI211_X1 g486(.A(KEYINPUT109), .B(new_n671), .C1(new_n478), .C2(new_n480), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n661), .B(KEYINPUT39), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n355), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n675), .B1(KEYINPUT40), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n609), .A2(new_n592), .ZN(new_n680));
  INV_X1    g494(.A(new_n678), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT40), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n298), .A2(new_n300), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT38), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n642), .B(KEYINPUT106), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n408), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n679), .A2(new_n605), .A3(new_n683), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G143), .ZN(G45));
  NAND3_X1  g505(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n692));
  AOI21_X1  g506(.A(G902), .B1(new_n614), .B2(new_n618), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n620), .B1(new_n693), .B2(G478), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n694), .A2(new_n556), .A3(new_n661), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(KEYINPUT110), .B1(new_n692), .B2(new_n696), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n604), .A2(new_n607), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n698), .A2(new_n699), .A3(new_n605), .A4(new_n695), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n502), .A2(new_n697), .A3(new_n700), .A4(new_n657), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  NOR2_X1   g516(.A1(new_n653), .A2(new_n654), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n344), .A2(G469), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n305), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n502), .A2(new_n622), .A3(new_n419), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NAND4_X1  g523(.A1(new_n502), .A2(new_n419), .A3(new_n631), .A4(new_n706), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT111), .B(G116), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G18));
  OAI211_X1 g526(.A(new_n688), .B(new_n306), .C1(new_n703), .C2(new_n704), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n692), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n502), .A2(new_n714), .A3(new_n601), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G119), .ZN(G21));
  NOR2_X1   g530(.A1(new_n692), .A2(new_n680), .ZN(new_n717));
  XOR2_X1   g531(.A(KEYINPUT112), .B(G472), .Z(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n474), .B2(new_n286), .ZN(new_n720));
  INV_X1    g534(.A(new_n475), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n466), .A2(new_n471), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT31), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n466), .A2(new_n471), .A3(KEYINPUT31), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n496), .A2(new_n458), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n721), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n408), .A2(new_n412), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n720), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n717), .A2(new_n706), .A3(new_n599), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(KEYINPUT113), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(new_n504), .ZN(G24));
  NOR2_X1   g547(.A1(new_n720), .A2(new_n728), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n714), .A2(new_n695), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  INV_X1    g550(.A(new_n486), .ZN(new_n737));
  INV_X1    g551(.A(new_n499), .ZN(new_n738));
  INV_X1    g552(.A(new_n489), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(G472), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n476), .B(KEYINPUT32), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n729), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n298), .A2(new_n605), .A3(new_n300), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n696), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n743), .A2(KEYINPUT42), .A3(new_n355), .A4(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n656), .A2(new_n744), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n502), .A2(new_n419), .A3(new_n695), .A4(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G131), .ZN(G33));
  NAND4_X1  g566(.A1(new_n502), .A2(new_n419), .A3(new_n662), .A4(new_n747), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G134), .ZN(G36));
  INV_X1    g568(.A(new_n694), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n556), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(KEYINPUT43), .Z(new_n757));
  OAI211_X1 g571(.A(new_n757), .B(new_n688), .C1(new_n624), .C2(new_n625), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n744), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n350), .A2(new_n353), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT45), .ZN(new_n765));
  OAI21_X1  g579(.A(G469), .B1(new_n765), .B2(G902), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT46), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT46), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n768), .B(G469), .C1(new_n765), .C2(G902), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n767), .B(new_n769), .C1(G469), .C2(new_n653), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n306), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n763), .B1(new_n771), .B2(new_n676), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n770), .A2(KEYINPUT114), .A3(new_n306), .A4(new_n677), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n762), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n758), .A2(new_n759), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(KEYINPUT115), .Z(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G137), .ZN(G39));
  INV_X1    g592(.A(KEYINPUT47), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT116), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n771), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n502), .A2(new_n419), .ZN(new_n782));
  XOR2_X1   g596(.A(KEYINPUT116), .B(KEYINPUT47), .Z(new_n783));
  NAND3_X1  g597(.A1(new_n770), .A2(new_n306), .A3(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n781), .A2(new_n745), .A3(new_n782), .A4(new_n784), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n785), .A2(KEYINPUT117), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(KEYINPUT117), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G140), .ZN(G42));
  NAND4_X1  g603(.A1(new_n707), .A2(new_n710), .A3(new_n715), .A4(new_n731), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(KEYINPUT122), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n790), .A2(KEYINPUT122), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n751), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT123), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT123), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n795), .B(new_n751), .C1(new_n791), .C2(new_n792), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n797));
  INV_X1    g611(.A(new_n717), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n799));
  INV_X1    g613(.A(new_n661), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n799), .B1(new_n645), .B2(new_n800), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n688), .A2(KEYINPUT120), .A3(new_n661), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n355), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n671), .B1(new_n478), .B2(new_n480), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT109), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI211_X1 g620(.A(new_n798), .B(new_n803), .C1(new_n806), .C2(new_n673), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n701), .A2(new_n664), .A3(new_n735), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n797), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n803), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n717), .B(new_n810), .C1(new_n672), .C2(new_n674), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n664), .A2(new_n735), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n811), .A2(new_n812), .A3(KEYINPUT52), .A4(new_n701), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n599), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n592), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n589), .A2(KEYINPUT119), .A3(new_n591), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI22_X1  g633(.A1(new_n621), .A2(KEYINPUT118), .B1(new_n819), .B2(new_n556), .ZN(new_n820));
  OR3_X1    g634(.A1(new_n694), .A2(new_n556), .A3(KEYINPUT118), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n815), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n822), .A2(new_n626), .A3(new_n301), .A4(new_n355), .ZN(new_n823));
  AND4_X1   g637(.A1(new_n602), .A2(new_n753), .A3(new_n647), .A4(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n609), .A2(new_n661), .ZN(new_n825));
  INV_X1    g639(.A(new_n819), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n502), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n734), .A2(new_n695), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n657), .A3(new_n761), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n824), .A2(KEYINPUT53), .A3(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n794), .A2(new_n796), .A3(new_n814), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n833));
  AND4_X1   g647(.A1(new_n707), .A2(new_n710), .A3(new_n715), .A4(new_n731), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n751), .A2(new_n834), .A3(new_n824), .A4(new_n830), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n814), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT121), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n839));
  AOI211_X1 g653(.A(new_n839), .B(KEYINPUT53), .C1(new_n835), .C2(new_n814), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n832), .B(new_n833), .C1(new_n838), .C2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n834), .A2(new_n824), .A3(new_n751), .A4(new_n830), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n842), .B1(new_n809), .B2(new_n813), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n814), .A2(new_n831), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n834), .A2(new_n751), .ZN(new_n845));
  OAI22_X1  g659(.A1(new_n843), .A2(KEYINPUT53), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT54), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n841), .A2(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n757), .A2(new_n658), .A3(new_n730), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n706), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n848), .B1(new_n692), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n623), .A2(new_n595), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n675), .A2(new_n706), .A3(new_n761), .A4(new_n852), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n853), .A2(new_n621), .ZN(new_n854));
  AND4_X1   g668(.A1(new_n658), .A2(new_n757), .A3(new_n706), .A4(new_n761), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n743), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT48), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n857), .A2(G952), .A3(new_n279), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n781), .A2(new_n784), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n705), .A2(new_n306), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n761), .B(new_n849), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n853), .A2(new_n609), .A3(new_n755), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n720), .A2(new_n645), .A3(new_n728), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n862), .B1(new_n855), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n686), .A2(new_n188), .ZN(new_n865));
  OR3_X1    g679(.A1(new_n850), .A2(KEYINPUT50), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT50), .B1(new_n850), .B2(new_n865), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n861), .A2(new_n864), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT124), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n868), .A2(new_n869), .A3(KEYINPUT51), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT51), .B1(new_n868), .B2(new_n869), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n854), .B(new_n858), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  OAI22_X1  g686(.A1(new_n851), .A2(new_n872), .B1(G952), .B2(G953), .ZN(new_n873));
  AOI211_X1 g687(.A(new_n756), .B(new_n685), .C1(KEYINPUT49), .C2(new_n705), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n874), .B(new_n675), .C1(KEYINPUT49), .C2(new_n705), .ZN(new_n875));
  OR4_X1    g689(.A1(new_n188), .A2(new_n875), .A3(new_n305), .A4(new_n729), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n873), .A2(new_n876), .ZN(G75));
  OAI21_X1  g691(.A(new_n839), .B1(new_n843), .B2(KEYINPUT53), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n836), .A2(KEYINPUT121), .A3(new_n837), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n286), .B1(new_n880), .B2(new_n832), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT56), .B1(new_n881), .B2(G210), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n251), .A2(new_n284), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(new_n282), .Z(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT55), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  AOI211_X1 g701(.A(KEYINPUT56), .B(new_n885), .C1(new_n881), .C2(G210), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n279), .A2(G952), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(G51));
  OAI21_X1  g704(.A(KEYINPUT57), .B1(new_n654), .B2(new_n286), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n833), .B1(new_n880), .B2(new_n832), .ZN(new_n892));
  INV_X1    g706(.A(new_n841), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n654), .A2(new_n286), .A3(KEYINPUT57), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n652), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n881), .A2(G469), .A3(new_n765), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n889), .B1(new_n896), .B2(new_n897), .ZN(G54));
  NAND3_X1  g712(.A1(new_n881), .A2(KEYINPUT58), .A3(G475), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(new_n550), .A3(new_n549), .ZN(new_n900));
  INV_X1    g714(.A(new_n889), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n881), .A2(KEYINPUT58), .A3(G475), .A4(new_n551), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(G60));
  NAND2_X1  g717(.A1(new_n614), .A2(new_n618), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(G478), .A2(G902), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT59), .Z(new_n907));
  NOR2_X1   g721(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n908), .B1(new_n892), .B2(new_n893), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n909), .A2(new_n910), .A3(new_n901), .ZN(new_n911));
  INV_X1    g725(.A(new_n908), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n832), .B1(new_n838), .B2(new_n840), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT54), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n912), .B1(new_n914), .B2(new_n841), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT125), .B1(new_n915), .B2(new_n889), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n905), .B1(new_n848), .B2(new_n907), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n911), .A2(new_n916), .A3(new_n917), .ZN(G63));
  NAND2_X1  g732(.A1(G217), .A2(G902), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT60), .Z(new_n920));
  NAND2_X1  g734(.A1(new_n913), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n400), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n889), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n640), .A2(new_n641), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(new_n921), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n923), .B(KEYINPUT61), .C1(new_n924), .C2(new_n921), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(G66));
  AOI21_X1  g743(.A(new_n279), .B1(new_n596), .B2(G224), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n834), .A2(new_n602), .A3(new_n647), .A4(new_n823), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n930), .B1(new_n931), .B2(new_n279), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n883), .B1(G898), .B2(new_n279), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n932), .B(new_n933), .Z(G69));
  AOI21_X1  g748(.A(new_n279), .B1(G227), .B2(G900), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT127), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n808), .B1(new_n786), .B2(new_n787), .ZN(new_n937));
  INV_X1    g751(.A(new_n751), .ZN(new_n938));
  INV_X1    g752(.A(new_n753), .ZN(new_n939));
  AOI211_X1 g753(.A(new_n938), .B(new_n939), .C1(new_n774), .C2(new_n776), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n772), .A2(new_n773), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n941), .A2(new_n717), .A3(new_n743), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n937), .A2(new_n940), .A3(new_n279), .A4(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(new_n543), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(G900), .B2(G953), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n936), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n808), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n690), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n690), .A2(KEYINPUT62), .A3(new_n951), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n820), .A2(new_n821), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n502), .A2(new_n419), .A3(new_n957), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n958), .A2(new_n678), .A3(new_n744), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n774), .B2(new_n776), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n788), .A2(new_n956), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n279), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n946), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n948), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n950), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n963), .B(new_n948), .C1(new_n949), .C2(new_n936), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(G72));
  NAND2_X1  g781(.A1(G472), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT63), .Z(new_n969));
  NAND3_X1  g783(.A1(new_n937), .A2(new_n940), .A3(new_n942), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n969), .B1(new_n970), .B2(new_n931), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n971), .A2(new_n447), .A3(new_n458), .A4(new_n466), .ZN(new_n972));
  INV_X1    g786(.A(new_n969), .ZN(new_n973));
  INV_X1    g787(.A(new_n487), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n973), .B1(new_n974), .B2(new_n722), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n889), .B1(new_n846), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n969), .B1(new_n961), .B2(new_n931), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n977), .A2(new_n457), .A3(new_n481), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n972), .A2(new_n976), .A3(new_n978), .ZN(G57));
endmodule


