//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G143), .B(G146), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT0), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  XOR2_X1   g005(.A(KEYINPUT0), .B(G128), .Z(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n188), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G131), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G137), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT11), .A2(G134), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT65), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n198));
  INV_X1    g012(.A(new_n196), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(G137), .ZN(new_n201));
  INV_X1    g015(.A(G137), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(KEYINPUT64), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n198), .B(new_n199), .C1(new_n201), .C2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n197), .A2(new_n204), .ZN(new_n205));
  OR2_X1    g019(.A1(KEYINPUT11), .A2(G134), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n199), .B1(new_n206), .B2(new_n202), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n194), .B1(new_n205), .B2(new_n208), .ZN(new_n209));
  AOI211_X1 g023(.A(G131), .B(new_n207), .C1(new_n197), .C2(new_n204), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n193), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT68), .ZN(new_n212));
  INV_X1    g026(.A(G119), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(G116), .ZN(new_n214));
  INV_X1    g028(.A(G116), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT68), .A3(G119), .ZN(new_n216));
  AOI22_X1  g030(.A1(new_n214), .A2(new_n216), .B1(G116), .B2(new_n213), .ZN(new_n217));
  NOR2_X1   g031(.A1(KEYINPUT2), .A2(G113), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT2), .A2(G113), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT67), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(KEYINPUT2), .A3(G113), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n218), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n217), .A2(KEYINPUT69), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(KEYINPUT69), .B1(new_n217), .B2(new_n223), .ZN(new_n225));
  OAI22_X1  g039(.A1(new_n224), .A2(new_n225), .B1(new_n223), .B2(new_n217), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n205), .A2(new_n194), .A3(new_n208), .ZN(new_n228));
  NAND2_X1  g042(.A1(G134), .A2(G137), .ZN(new_n229));
  OAI211_X1 g043(.A(G131), .B(new_n229), .C1(new_n195), .C2(G134), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT1), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n188), .A2(new_n231), .A3(G128), .ZN(new_n232));
  INV_X1    g046(.A(G146), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G143), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT1), .ZN(new_n235));
  INV_X1    g049(.A(G143), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(G146), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n190), .B1(new_n237), .B2(new_n234), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n232), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n228), .A2(new_n230), .A3(new_n239), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n211), .A2(new_n227), .A3(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(KEYINPUT28), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n211), .A2(KEYINPUT66), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n245), .B(new_n193), .C1(new_n209), .C2(new_n210), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n244), .A2(new_n240), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n241), .B1(new_n247), .B2(new_n226), .ZN(new_n248));
  XOR2_X1   g062(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n249));
  OAI21_X1  g063(.A(new_n243), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(G237), .A2(G953), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G210), .ZN(new_n252));
  XOR2_X1   g066(.A(new_n252), .B(G101), .Z(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n254));
  XOR2_X1   g068(.A(new_n253), .B(new_n254), .Z(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n250), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT30), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n247), .A2(new_n258), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n211), .A2(KEYINPUT30), .A3(new_n240), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n259), .A2(new_n226), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT31), .ZN(new_n263));
  INV_X1    g077(.A(new_n241), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n262), .A2(new_n263), .A3(new_n255), .A4(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n257), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n260), .B1(new_n247), .B2(new_n258), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n241), .B1(new_n267), .B2(new_n226), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n263), .B1(new_n268), .B2(new_n255), .ZN(new_n269));
  OAI211_X1 g083(.A(KEYINPUT32), .B(new_n187), .C1(new_n266), .C2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n187), .B1(new_n266), .B2(new_n269), .ZN(new_n271));
  XOR2_X1   g085(.A(KEYINPUT71), .B(KEYINPUT32), .Z(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n243), .B(new_n255), .C1(new_n248), .C2(new_n249), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT29), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n276), .B(new_n277), .C1(new_n268), .C2(new_n255), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n227), .B1(new_n211), .B2(new_n240), .ZN(new_n279));
  OR2_X1    g093(.A1(new_n241), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n242), .B1(new_n280), .B2(KEYINPUT28), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n256), .A2(new_n277), .ZN(new_n282));
  AOI21_X1  g096(.A(G902), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n275), .B1(new_n284), .B2(G472), .ZN(new_n285));
  INV_X1    g099(.A(G472), .ZN(new_n286));
  AOI211_X1 g100(.A(KEYINPUT72), .B(new_n286), .C1(new_n278), .C2(new_n283), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n270), .B(new_n274), .C1(new_n285), .C2(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(KEYINPUT74), .B(G125), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n191), .B(new_n289), .C1(new_n188), .C2(new_n192), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n290), .B1(new_n239), .B2(new_n289), .ZN(new_n291));
  INV_X1    g105(.A(G224), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n292), .A2(G953), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n293), .B(KEYINPUT85), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n291), .B(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n217), .A2(new_n223), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT69), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n217), .A2(new_n223), .A3(KEYINPUT69), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G104), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G107), .ZN(new_n302));
  INV_X1    g116(.A(G107), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G104), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G101), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT3), .B1(new_n301), .B2(G107), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT3), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(new_n303), .A3(G104), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n307), .A2(new_n309), .A3(new_n302), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT79), .B(G101), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n306), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n213), .A2(G116), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n215), .A2(KEYINPUT68), .A3(G119), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT68), .B1(new_n215), .B2(G119), .ZN(new_n316));
  OAI211_X1 g130(.A(KEYINPUT5), .B(new_n314), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  OR2_X1    g131(.A1(new_n314), .A2(KEYINPUT5), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(G113), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT82), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT82), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n317), .A2(new_n321), .A3(G113), .A4(new_n318), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n300), .A2(new_n313), .A3(new_n320), .A4(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT4), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n310), .A2(new_n324), .A3(G101), .ZN(new_n325));
  AND3_X1   g139(.A1(new_n307), .A2(new_n309), .A3(new_n302), .ZN(new_n326));
  INV_X1    g140(.A(new_n311), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n310), .A2(G101), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n226), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n323), .A2(new_n331), .ZN(new_n332));
  XOR2_X1   g146(.A(G110), .B(G122), .Z(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n333), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n323), .A2(new_n331), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(KEYINPUT6), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT83), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT6), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  AOI211_X1 g154(.A(new_n335), .B(new_n340), .C1(new_n323), .C2(new_n331), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n338), .A2(KEYINPUT6), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT84), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n332), .A2(new_n343), .A3(new_n333), .A4(new_n339), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT84), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n295), .B(new_n337), .C1(new_n344), .C2(new_n347), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n300), .A2(new_n312), .A3(new_n320), .A4(new_n322), .ZN(new_n349));
  XOR2_X1   g163(.A(new_n333), .B(KEYINPUT8), .Z(new_n350));
  AND2_X1   g164(.A1(new_n300), .A2(new_n319), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n349), .B(new_n350), .C1(new_n351), .C2(new_n312), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n352), .A2(new_n336), .ZN(new_n353));
  INV_X1    g167(.A(new_n290), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT7), .ZN(new_n355));
  OAI22_X1  g169(.A1(new_n354), .A2(KEYINPUT86), .B1(new_n355), .B2(new_n293), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(new_n291), .ZN(new_n357));
  AOI21_X1  g171(.A(G902), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n348), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(G210), .B1(G237), .B2(G902), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT87), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n348), .A2(new_n360), .A3(new_n358), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(G214), .B1(G237), .B2(G902), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n348), .A2(KEYINPUT87), .A3(new_n360), .A4(new_n358), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT16), .ZN(new_n369));
  INV_X1    g183(.A(G140), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n289), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(G125), .A2(G140), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n372), .B1(new_n289), .B2(G140), .ZN(new_n373));
  OAI211_X1 g187(.A(G146), .B(new_n371), .C1(new_n373), .C2(new_n369), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n251), .A2(G143), .A3(G214), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(G143), .B1(new_n251), .B2(G214), .ZN(new_n377));
  OAI21_X1  g191(.A(G131), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n377), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n194), .A3(new_n375), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n373), .A2(KEYINPUT19), .ZN(new_n382));
  XNOR2_X1  g196(.A(G125), .B(G140), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT19), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n374), .B(new_n381), .C1(new_n386), .C2(G146), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(new_n233), .ZN(new_n388));
  INV_X1    g202(.A(new_n373), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n388), .B1(new_n389), .B2(new_n233), .ZN(new_n390));
  NAND2_X1  g204(.A1(KEYINPUT18), .A2(G131), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n379), .A2(new_n375), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n379), .A2(new_n375), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(KEYINPUT18), .A3(G131), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n390), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n387), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(G113), .B(G122), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(new_n301), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n398), .B(KEYINPUT89), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n371), .B1(new_n373), .B2(new_n369), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n233), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n374), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n393), .A2(KEYINPUT17), .A3(G131), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n381), .B2(KEYINPUT17), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n401), .B(new_n395), .C1(new_n404), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n400), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(G475), .A2(G902), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n409), .B(KEYINPUT91), .Z(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(KEYINPUT20), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n408), .A2(KEYINPUT90), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT90), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n400), .A2(new_n414), .A3(new_n407), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n410), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n412), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n407), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n395), .B1(new_n404), .B2(new_n406), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT92), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n398), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n395), .B(KEYINPUT92), .C1(new_n404), .C2(new_n406), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n420), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(G475), .B1(new_n425), .B2(G902), .ZN(new_n426));
  NAND2_X1  g240(.A1(G234), .A2(G237), .ZN(new_n427));
  INV_X1    g241(.A(G953), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(G952), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  XOR2_X1   g244(.A(KEYINPUT21), .B(G898), .Z(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n427), .A2(G902), .A3(G953), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n430), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n419), .A2(new_n426), .A3(new_n436), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n232), .A2(new_n235), .A3(new_n238), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT80), .B1(new_n438), .B2(new_n312), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT80), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n313), .A2(new_n440), .A3(new_n239), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT10), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n439), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n313), .A2(KEYINPUT10), .A3(new_n239), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n330), .A2(new_n193), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n209), .A2(new_n210), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n443), .A2(new_n447), .A3(new_n444), .A4(new_n445), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G110), .B(G140), .ZN(new_n452));
  INV_X1    g266(.A(G227), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(G953), .ZN(new_n454));
  XOR2_X1   g268(.A(new_n452), .B(new_n454), .Z(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(KEYINPUT81), .B1(new_n313), .B2(new_n239), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT81), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n438), .A2(new_n459), .A3(new_n312), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n458), .A2(new_n439), .A3(new_n441), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n448), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT12), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT12), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n461), .A2(new_n448), .A3(new_n464), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n463), .A2(new_n450), .A3(new_n455), .A4(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(G902), .B1(new_n457), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G469), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(G469), .A2(G902), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n463), .A2(new_n450), .A3(new_n465), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n456), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n449), .A2(new_n450), .A3(new_n455), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(G469), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n469), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G221), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT9), .B(G234), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT78), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G902), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n476), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT97), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT96), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT15), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n485), .A3(G478), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n236), .A2(G128), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n190), .A2(G143), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OR2_X1    g303(.A1(new_n489), .A2(KEYINPUT94), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(KEYINPUT94), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(G134), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n490), .A2(G134), .A3(new_n491), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n215), .A2(G122), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n215), .A2(G122), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n498), .A3(new_n303), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  OR3_X1    g314(.A1(new_n498), .A2(KEYINPUT95), .A3(KEYINPUT14), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n498), .A2(KEYINPUT14), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT95), .B1(new_n498), .B2(KEYINPUT14), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n501), .A2(new_n497), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n500), .B1(new_n504), .B2(G107), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n496), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT13), .B1(new_n236), .B2(G128), .ZN(new_n507));
  OR2_X1    g321(.A1(new_n507), .A2(KEYINPUT93), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(KEYINPUT93), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n236), .A2(KEYINPUT13), .A3(G128), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n508), .A2(new_n509), .A3(new_n488), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(G134), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n303), .B1(new_n497), .B2(new_n498), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n494), .B(new_n512), .C1(new_n513), .C2(new_n500), .ZN(new_n514));
  INV_X1    g328(.A(G217), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n478), .A2(new_n515), .A3(G953), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n506), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n516), .B1(new_n506), .B2(new_n514), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n480), .B(new_n486), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n484), .B1(new_n485), .B2(G478), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n483), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n506), .A2(new_n514), .ZN(new_n523));
  INV_X1    g337(.A(new_n516), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(G902), .B1(new_n525), .B2(new_n517), .ZN(new_n526));
  INV_X1    g340(.A(new_n521), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n526), .A2(KEYINPUT97), .A3(new_n527), .A4(new_n486), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n518), .A2(new_n519), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n485), .B(G478), .C1(new_n529), .C2(G902), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n522), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n437), .A2(new_n475), .A3(new_n482), .A4(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n368), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n190), .A2(G119), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(KEYINPUT23), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n213), .A2(G128), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT75), .B(G110), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(KEYINPUT76), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n537), .A2(new_n535), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT24), .B(G110), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n374), .B(new_n388), .C1(new_n541), .C2(new_n544), .ZN(new_n545));
  XOR2_X1   g359(.A(new_n538), .B(KEYINPUT73), .Z(new_n546));
  INV_X1    g360(.A(G110), .ZN(new_n547));
  OAI221_X1 g361(.A(new_n404), .B1(new_n542), .B2(new_n543), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT22), .B(G137), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n428), .A2(G221), .A3(G234), .ZN(new_n551));
  XOR2_X1   g365(.A(new_n550), .B(new_n551), .Z(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n545), .A2(new_n548), .A3(new_n552), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n480), .A3(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT25), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(KEYINPUT77), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT77), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(KEYINPUT25), .ZN(new_n560));
  OR3_X1    g374(.A1(new_n556), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n554), .A2(new_n555), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n559), .B(KEYINPUT25), .C1(new_n562), .C2(G902), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n515), .B1(G234), .B2(new_n480), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n561), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n564), .A2(G902), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n554), .A2(new_n555), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n288), .A2(new_n534), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(new_n311), .ZN(G3));
  NAND3_X1  g385(.A1(new_n262), .A2(new_n255), .A3(new_n264), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT31), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(new_n265), .A3(new_n257), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n286), .B1(new_n574), .B2(new_n480), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT98), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n271), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n575), .A2(new_n577), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AND4_X1   g397(.A1(new_n569), .A2(new_n583), .A3(new_n482), .A4(new_n475), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT99), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n362), .A2(new_n585), .A3(new_n364), .ZN(new_n586));
  INV_X1    g400(.A(new_n366), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n360), .B1(new_n348), .B2(new_n358), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n587), .B1(new_n588), .B2(KEYINPUT99), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n419), .A2(new_n426), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(G478), .A2(G902), .ZN(new_n593));
  INV_X1    g407(.A(G478), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n526), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n525), .A2(KEYINPUT100), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n596), .B(KEYINPUT33), .C1(new_n518), .C2(new_n519), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n525), .B(new_n517), .C1(KEYINPUT100), .C2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n593), .B(new_n595), .C1(new_n600), .C2(new_n594), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n592), .A2(new_n601), .A3(new_n435), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n584), .A2(new_n590), .A3(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT34), .B(G104), .Z(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G6));
  INV_X1    g419(.A(KEYINPUT101), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n426), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g421(.A(KEYINPUT101), .B(G475), .C1(new_n425), .C2(G902), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n416), .A2(new_n418), .ZN(new_n609));
  AOI211_X1 g423(.A(new_n410), .B(new_n417), .C1(new_n413), .C2(new_n415), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n607), .B(new_n608), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(new_n532), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n612), .A2(new_n586), .A3(new_n589), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n584), .A2(new_n436), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(new_n303), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT102), .B(KEYINPUT35), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G9));
  NOR2_X1   g431(.A1(new_n553), .A2(KEYINPUT36), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n549), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n566), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n565), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n534), .A2(new_n579), .A3(new_n581), .A4(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(new_n547), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT103), .B(KEYINPUT37), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G12));
  AND2_X1   g439(.A1(new_n565), .A2(new_n620), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n286), .B1(new_n278), .B2(new_n283), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(new_n275), .ZN(new_n628));
  INV_X1    g442(.A(new_n270), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n272), .B1(new_n574), .B2(new_n187), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n626), .B1(new_n628), .B2(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n475), .A2(new_n482), .ZN(new_n633));
  INV_X1    g447(.A(G900), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n434), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n429), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n611), .A2(new_n532), .A3(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n632), .A2(new_n633), .A3(new_n590), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G128), .ZN(G30));
  NAND2_X1  g454(.A1(new_n591), .A2(new_n531), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n636), .B(KEYINPUT39), .Z(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n633), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n642), .B1(new_n645), .B2(KEYINPUT40), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(KEYINPUT40), .B2(new_n645), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n365), .A2(new_n367), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(KEYINPUT38), .Z(new_n649));
  NOR2_X1   g463(.A1(new_n621), .A2(new_n587), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n268), .A2(new_n256), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n480), .B1(new_n280), .B2(new_n255), .ZN(new_n652));
  OAI21_X1  g466(.A(G472), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n631), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n647), .A2(new_n649), .A3(new_n650), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G143), .ZN(G45));
  NOR3_X1   g470(.A1(new_n592), .A2(new_n601), .A3(new_n637), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n632), .A2(new_n633), .A3(new_n590), .A4(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G146), .ZN(G48));
  NAND2_X1  g473(.A1(KEYINPUT104), .A2(G469), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n467), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n660), .ZN(new_n662));
  AOI211_X1 g476(.A(G902), .B(new_n662), .C1(new_n457), .C2(new_n466), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n661), .A2(new_n663), .A3(new_n481), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n586), .A2(new_n664), .A3(new_n589), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n288), .A2(new_n569), .A3(new_n602), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT41), .B(G113), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT105), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n666), .B(new_n668), .ZN(G15));
  INV_X1    g483(.A(new_n664), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n435), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n288), .A2(new_n613), .A3(new_n569), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G116), .ZN(G18));
  NOR3_X1   g487(.A1(new_n591), .A2(new_n531), .A3(new_n435), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n288), .A2(new_n674), .A3(new_n621), .A4(new_n665), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G119), .ZN(G21));
  AND3_X1   g490(.A1(new_n642), .A2(new_n586), .A3(new_n589), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n574), .A2(new_n480), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n573), .B(new_n265), .C1(new_n255), .C2(new_n281), .ZN(new_n679));
  AOI22_X1  g493(.A1(new_n678), .A2(G472), .B1(new_n679), .B2(new_n187), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n677), .A2(new_n569), .A3(new_n671), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G122), .ZN(G24));
  INV_X1    g496(.A(new_n680), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n626), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n684), .A2(new_n657), .A3(new_n665), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G125), .ZN(G27));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n472), .B(KEYINPUT106), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(G469), .A3(new_n473), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n469), .A2(new_n470), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n481), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n587), .B1(new_n365), .B2(new_n367), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n288), .A2(new_n569), .A3(new_n691), .A4(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n657), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n687), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT107), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI211_X1 g511(.A(KEYINPUT107), .B(new_n687), .C1(new_n693), .C2(new_n694), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n285), .A2(new_n287), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(KEYINPUT108), .B2(new_n270), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n270), .A2(KEYINPUT108), .ZN(new_n702));
  INV_X1    g516(.A(new_n187), .ZN(new_n703));
  AOI211_X1 g517(.A(new_n256), .B(new_n241), .C1(new_n267), .C2(new_n226), .ZN(new_n704));
  AOI22_X1  g518(.A1(new_n704), .A2(new_n263), .B1(new_n256), .B2(new_n250), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n703), .B1(new_n705), .B2(new_n573), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n701), .B(new_n702), .C1(KEYINPUT32), .C2(new_n706), .ZN(new_n707));
  AND4_X1   g521(.A1(KEYINPUT42), .A2(new_n692), .A3(new_n657), .A4(new_n691), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n707), .A2(new_n569), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n699), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G131), .ZN(G33));
  INV_X1    g525(.A(new_n638), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n693), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n493), .ZN(G36));
  NOR2_X1   g528(.A1(new_n601), .A2(new_n591), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT43), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n716), .B(new_n621), .C1(new_n580), .C2(new_n582), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n688), .A2(KEYINPUT45), .A3(new_n473), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n472), .A2(new_n473), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n721), .A2(KEYINPUT45), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n720), .A2(G469), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT46), .B1(new_n723), .B2(new_n470), .ZN(new_n724));
  INV_X1    g538(.A(new_n469), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n723), .A2(KEYINPUT46), .A3(new_n470), .ZN(new_n727));
  AOI211_X1 g541(.A(new_n481), .B(new_n643), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n717), .A2(new_n718), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n719), .A2(new_n728), .A3(new_n692), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G137), .ZN(G39));
  NOR2_X1   g545(.A1(new_n288), .A2(new_n569), .ZN(new_n732));
  INV_X1    g546(.A(new_n692), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n694), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n726), .A2(new_n727), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT47), .B1(new_n735), .B2(new_n482), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT47), .ZN(new_n737));
  AOI211_X1 g551(.A(new_n737), .B(new_n481), .C1(new_n726), .C2(new_n727), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n732), .B(new_n734), .C1(new_n736), .C2(new_n738), .ZN(new_n739));
  XOR2_X1   g553(.A(KEYINPUT109), .B(G140), .Z(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G42));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n716), .A2(new_n430), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n683), .A2(new_n568), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n587), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n649), .A2(new_n670), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n742), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n743), .A2(new_n744), .ZN(new_n751));
  AOI21_X1  g565(.A(KEYINPUT112), .B1(new_n716), .B2(new_n430), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n746), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n755), .A2(KEYINPUT50), .A3(new_n587), .A4(new_n748), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n692), .A2(new_n664), .ZN(new_n757));
  NOR4_X1   g571(.A1(new_n654), .A2(new_n757), .A3(new_n568), .A4(new_n429), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n592), .A3(new_n601), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT114), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n759), .A2(KEYINPUT114), .ZN(new_n761));
  AOI22_X1  g575(.A1(new_n750), .A2(new_n756), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n757), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n745), .A2(new_n684), .A3(new_n763), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n746), .B(new_n692), .C1(new_n751), .C2(new_n752), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n736), .A2(new_n738), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n661), .A2(new_n663), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n482), .ZN(new_n772));
  OAI22_X1  g586(.A1(new_n767), .A2(new_n768), .B1(new_n769), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n762), .A2(new_n764), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n762), .A2(KEYINPUT51), .A3(new_n764), .A4(new_n773), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n745), .A2(new_n569), .A3(new_n707), .A4(new_n763), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT48), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n592), .A2(new_n601), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n758), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(G952), .A3(new_n428), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n780), .A2(new_n781), .A3(new_n784), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n776), .A2(new_n777), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n621), .A2(new_n637), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n654), .A2(new_n677), .A3(new_n691), .A4(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n639), .A2(new_n658), .A3(new_n685), .A4(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AND4_X1   g606(.A1(new_n288), .A2(new_n633), .A3(new_n590), .A4(new_n621), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n793), .B1(new_n638), .B2(new_n657), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n794), .A2(KEYINPUT52), .A3(new_n685), .A4(new_n789), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT53), .B1(new_n796), .B2(KEYINPUT111), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n666), .A2(new_n672), .A3(new_n675), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n622), .A2(new_n570), .A3(new_n681), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n782), .B1(new_n531), .B2(new_n592), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n800), .A2(new_n368), .A3(new_n435), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n583), .A2(new_n801), .A3(new_n569), .A4(new_n633), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n798), .A2(new_n799), .A3(new_n802), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n611), .A2(new_n531), .A3(new_n637), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n270), .B1(new_n706), .B2(new_n272), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n633), .B(new_n804), .C1(new_n700), .C2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n680), .A2(new_n657), .A3(new_n691), .ZN(new_n807));
  AOI211_X1 g621(.A(new_n626), .B(new_n733), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(KEYINPUT110), .B1(new_n808), .B2(new_n713), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n806), .A2(new_n807), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n621), .A3(new_n692), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT110), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n693), .A2(new_n712), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n803), .B1(new_n809), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n815), .A2(new_n796), .A3(new_n710), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n797), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n797), .A2(new_n816), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n787), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND4_X1   g633(.A1(KEYINPUT53), .A2(new_n815), .A3(new_n710), .A4(new_n796), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n792), .A2(new_n795), .B1(new_n699), .B2(new_n709), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT53), .B1(new_n821), .B2(new_n815), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n820), .A2(new_n822), .A3(KEYINPUT54), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n755), .A2(new_n665), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT115), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n786), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n827), .B1(G952), .B2(G953), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n771), .A2(KEYINPUT49), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n771), .A2(KEYINPUT49), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(new_n569), .A3(new_n366), .A4(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n831), .A2(new_n481), .A3(new_n654), .ZN(new_n832));
  INV_X1    g646(.A(new_n649), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(new_n833), .A3(new_n715), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n828), .A2(new_n834), .ZN(G75));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n816), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n821), .A2(KEYINPUT53), .A3(new_n815), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(G902), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(G210), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n337), .B1(new_n344), .B2(new_n347), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(new_n295), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT55), .ZN(new_n845));
  XOR2_X1   g659(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n846));
  AND3_X1   g660(.A1(new_n842), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT56), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n845), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n428), .A2(G952), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(G51));
  XOR2_X1   g665(.A(new_n470), .B(KEYINPUT117), .Z(new_n852));
  XOR2_X1   g666(.A(new_n852), .B(KEYINPUT57), .Z(new_n853));
  AOI21_X1  g667(.A(new_n787), .B1(new_n837), .B2(new_n838), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(new_n823), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n457), .A2(new_n466), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n853), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT54), .B1(new_n820), .B2(new_n822), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n837), .A2(new_n787), .A3(new_n838), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT118), .B1(new_n863), .B2(new_n857), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n840), .A2(new_n723), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n859), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n850), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(G54));
  NAND3_X1  g682(.A1(new_n841), .A2(KEYINPUT58), .A3(G475), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n413), .A2(new_n415), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n869), .A2(new_n871), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n872), .A2(new_n873), .A3(new_n850), .ZN(G60));
  XNOR2_X1  g688(.A(new_n600), .B(KEYINPUT119), .ZN(new_n875));
  XNOR2_X1  g689(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(new_n593), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n875), .B(new_n878), .C1(new_n861), .C2(new_n862), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n877), .B1(new_n819), .B2(new_n823), .ZN(new_n880));
  AOI211_X1 g694(.A(new_n850), .B(new_n879), .C1(new_n875), .C2(new_n880), .ZN(G63));
  NAND2_X1  g695(.A1(G217), .A2(G902), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT60), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n839), .A2(new_n619), .A3(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n884), .B1(new_n820), .B2(new_n822), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n850), .B1(new_n888), .B2(new_n562), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n839), .A2(KEYINPUT121), .A3(new_n619), .A4(new_n884), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT61), .B1(new_n889), .B2(KEYINPUT122), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n891), .B(new_n892), .ZN(G66));
  OAI21_X1  g707(.A(G953), .B1(new_n432), .B2(new_n292), .ZN(new_n894));
  INV_X1    g708(.A(new_n803), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n894), .B1(new_n895), .B2(G953), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT123), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n843), .B1(G898), .B2(new_n428), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n897), .B(new_n898), .ZN(G69));
  AND2_X1   g713(.A1(new_n699), .A2(new_n709), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n794), .A2(new_n685), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n707), .A2(new_n569), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n728), .A2(new_n677), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n739), .A2(new_n730), .A3(new_n813), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n428), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n428), .A2(G900), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n908), .A2(KEYINPUT125), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT125), .ZN(new_n912));
  AOI21_X1  g726(.A(G953), .B1(new_n905), .B2(new_n906), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n912), .B1(new_n913), .B2(new_n909), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n267), .B(new_n386), .Z(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(G953), .B1(new_n453), .B2(new_n634), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n739), .A2(new_n730), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n901), .A2(new_n655), .ZN(new_n920));
  XNOR2_X1  g734(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n800), .A2(new_n645), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n923), .A2(new_n288), .A3(new_n569), .A4(new_n692), .ZN(new_n924));
  NAND2_X1  g738(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n901), .A2(new_n655), .A3(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n919), .A2(new_n922), .A3(new_n924), .A4(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n916), .A2(G953), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n917), .A2(KEYINPUT126), .A3(new_n918), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n918), .A2(KEYINPUT126), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n918), .A2(KEYINPUT126), .ZN(new_n932));
  INV_X1    g746(.A(new_n916), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n911), .B2(new_n914), .ZN(new_n934));
  INV_X1    g748(.A(new_n929), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n931), .B(new_n932), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n930), .A2(new_n936), .ZN(G72));
  NAND2_X1  g751(.A1(new_n268), .A2(new_n256), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n907), .A2(new_n803), .ZN(new_n940));
  NAND2_X1  g754(.A1(G472), .A2(G902), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT63), .Z(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT127), .Z(new_n943));
  OAI21_X1  g757(.A(new_n939), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n927), .A2(new_n803), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n651), .B1(new_n945), .B2(new_n943), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n944), .A2(new_n946), .A3(new_n867), .ZN(new_n947));
  AOI211_X1 g761(.A(new_n651), .B(new_n939), .C1(new_n817), .C2(new_n818), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n947), .B1(new_n942), .B2(new_n948), .ZN(G57));
endmodule


