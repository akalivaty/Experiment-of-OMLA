//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 0 0 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967;
  XOR2_X1   g000(.A(G141gat), .B(G148gat), .Z(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  INV_X1    g002(.A(G162gat), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT2), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n202), .A2(KEYINPUT77), .A3(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G155gat), .B(G162gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND4_X1  g008(.A1(new_n202), .A2(KEYINPUT77), .A3(new_n207), .A4(new_n205), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G197gat), .B(G204gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT75), .B(G218gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(new_n214), .B2(KEYINPUT22), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G211gat), .ZN(new_n216));
  INV_X1    g015(.A(G211gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n213), .A2(KEYINPUT22), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G218gat), .ZN(new_n220));
  INV_X1    g019(.A(G218gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n216), .A2(new_n221), .A3(new_n218), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT84), .B1(new_n223), .B2(KEYINPUT29), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR3_X1   g025(.A1(new_n223), .A2(KEYINPUT84), .A3(KEYINPUT29), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n212), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G228gat), .A2(G233gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT78), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n211), .A2(new_n231), .A3(new_n225), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n209), .A2(new_n225), .A3(new_n210), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT78), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT29), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n223), .ZN(new_n236));
  OR2_X1    g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n228), .A2(new_n230), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT29), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(new_n239), .A3(new_n212), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n212), .A2(KEYINPUT3), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n240), .B(new_n241), .C1(new_n235), .C2(new_n236), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n229), .B(KEYINPUT82), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n242), .A2(KEYINPUT83), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT83), .B1(new_n242), .B2(new_n243), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n238), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G22gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT85), .ZN(new_n248));
  XOR2_X1   g047(.A(G78gat), .B(G106gat), .Z(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT31), .ZN(new_n250));
  INV_X1    g049(.A(G50gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G22gat), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n254), .B(new_n238), .C1(new_n244), .C2(new_n245), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n247), .A2(new_n248), .A3(new_n253), .A4(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n245), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT83), .A3(new_n243), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n228), .A2(new_n237), .ZN(new_n259));
  AOI22_X1  g058(.A1(new_n257), .A2(new_n258), .B1(new_n259), .B2(new_n230), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n260), .B(new_n254), .C1(KEYINPUT85), .C2(new_n252), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n246), .A2(G22gat), .A3(new_n252), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n256), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT5), .ZN(new_n265));
  INV_X1    g064(.A(G120gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G113gat), .ZN(new_n267));
  INV_X1    g066(.A(G113gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G120gat), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT1), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(G127gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G134gat), .ZN(new_n272));
  INV_X1    g071(.A(G127gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n270), .B(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G134gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(new_n212), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n211), .A2(new_n272), .A3(new_n276), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G225gat), .A2(G233gat), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n265), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n279), .A2(KEYINPUT4), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n232), .A2(new_n234), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(new_n277), .A3(new_n241), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n281), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n279), .A2(KEYINPUT4), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n283), .B(new_n284), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT80), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n284), .A2(new_n290), .A3(new_n288), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n279), .A2(KEYINPUT80), .A3(KEYINPUT4), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n282), .A2(KEYINPUT5), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n291), .A2(new_n286), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(G1gat), .B(G29gat), .Z(new_n296));
  XNOR2_X1  g095(.A(G57gat), .B(G85gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n299));
  XOR2_X1   g098(.A(new_n298), .B(new_n299), .Z(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT6), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT28), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n306), .A2(G190gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n310));
  NOR3_X1   g109(.A1(new_n309), .A2(new_n310), .A3(KEYINPUT65), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT65), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT27), .ZN(new_n313));
  INV_X1    g112(.A(G183gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n312), .B1(new_n315), .B2(new_n308), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n307), .B1(new_n311), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT66), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(KEYINPUT64), .B(G183gat), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n310), .B1(new_n320), .B2(KEYINPUT27), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n306), .B1(new_n321), .B2(G190gat), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT65), .B1(new_n309), .B2(new_n310), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n315), .A2(new_n312), .A3(new_n308), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n325), .A2(KEYINPUT66), .A3(new_n307), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n319), .A2(new_n322), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(G169gat), .A2(G176gat), .ZN(new_n329));
  OR3_X1    g128(.A1(new_n328), .A2(new_n329), .A3(KEYINPUT67), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT26), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT67), .B1(new_n328), .B2(new_n329), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n327), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n335), .B(KEYINPUT24), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(G183gat), .B2(G190gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n329), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n341), .A2(new_n342), .B1(G169gat), .B2(G176gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT25), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n320), .ZN(new_n347));
  INV_X1    g146(.A(G190gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n345), .B1(new_n349), .B2(new_n338), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n343), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G226gat), .A2(G233gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n239), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT68), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n327), .A2(new_n358), .A3(new_n336), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(new_n327), .B2(new_n336), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n352), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n357), .B1(new_n361), .B2(new_n354), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n236), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n356), .ZN(new_n364));
  OR2_X1    g163(.A1(new_n353), .A2(new_n354), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n365), .A3(new_n223), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n363), .A2(new_n366), .A3(KEYINPUT76), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n364), .A2(new_n368), .A3(new_n365), .A4(new_n223), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G8gat), .B(G36gat), .ZN(new_n371));
  INV_X1    g170(.A(G64gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(G92gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n370), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n302), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n303), .B1(new_n295), .B2(new_n301), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n305), .B(new_n377), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT86), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n367), .A2(new_n369), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n381), .B1(new_n382), .B2(KEYINPUT37), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT37), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n370), .A2(KEYINPUT86), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n367), .A2(KEYINPUT37), .A3(new_n369), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n375), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT87), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n387), .A2(KEYINPUT87), .A3(new_n375), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n386), .A2(KEYINPUT38), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n362), .A2(new_n223), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n364), .A2(new_n365), .A3(new_n236), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(KEYINPUT37), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT86), .B1(new_n370), .B2(new_n384), .ZN(new_n396));
  AOI211_X1 g195(.A(new_n381), .B(KEYINPUT37), .C1(new_n367), .C2(new_n369), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n375), .B(new_n395), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT38), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n380), .B1(new_n392), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n382), .A2(new_n375), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(KEYINPUT30), .A3(new_n377), .ZN(new_n403));
  OR3_X1    g202(.A1(new_n382), .A2(KEYINPUT30), .A3(new_n375), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n291), .A2(new_n286), .A3(new_n292), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n282), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n300), .B1(new_n407), .B2(KEYINPUT39), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n278), .A2(new_n279), .A3(new_n281), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n408), .B1(KEYINPUT39), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT40), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n302), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n411), .A2(KEYINPUT40), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n405), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n264), .B1(new_n401), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT81), .B1(new_n295), .B2(new_n301), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT81), .ZN(new_n418));
  AOI211_X1 g217(.A(new_n418), .B(new_n300), .C1(new_n289), .C2(new_n294), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n379), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n304), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n422), .B1(new_n404), .B2(new_n403), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n263), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n416), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n361), .A2(new_n277), .ZN(new_n426));
  NAND2_X1  g225(.A1(G227gat), .A2(G233gat), .ZN(new_n427));
  INV_X1    g226(.A(new_n277), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n428), .B(new_n352), .C1(new_n359), .C2(new_n360), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT72), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT34), .ZN(new_n433));
  INV_X1    g232(.A(new_n427), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n337), .A2(KEYINPUT68), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n327), .A2(new_n358), .A3(new_n336), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n428), .B1(new_n437), .B2(new_n352), .ZN(new_n438));
  INV_X1    g237(.A(new_n429), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n434), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(KEYINPUT69), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT69), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n427), .B1(new_n426), .B2(new_n429), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n443), .B1(new_n444), .B2(KEYINPUT33), .ZN(new_n445));
  XNOR2_X1  g244(.A(KEYINPUT70), .B(G71gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(G99gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(G15gat), .B(G43gat), .ZN(new_n448));
  XOR2_X1   g247(.A(new_n447), .B(new_n448), .Z(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n440), .A2(KEYINPUT32), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n442), .A2(new_n445), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n440), .B(KEYINPUT32), .C1(new_n441), .C2(new_n449), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT71), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT71), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n452), .A2(new_n456), .A3(new_n453), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n433), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n433), .A2(new_n452), .A3(new_n453), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT36), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT73), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n433), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n454), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT74), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(new_n464), .A3(new_n459), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT36), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n454), .A2(new_n462), .A3(KEYINPUT74), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n452), .A2(new_n456), .A3(new_n453), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n456), .B1(new_n452), .B2(new_n453), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n462), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n460), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT73), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n461), .A2(new_n468), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n425), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n459), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n263), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n423), .A2(new_n478), .A3(new_n471), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT35), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n467), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n305), .B1(new_n378), .B2(new_n379), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT35), .B1(new_n403), .B2(new_n404), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n481), .A2(new_n482), .A3(new_n264), .A4(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n476), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT18), .ZN(new_n487));
  XNOR2_X1  g286(.A(G15gat), .B(G22gat), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT16), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n488), .B1(new_n489), .B2(G1gat), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n490), .B1(G1gat), .B2(new_n488), .ZN(new_n491));
  INV_X1    g290(.A(G8gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(G43gat), .B(G50gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT15), .ZN(new_n495));
  OR3_X1    g294(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT88), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n496), .A2(new_n497), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G29gat), .A2(G36gat), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n495), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n494), .A2(KEYINPUT15), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT89), .B1(new_n494), .B2(KEYINPUT15), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT90), .B1(G29gat), .B2(G36gat), .ZN(new_n507));
  AND3_X1   g306(.A1(KEYINPUT90), .A2(G29gat), .A3(G36gat), .ZN(new_n508));
  AOI211_X1 g307(.A(new_n507), .B(new_n508), .C1(new_n496), .C2(new_n499), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT91), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT91), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n506), .A2(new_n512), .A3(new_n509), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n503), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT17), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI211_X1 g315(.A(KEYINPUT17), .B(new_n503), .C1(new_n511), .C2(new_n513), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n493), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n514), .A2(new_n493), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G229gat), .A2(G233gat), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n487), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(KEYINPUT11), .B(G169gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(G197gat), .ZN(new_n526));
  XOR2_X1   g325(.A(G113gat), .B(G141gat), .Z(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT12), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n522), .B(KEYINPUT13), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n514), .A2(new_n493), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n531), .B1(new_n532), .B2(new_n519), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n518), .A2(KEYINPUT18), .A3(new_n520), .A4(new_n522), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n524), .A2(new_n529), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT92), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n524), .A2(new_n533), .A3(new_n534), .ZN(new_n538));
  INV_X1    g337(.A(new_n529), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G134gat), .B(G162gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(G190gat), .B(G218gat), .ZN(new_n543));
  AND2_X1   g342(.A1(G232gat), .A2(G233gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT41), .ZN(new_n545));
  NAND2_X1  g344(.A1(G85gat), .A2(G92gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT7), .ZN(new_n547));
  INV_X1    g346(.A(G99gat), .ZN(new_n548));
  INV_X1    g347(.A(G106gat), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT8), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n547), .B(new_n550), .C1(G85gat), .C2(G92gat), .ZN(new_n551));
  XOR2_X1   g350(.A(G99gat), .B(G106gat), .Z(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n545), .B1(new_n514), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT98), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n544), .A2(KEYINPUT41), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n553), .B1(new_n516), .B2(new_n517), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n555), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n557), .B1(new_n555), .B2(new_n558), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n543), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n561), .ZN(new_n563));
  INV_X1    g362(.A(new_n543), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(new_n559), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n542), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n562), .A2(new_n565), .A3(new_n542), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G127gat), .B(G155gat), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n570), .B(KEYINPUT20), .Z(new_n571));
  OR2_X1    g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(G71gat), .A2(G78gat), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n573), .B(KEYINPUT93), .Z(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT94), .B(G64gat), .ZN(new_n575));
  INV_X1    g374(.A(G57gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n572), .B(new_n574), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n578), .B1(new_n572), .B2(new_n573), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n372), .B1(new_n576), .B2(KEYINPUT95), .ZN(new_n582));
  OR3_X1    g381(.A1(new_n576), .A2(new_n372), .A3(KEYINPUT95), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n579), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n580), .B1(new_n579), .B2(new_n584), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT21), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n217), .B1(new_n588), .B2(new_n493), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n587), .A2(KEYINPUT21), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n588), .A2(new_n217), .A3(new_n493), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n591), .B1(new_n590), .B2(new_n592), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n571), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n595), .ZN(new_n597));
  INV_X1    g396(.A(new_n571), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(new_n593), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT19), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT97), .B(G183gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  AND3_X1   g402(.A1(new_n596), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n603), .B1(new_n596), .B2(new_n599), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT99), .B1(new_n569), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT99), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n567), .A2(new_n606), .A3(new_n568), .A4(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G120gat), .B(G148gat), .ZN(new_n611));
  INV_X1    g410(.A(G176gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n613), .B(G204gat), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT102), .ZN(new_n615));
  INV_X1    g414(.A(new_n553), .ZN(new_n616));
  OAI211_X1 g415(.A(KEYINPUT10), .B(new_n616), .C1(new_n585), .C2(new_n586), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n617), .A2(KEYINPUT100), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(KEYINPUT100), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n553), .B1(new_n579), .B2(new_n584), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n620), .B1(new_n587), .B2(new_n553), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n618), .B(new_n619), .C1(new_n621), .C2(KEYINPUT10), .ZN(new_n622));
  NAND2_X1  g421(.A1(G230gat), .A2(G233gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n623), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n615), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n628), .B1(new_n622), .B2(new_n623), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT101), .ZN(new_n631));
  INV_X1    g430(.A(new_n614), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n631), .B1(new_n630), .B2(new_n632), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n629), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n608), .A2(new_n610), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n486), .A2(new_n541), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT103), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n422), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G1gat), .ZN(G1324gat));
  INV_X1    g442(.A(new_n405), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n489), .A2(new_n492), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n489), .A2(new_n492), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n641), .A2(new_n644), .A3(new_n646), .A4(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT104), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT105), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT42), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n641), .A2(new_n644), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(G8gat), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT42), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n654), .B1(new_n648), .B2(KEYINPUT105), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT105), .B1(new_n648), .B2(KEYINPUT104), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n651), .B(new_n653), .C1(new_n655), .C2(new_n656), .ZN(G1325gat));
  AOI21_X1  g456(.A(G15gat), .B1(new_n641), .B2(new_n481), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT106), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n475), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n461), .A2(new_n468), .A3(new_n474), .A4(KEYINPUT106), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n641), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n658), .B1(G15gat), .B2(new_n664), .ZN(G1326gat));
  NAND2_X1  g464(.A1(new_n641), .A2(new_n263), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT43), .B(G22gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1327gat));
  NAND2_X1  g467(.A1(new_n486), .A2(new_n541), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n567), .A2(new_n568), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n607), .A2(new_n637), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n422), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n673), .A2(G29gat), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(KEYINPUT45), .Z(new_n676));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n480), .A2(new_n484), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n678), .B1(new_n662), .B2(new_n425), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n677), .B1(new_n679), .B2(new_n670), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT107), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n537), .A2(new_n681), .A3(new_n540), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n681), .B1(new_n537), .B2(new_n540), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(new_n671), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n486), .A2(KEYINPUT44), .A3(new_n569), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n680), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(G29gat), .B1(new_n689), .B2(new_n674), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n676), .A2(new_n690), .ZN(G1328gat));
  NOR3_X1   g490(.A1(new_n673), .A2(G36gat), .A3(new_n405), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT46), .ZN(new_n693));
  OAI21_X1  g492(.A(G36gat), .B1(new_n689), .B2(new_n405), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(G1329gat));
  NAND3_X1  g494(.A1(new_n688), .A2(G43gat), .A3(new_n663), .ZN(new_n696));
  INV_X1    g495(.A(new_n481), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n673), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n696), .B1(new_n698), .B2(G43gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g499(.A1(new_n680), .A2(new_n263), .A3(new_n687), .A4(new_n686), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(G50gat), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n702), .A2(KEYINPUT108), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT48), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n672), .A2(new_n251), .A3(new_n263), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n706), .B1(new_n702), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n702), .A2(new_n707), .A3(new_n706), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n705), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n710), .ZN(new_n712));
  OAI22_X1  g511(.A1(new_n712), .A2(new_n708), .B1(new_n703), .B2(new_n704), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(G1331gat));
  INV_X1    g513(.A(new_n685), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n679), .A2(new_n715), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n608), .A2(new_n610), .A3(new_n636), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(new_n674), .ZN(new_n719));
  XOR2_X1   g518(.A(KEYINPUT110), .B(G57gat), .Z(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1332gat));
  XNOR2_X1  g520(.A(new_n405), .B(KEYINPUT111), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  AND2_X1   g524(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(new_n724), .B2(new_n725), .ZN(G1333gat));
  INV_X1    g527(.A(new_n718), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n729), .A2(G71gat), .A3(new_n663), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n718), .A2(new_n697), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(G71gat), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g532(.A1(new_n729), .A2(new_n263), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g534(.A1(new_n715), .A2(new_n606), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n680), .A2(new_n636), .A3(new_n687), .A4(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(G85gat), .B1(new_n737), .B2(new_n674), .ZN(new_n738));
  AOI22_X1  g537(.A1(new_n660), .A2(new_n661), .B1(new_n416), .B2(new_n424), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n569), .B(new_n736), .C1(new_n739), .C2(new_n678), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT51), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n637), .A2(G85gat), .A3(new_n674), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT112), .Z(new_n746));
  OAI21_X1  g545(.A(new_n738), .B1(new_n744), .B2(new_n746), .ZN(G1336gat));
  NOR2_X1   g546(.A1(new_n744), .A2(new_n637), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n723), .A2(G92gat), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751));
  OAI21_X1  g550(.A(G92gat), .B1(new_n737), .B2(new_n723), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  AND4_X1   g552(.A1(new_n636), .A2(new_n680), .A3(new_n687), .A4(new_n736), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n374), .B1(new_n754), .B2(new_n644), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT113), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n742), .B2(new_n743), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n756), .B1(new_n740), .B2(new_n741), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n637), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n755), .B1(new_n760), .B2(new_n749), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n753), .B1(new_n761), .B2(new_n751), .ZN(G1337gat));
  NOR3_X1   g561(.A1(new_n737), .A2(new_n548), .A3(new_n662), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n481), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n764), .B2(new_n548), .ZN(G1338gat));
  NOR2_X1   g564(.A1(new_n264), .A2(G106gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n636), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n767), .B1(new_n757), .B2(new_n759), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n549), .B1(new_n754), .B2(new_n263), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT53), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n771));
  OAI21_X1  g570(.A(G106gat), .B1(new_n737), .B2(new_n264), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n636), .B(new_n766), .C1(new_n742), .C2(new_n743), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n770), .A2(new_n771), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n767), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n662), .A2(new_n425), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n485), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n779), .A2(KEYINPUT51), .A3(new_n569), .A4(new_n736), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n740), .A2(new_n741), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT113), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n777), .B1(new_n782), .B2(new_n758), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n773), .B1(new_n783), .B2(new_n772), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n785));
  OAI21_X1  g584(.A(KEYINPUT114), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n776), .A2(new_n786), .ZN(G1339gat));
  OAI21_X1  g586(.A(KEYINPUT54), .B1(new_n622), .B2(new_n623), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n625), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n614), .B1(new_n624), .B2(KEYINPUT54), .ZN(new_n791));
  OR3_X1    g590(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n635), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n633), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n790), .B1(new_n789), .B2(new_n791), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n792), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n541), .A2(KEYINPUT107), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n796), .B1(new_n797), .B2(new_n682), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799));
  INV_X1    g598(.A(new_n521), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n800), .B2(new_n522), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n521), .A2(KEYINPUT115), .A3(new_n523), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n532), .A2(new_n519), .A3(new_n531), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n528), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n535), .A2(new_n536), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n535), .A2(new_n536), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n636), .B(new_n805), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n670), .B1(new_n798), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n537), .A2(new_n805), .ZN(new_n812));
  INV_X1    g611(.A(new_n796), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n569), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n606), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n685), .A2(new_n608), .A3(new_n610), .A4(new_n637), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(new_n697), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n722), .A2(new_n674), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(new_n264), .A3(new_n820), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n535), .A2(new_n536), .ZN(new_n822));
  AOI22_X1  g621(.A1(new_n822), .A2(new_n806), .B1(new_n539), .B2(new_n538), .ZN(new_n823));
  OAI21_X1  g622(.A(G113gat), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n813), .B1(new_n683), .B2(new_n684), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n569), .B1(new_n825), .B2(new_n809), .ZN(new_n826));
  INV_X1    g625(.A(new_n814), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n607), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n816), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n458), .A2(new_n477), .A3(new_n263), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n422), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(new_n722), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n715), .A2(new_n268), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT116), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n824), .B1(new_n833), .B2(new_n835), .ZN(G1340gat));
  NAND3_X1  g635(.A1(new_n832), .A2(new_n266), .A3(new_n636), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n637), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n837), .B1(new_n838), .B2(new_n266), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT117), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n837), .B(new_n841), .C1(new_n838), .C2(new_n266), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(G1341gat));
  NOR3_X1   g642(.A1(new_n821), .A2(new_n273), .A3(new_n607), .ZN(new_n844));
  AOI21_X1  g643(.A(G127gat), .B1(new_n832), .B2(new_n606), .ZN(new_n845));
  OR3_X1    g644(.A1(new_n844), .A2(new_n845), .A3(KEYINPUT118), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT118), .B1(new_n844), .B2(new_n845), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(G1342gat));
  INV_X1    g647(.A(new_n831), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n569), .A2(new_n405), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT119), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n275), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT56), .ZN(new_n853));
  OAI21_X1  g652(.A(G134gat), .B1(new_n821), .B2(new_n670), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT56), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n849), .A2(new_n855), .A3(new_n275), .A4(new_n851), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT120), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n853), .A2(new_n854), .A3(new_n859), .A4(new_n856), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(G1343gat));
  INV_X1    g660(.A(G141gat), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n818), .A2(new_n674), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n663), .A2(new_n264), .ZN(new_n864));
  AND4_X1   g663(.A1(new_n862), .A2(new_n863), .A3(new_n723), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n541), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT58), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n809), .B1(new_n823), .B2(new_n796), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n670), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n606), .B1(new_n870), .B2(new_n814), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n816), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI211_X1 g672(.A(KEYINPUT122), .B(new_n606), .C1(new_n870), .C2(new_n814), .ZN(new_n874));
  OAI211_X1 g673(.A(KEYINPUT57), .B(new_n263), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n264), .B1(new_n828), .B2(new_n816), .ZN(new_n876));
  XOR2_X1   g675(.A(KEYINPUT121), .B(KEYINPUT57), .Z(new_n877));
  OAI21_X1  g676(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n662), .A2(new_n820), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n862), .B1(new_n880), .B2(new_n541), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n878), .A2(new_n715), .A3(new_n879), .ZN(new_n882));
  AOI22_X1  g681(.A1(new_n865), .A2(new_n541), .B1(new_n882), .B2(G141gat), .ZN(new_n883));
  OAI22_X1  g682(.A1(new_n868), .A2(new_n881), .B1(new_n883), .B2(new_n867), .ZN(G1344gat));
  NAND3_X1  g683(.A1(new_n878), .A2(new_n636), .A3(new_n879), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n886), .A3(G148gat), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT123), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n263), .B(new_n877), .C1(new_n815), .C2(new_n817), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n638), .A2(new_n541), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n263), .B1(new_n890), .B2(new_n871), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n637), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n894), .A2(new_n879), .ZN(new_n895));
  INV_X1    g694(.A(G148gat), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT59), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n885), .A2(new_n898), .A3(new_n886), .A4(G148gat), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n888), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n863), .A2(new_n864), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n901), .A2(new_n723), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n896), .A3(new_n636), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n900), .A2(new_n903), .ZN(G1345gat));
  AOI21_X1  g703(.A(G155gat), .B1(new_n902), .B2(new_n606), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n607), .A2(new_n203), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n905), .B1(new_n880), .B2(new_n906), .ZN(G1346gat));
  NAND3_X1  g706(.A1(new_n901), .A2(new_n204), .A3(new_n851), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n880), .A2(new_n569), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n909), .B2(new_n204), .ZN(G1347gat));
  NAND4_X1  g709(.A1(new_n829), .A2(new_n674), .A3(new_n830), .A4(new_n722), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(G169gat), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n913), .A3(new_n715), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n819), .A2(new_n264), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n644), .A2(new_n674), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n915), .A2(new_n823), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n914), .B1(new_n917), .B2(new_n913), .ZN(G1348gat));
  AOI21_X1  g717(.A(G176gat), .B1(new_n912), .B2(new_n636), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n915), .A2(new_n916), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n637), .A2(new_n612), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(G1349gat));
  NAND3_X1  g721(.A1(new_n912), .A2(new_n325), .A3(new_n606), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n915), .A2(new_n607), .A3(new_n916), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n924), .B2(new_n347), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT60), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n923), .B(new_n927), .C1(new_n924), .C2(new_n347), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(G1350gat));
  NOR3_X1   g728(.A1(new_n915), .A2(new_n670), .A3(new_n916), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n930), .A2(new_n348), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n931), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n912), .A2(new_n348), .A3(new_n569), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n932), .B(new_n933), .C1(new_n930), .C2(new_n348), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(G1351gat));
  AOI211_X1 g738(.A(new_n663), .B(new_n916), .C1(new_n889), .C2(new_n893), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(new_n541), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT126), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n940), .A2(new_n943), .A3(new_n541), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n942), .A2(G197gat), .A3(new_n944), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n663), .A2(new_n264), .A3(new_n723), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT125), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n818), .A2(new_n422), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n685), .A2(G197gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n945), .B1(new_n949), .B2(new_n950), .ZN(G1352gat));
  XOR2_X1   g750(.A(KEYINPUT127), .B(G204gat), .Z(new_n952));
  NOR3_X1   g751(.A1(new_n949), .A2(new_n637), .A3(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n894), .A2(new_n674), .A3(new_n644), .A4(new_n662), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(new_n952), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n953), .A2(new_n954), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n955), .A2(new_n957), .A3(new_n958), .ZN(G1353gat));
  INV_X1    g758(.A(new_n949), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n960), .A2(new_n217), .A3(new_n606), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n940), .A2(new_n606), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n962), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT63), .B1(new_n962), .B2(G211gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1354gat));
  AOI21_X1  g764(.A(G218gat), .B1(new_n960), .B2(new_n569), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n569), .A2(new_n214), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n966), .B1(new_n940), .B2(new_n967), .ZN(G1355gat));
endmodule


