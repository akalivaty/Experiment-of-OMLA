//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 0 1 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT0), .A2(G128), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G143), .B(G146), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n194), .B1(KEYINPUT0), .B2(G128), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n192), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT0), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  AOI21_X1  g017(.A(KEYINPUT64), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n201), .A2(new_n191), .A3(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n196), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G125), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(KEYINPUT88), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n207), .A2(KEYINPUT88), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n193), .A2(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n203), .B1(new_n198), .B2(KEYINPUT1), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(new_n193), .ZN(new_n213));
  OR2_X1    g027(.A1(new_n213), .A2(G125), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n208), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G953), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G224), .ZN(new_n217));
  XOR2_X1   g031(.A(new_n215), .B(new_n217), .Z(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT86), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT6), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(KEYINPUT78), .A2(G104), .ZN(new_n224));
  NOR2_X1   g038(.A1(KEYINPUT78), .A2(G104), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(G101), .B1(new_n226), .B2(G107), .ZN(new_n227));
  INV_X1    g041(.A(G107), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n228), .B1(new_n224), .B2(new_n225), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT3), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(new_n228), .A3(G104), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT79), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT79), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n234), .A2(new_n231), .A3(new_n228), .A4(G104), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n227), .A2(new_n230), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G101), .ZN(new_n238));
  INV_X1    g052(.A(G104), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G107), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n238), .B1(new_n229), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(G116), .B(G119), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT5), .ZN(new_n245));
  INV_X1    g059(.A(G119), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G116), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n245), .B(G113), .C1(KEYINPUT5), .C2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT2), .ZN(new_n250));
  INV_X1    g064(.A(G113), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(KEYINPUT2), .A2(G113), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(new_n244), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n248), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n243), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT80), .ZN(new_n259));
  AOI22_X1  g073(.A1(KEYINPUT3), .A2(new_n229), .B1(new_n233), .B2(new_n235), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n226), .A2(G107), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n238), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n237), .A2(KEYINPUT4), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n259), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n265), .B1(new_n260), .B2(new_n227), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n230), .A2(new_n236), .A3(new_n261), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G101), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n266), .A2(new_n268), .A3(KEYINPUT80), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n254), .A2(new_n255), .A3(new_n244), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n244), .B1(new_n254), .B2(new_n255), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n253), .ZN(new_n275));
  NOR3_X1   g089(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n255), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n244), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(new_n256), .A3(KEYINPUT68), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n265), .A2(new_n262), .B1(new_n274), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n258), .B1(new_n270), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(G110), .B(G122), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n223), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n266), .A2(new_n268), .A3(KEYINPUT80), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT80), .B1(new_n266), .B2(new_n268), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n281), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n258), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n283), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(new_n290), .A3(new_n222), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n287), .A2(new_n283), .A3(new_n288), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT87), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n282), .A2(KEYINPUT87), .A3(new_n283), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n296), .A3(KEYINPUT6), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n219), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n295), .A2(new_n296), .ZN(new_n299));
  XOR2_X1   g113(.A(new_n283), .B(KEYINPUT8), .Z(new_n300));
  NAND2_X1  g114(.A1(new_n243), .A2(new_n257), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n300), .B1(new_n288), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n215), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n217), .A2(KEYINPUT7), .ZN(new_n304));
  NAND2_X1  g118(.A1(KEYINPUT89), .A2(KEYINPUT7), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  OAI211_X1 g120(.A(KEYINPUT7), .B(new_n217), .C1(new_n215), .C2(KEYINPUT89), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n302), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n299), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G902), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n190), .B1(new_n298), .B2(new_n311), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n295), .A2(new_n296), .A3(KEYINPUT6), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n284), .A2(new_n291), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n218), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(G902), .B1(new_n299), .B2(new_n308), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n189), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n188), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G469), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(new_n310), .ZN(new_n321));
  XNOR2_X1  g135(.A(G110), .B(G140), .ZN(new_n322));
  INV_X1    g136(.A(G227), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(G953), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n322), .B(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n241), .B1(new_n260), .B2(new_n227), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(KEYINPUT10), .A3(new_n213), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT1), .B1(new_n199), .B2(G146), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT81), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n198), .A2(KEYINPUT81), .A3(KEYINPUT1), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(G128), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n201), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n211), .ZN(new_n334));
  AOI211_X1 g148(.A(KEYINPUT82), .B(KEYINPUT10), .C1(new_n326), .C2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT82), .ZN(new_n336));
  INV_X1    g150(.A(new_n211), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n203), .B1(new_n328), .B2(new_n329), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n193), .B1(new_n338), .B2(new_n331), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n237), .B(new_n242), .C1(new_n337), .C2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT10), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n336), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n327), .B1(new_n335), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT69), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n193), .A2(new_n192), .A3(new_n195), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n191), .B1(new_n201), .B2(new_n204), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n196), .A2(new_n205), .A3(KEYINPUT69), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n349), .B1(KEYINPUT4), .B2(new_n268), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n350), .B1(new_n264), .B2(new_n269), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT11), .ZN(new_n352));
  INV_X1    g166(.A(G134), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n352), .B1(new_n353), .B2(G137), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(G137), .ZN(new_n355));
  INV_X1    g169(.A(G137), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(KEYINPUT11), .A3(G134), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n354), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT65), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(G131), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(G131), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n354), .A2(new_n357), .A3(new_n361), .A4(new_n355), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n343), .A2(new_n351), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n363), .ZN(new_n365));
  INV_X1    g179(.A(new_n327), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n337), .B1(new_n332), .B2(new_n201), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n341), .B1(new_n243), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT82), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n340), .A2(new_n336), .A3(new_n341), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n366), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n262), .A2(new_n265), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n349), .B(new_n372), .C1(new_n285), .C2(new_n286), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n365), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n325), .B1(new_n364), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n213), .B1(new_n237), .B2(new_n242), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT83), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n340), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NOR3_X1   g192(.A1(new_n326), .A2(KEYINPUT83), .A3(new_n213), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n363), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT12), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI211_X1 g196(.A(KEYINPUT12), .B(new_n363), .C1(new_n378), .C2(new_n379), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n371), .A2(new_n365), .A3(new_n373), .ZN(new_n385));
  INV_X1    g199(.A(new_n325), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(G902), .B1(new_n375), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n321), .B1(new_n388), .B2(new_n320), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT84), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n363), .B1(new_n343), .B2(new_n351), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n391), .A2(new_n385), .A3(new_n386), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n386), .B1(new_n384), .B2(new_n385), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n390), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(new_n385), .A3(new_n386), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n343), .A2(new_n351), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n396), .A2(new_n365), .B1(new_n383), .B2(new_n382), .ZN(new_n397));
  OAI211_X1 g211(.A(KEYINPUT84), .B(new_n395), .C1(new_n397), .C2(new_n386), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n394), .A2(new_n398), .A3(G469), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n389), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT9), .B(G234), .ZN(new_n401));
  OAI21_X1  g215(.A(G221), .B1(new_n401), .B2(G902), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT85), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT85), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n400), .A2(new_n405), .A3(new_n402), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n319), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(G113), .B(G122), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n408), .B(new_n239), .ZN(new_n409));
  XNOR2_X1  g223(.A(G125), .B(G140), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(new_n197), .ZN(new_n411));
  NOR2_X1   g225(.A1(G237), .A2(G953), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(G143), .A3(G214), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(G143), .B1(new_n412), .B2(G214), .ZN(new_n415));
  OAI211_X1 g229(.A(KEYINPUT18), .B(G131), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n415), .ZN(new_n417));
  NAND2_X1  g231(.A1(KEYINPUT18), .A2(G131), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n413), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n411), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n410), .A2(KEYINPUT16), .ZN(new_n421));
  INV_X1    g235(.A(G125), .ZN(new_n422));
  OR3_X1    g236(.A1(new_n422), .A2(KEYINPUT16), .A3(G140), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n197), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n421), .A2(G146), .A3(new_n423), .ZN(new_n426));
  OAI21_X1  g240(.A(G131), .B1(new_n414), .B2(new_n415), .ZN(new_n427));
  INV_X1    g241(.A(G131), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n417), .A2(new_n428), .A3(new_n413), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n425), .B(new_n426), .C1(new_n430), .C2(KEYINPUT17), .ZN(new_n431));
  OAI211_X1 g245(.A(KEYINPUT17), .B(G131), .C1(new_n414), .C2(new_n415), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(KEYINPUT91), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n409), .B(new_n420), .C1(new_n431), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n430), .A2(new_n426), .ZN(new_n435));
  NAND2_X1  g249(.A1(KEYINPUT90), .A2(KEYINPUT19), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(KEYINPUT90), .A2(KEYINPUT19), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n410), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n410), .A2(KEYINPUT90), .A3(KEYINPUT19), .ZN(new_n441));
  AOI21_X1  g255(.A(G146), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n420), .B1(new_n435), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n409), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n434), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(G475), .A2(G902), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT20), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT20), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n446), .A2(new_n450), .A3(new_n447), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n420), .B1(new_n431), .B2(new_n433), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(new_n409), .ZN(new_n454));
  OAI21_X1  g268(.A(G475), .B1(new_n454), .B2(G902), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G128), .B(G143), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT13), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n199), .A2(G128), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n458), .B(G134), .C1(KEYINPUT13), .C2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G116), .B(G122), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(new_n228), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n457), .A2(new_n353), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n457), .A2(new_n353), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n465), .A2(KEYINPUT92), .A3(new_n463), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT14), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G122), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(G116), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n228), .B1(new_n470), .B2(KEYINPUT14), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n468), .A2(new_n471), .B1(new_n228), .B2(new_n461), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT92), .B1(new_n465), .B2(new_n463), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n464), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G217), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n401), .A2(new_n476), .A3(G953), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n475), .A2(new_n478), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n310), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G478), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(KEYINPUT15), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n481), .B(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G952), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n485), .A2(KEYINPUT93), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(KEYINPUT93), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n216), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n488), .B1(G234), .B2(G237), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(G234), .A2(G237), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(G902), .A3(G953), .ZN(new_n492));
  XOR2_X1   g306(.A(new_n492), .B(KEYINPUT94), .Z(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT21), .B(G898), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n490), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT95), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NOR3_X1   g312(.A1(new_n456), .A2(new_n484), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n407), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n476), .B1(G234), .B2(new_n310), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT23), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n503), .B1(new_n246), .B2(G128), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n203), .A2(KEYINPUT23), .A3(G119), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n504), .B(new_n505), .C1(G119), .C2(new_n203), .ZN(new_n506));
  XNOR2_X1  g320(.A(G119), .B(G128), .ZN(new_n507));
  XOR2_X1   g321(.A(KEYINPUT24), .B(G110), .Z(new_n508));
  OAI22_X1  g322(.A1(new_n506), .A2(G110), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n410), .A2(new_n197), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n426), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n508), .A2(new_n507), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT75), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n506), .A2(G110), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n425), .A2(new_n426), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n511), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n216), .A2(G221), .A3(G234), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT22), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(G137), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n511), .B(new_n520), .C1(new_n515), .C2(new_n516), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n310), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT76), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT25), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n524), .A2(new_n526), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT76), .B1(new_n524), .B2(new_n526), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n502), .B(new_n527), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n522), .A2(new_n523), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n502), .A2(G902), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(KEYINPUT77), .ZN(new_n536));
  INV_X1    g350(.A(new_n348), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT69), .B1(new_n196), .B2(new_n205), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n363), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n354), .A2(new_n357), .A3(new_n428), .A4(new_n355), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n353), .A2(G137), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n356), .A2(G134), .ZN(new_n542));
  OAI21_X1  g356(.A(G131), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n213), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n539), .A2(KEYINPUT30), .A3(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n345), .A2(new_n346), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n547), .A2(new_n363), .B1(new_n544), .B2(new_n213), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT66), .B1(new_n548), .B2(KEYINPUT30), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT66), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT30), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n206), .B1(new_n360), .B2(new_n362), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n544), .A2(new_n213), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n550), .B(new_n551), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n274), .A2(new_n280), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n546), .A2(new_n549), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT70), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n272), .A2(new_n273), .A3(new_n271), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT68), .B1(new_n279), .B2(new_n256), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n274), .A2(new_n280), .A3(KEYINPUT70), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n560), .A2(new_n561), .A3(new_n539), .A4(new_n545), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n412), .A2(G210), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT27), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(KEYINPUT26), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(new_n238), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n556), .A2(new_n562), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT31), .ZN(new_n569));
  INV_X1    g383(.A(new_n567), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT28), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n555), .B1(new_n553), .B2(new_n552), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n571), .B1(new_n562), .B2(new_n572), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n274), .A2(KEYINPUT70), .A3(new_n280), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT70), .B1(new_n274), .B2(new_n280), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n553), .B1(new_n349), .B2(new_n363), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT28), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n570), .B1(new_n573), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT31), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n556), .A2(new_n580), .A3(new_n562), .A4(new_n567), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n569), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G472), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n583), .A3(new_n310), .ZN(new_n584));
  XOR2_X1   g398(.A(KEYINPUT71), .B(KEYINPUT32), .Z(new_n585));
  AND3_X1   g399(.A1(new_n584), .A2(KEYINPUT72), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT72), .B1(new_n584), .B2(new_n585), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n562), .A2(new_n571), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n562), .A2(new_n572), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n589), .B(new_n567), .C1(new_n590), .C2(new_n571), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT29), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n556), .A2(new_n562), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT73), .B1(new_n594), .B2(new_n570), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n594), .A2(KEYINPUT73), .A3(new_n570), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n593), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n539), .A2(new_n545), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n598), .B1(new_n575), .B2(new_n574), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n562), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(KEYINPUT28), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT74), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n571), .B1(new_n599), .B2(new_n562), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT74), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n570), .A2(new_n592), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n602), .A2(new_n589), .A3(new_n605), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n310), .ZN(new_n608));
  OAI21_X1  g422(.A(G472), .B1(new_n597), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT32), .ZN(new_n610));
  OR2_X1    g424(.A1(new_n584), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n536), .B1(new_n588), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n501), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  NAND2_X1  g430(.A1(new_n404), .A2(new_n406), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n318), .A2(new_n497), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  OR3_X1    g433(.A1(new_n479), .A2(new_n480), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n619), .B1(new_n479), .B2(new_n480), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n620), .A2(G478), .A3(new_n310), .A4(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT96), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n481), .A2(new_n482), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n623), .B1(new_n622), .B2(new_n624), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n456), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n618), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n536), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n583), .B1(new_n582), .B2(new_n310), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n584), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n617), .A2(new_n631), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT34), .B(G104), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G6));
  INV_X1    g453(.A(KEYINPUT97), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n449), .A2(new_n640), .A3(new_n451), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n450), .B1(new_n446), .B2(new_n447), .ZN(new_n642));
  INV_X1    g456(.A(new_n447), .ZN(new_n643));
  AOI211_X1 g457(.A(KEYINPUT20), .B(new_n643), .C1(new_n434), .C2(new_n445), .ZN(new_n644));
  OAI21_X1  g458(.A(KEYINPUT97), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n646), .A2(new_n455), .A3(new_n484), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n318), .A2(new_n497), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n617), .A2(new_n636), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT35), .B(G107), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  NAND3_X1  g465(.A1(new_n532), .A2(KEYINPUT25), .A3(new_n310), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n652), .A2(KEYINPUT76), .A3(new_n528), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n527), .A2(new_n502), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n521), .A2(KEYINPUT36), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n517), .B(new_n655), .ZN(new_n656));
  AOI22_X1  g470(.A1(new_n653), .A2(new_n654), .B1(new_n533), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n635), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n501), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT37), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  INV_X1    g475(.A(KEYINPUT98), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n490), .B1(new_n493), .B2(G900), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n646), .A2(new_n455), .A3(new_n484), .A4(new_n663), .ZN(new_n664));
  AOI211_X1 g478(.A(new_n188), .B(new_n664), .C1(new_n312), .C2(new_n317), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n405), .B1(new_n400), .B2(new_n402), .ZN(new_n666));
  INV_X1    g480(.A(new_n402), .ZN(new_n667));
  AOI211_X1 g481(.A(KEYINPUT85), .B(new_n667), .C1(new_n389), .C2(new_n399), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n665), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n656), .A2(new_n533), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n531), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n671), .B1(new_n588), .B2(new_n612), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n662), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n609), .A2(new_n611), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n584), .A2(new_n585), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT72), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n584), .A2(KEYINPUT72), .A3(new_n585), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n657), .B1(new_n674), .B2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n617), .A2(KEYINPUT98), .A3(new_n680), .A4(new_n665), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n673), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  NOR2_X1   g497(.A1(new_n584), .A2(new_n610), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n594), .A2(new_n567), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n685), .B(new_n310), .C1(new_n567), .C2(new_n600), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n684), .B1(G472), .B2(new_n686), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n679), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n312), .A2(new_n317), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT38), .ZN(new_n691));
  AND4_X1   g505(.A1(new_n456), .A2(new_n657), .A3(new_n484), .A4(new_n187), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT40), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT99), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n663), .B(KEYINPUT39), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n617), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n695), .B1(new_n617), .B2(new_n696), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n694), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n617), .A2(new_n696), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT99), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(KEYINPUT40), .A3(new_n697), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n693), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n199), .ZN(G45));
  OAI211_X1 g519(.A(new_n456), .B(new_n663), .C1(new_n625), .C2(new_n626), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n318), .B(new_n707), .C1(new_n666), .C2(new_n668), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n680), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT100), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n197), .ZN(G48));
  NAND2_X1  g526(.A1(new_n375), .A2(new_n387), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n310), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(G469), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n388), .A2(new_n320), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n667), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n614), .A2(new_n631), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  NAND3_X1  g535(.A1(new_n614), .A2(new_n648), .A3(new_n718), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  AND3_X1   g537(.A1(new_n718), .A2(new_n499), .A3(new_n318), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n680), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  NAND3_X1  g540(.A1(new_n318), .A2(new_n456), .A3(new_n484), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n715), .A2(new_n716), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n497), .A3(new_n402), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(G472), .A2(G902), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n605), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n589), .B1(new_n603), .B2(new_n604), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n570), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n569), .A2(new_n581), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n732), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n633), .ZN(new_n738));
  INV_X1    g552(.A(new_n535), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT101), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT101), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n738), .A2(new_n742), .A3(new_n739), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n730), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G122), .ZN(G24));
  INV_X1    g560(.A(KEYINPUT103), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT102), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n748), .B1(new_n738), .B2(new_n671), .ZN(new_n749));
  NOR4_X1   g563(.A1(new_n737), .A2(new_n657), .A3(new_n633), .A4(KEYINPUT102), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n707), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n718), .A2(new_n318), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n747), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n735), .A2(new_n736), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n634), .B(new_n671), .C1(new_n754), .C2(new_n732), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT102), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n738), .A2(new_n748), .A3(new_n671), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n706), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n718), .A2(new_n318), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n759), .A3(KEYINPUT103), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n753), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G125), .ZN(G27));
  NAND3_X1  g576(.A1(new_n312), .A2(new_n317), .A3(new_n187), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT104), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n312), .A2(new_n317), .A3(KEYINPUT104), .A4(new_n187), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n392), .A2(new_n393), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(G469), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n667), .B1(new_n389), .B2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT42), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n706), .A2(new_n770), .ZN(new_n771));
  AND4_X1   g585(.A1(new_n765), .A2(new_n766), .A3(new_n769), .A4(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT105), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n584), .A2(new_n610), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT106), .ZN(new_n775));
  OAI22_X1  g589(.A1(new_n684), .A2(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n584), .A2(KEYINPUT105), .A3(new_n610), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n774), .A2(new_n775), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n779), .A2(new_n609), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n535), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n772), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n765), .A2(new_n766), .A3(new_n769), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n783), .A2(new_n613), .A3(new_n706), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n782), .B1(new_n784), .B2(KEYINPUT42), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G131), .ZN(G33));
  OR3_X1    g600(.A1(new_n783), .A2(new_n613), .A3(new_n664), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G134), .ZN(G36));
  AND2_X1   g602(.A1(new_n765), .A2(new_n766), .ZN(new_n789));
  XOR2_X1   g603(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n790));
  OR3_X1    g604(.A1(new_n627), .A2(new_n456), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n792), .B1(new_n627), .B2(new_n456), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n635), .A3(new_n671), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT44), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n789), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT108), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n767), .A2(KEYINPUT45), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(G469), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT45), .B1(new_n394), .B2(new_n398), .ZN(new_n801));
  OAI22_X1  g615(.A1(new_n800), .A2(new_n801), .B1(new_n320), .B2(new_n310), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT46), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n802), .A2(new_n803), .B1(new_n320), .B2(new_n388), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n804), .B1(new_n803), .B2(new_n802), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n402), .A3(new_n696), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n806), .B1(new_n796), .B2(new_n795), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n798), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G137), .ZN(G39));
  XNOR2_X1  g623(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n805), .A2(new_n402), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n812), .B1(new_n805), .B2(new_n402), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n789), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n674), .A2(new_n679), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n815), .A2(new_n816), .A3(new_n536), .A4(new_n706), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G140), .ZN(G42));
  NOR2_X1   g633(.A1(new_n627), .A2(new_n456), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n717), .A2(KEYINPUT49), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n717), .A2(KEYINPUT49), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n535), .A2(new_n667), .A3(new_n188), .ZN(new_n823));
  AND4_X1   g637(.A1(new_n820), .A2(new_n821), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT38), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n690), .B(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n824), .A2(new_n688), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n707), .B(new_n769), .C1(new_n749), .C2(new_n750), .ZN(new_n829));
  INV_X1    g643(.A(new_n484), .ZN(new_n830));
  AND4_X1   g644(.A1(new_n455), .A2(new_n646), .A3(new_n830), .A4(new_n663), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n831), .B1(new_n666), .B2(new_n668), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n829), .B1(new_n832), .B2(new_n672), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n789), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n785), .A2(new_n834), .A3(new_n787), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n407), .B(new_n499), .C1(new_n614), .C2(new_n658), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n744), .A2(new_n730), .B1(new_n724), .B2(new_n680), .ZN(new_n837));
  INV_X1    g651(.A(new_n618), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n630), .B1(new_n456), .B2(new_n830), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n617), .A2(new_n636), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n614), .B(new_n718), .C1(new_n631), .C2(new_n648), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n836), .A2(new_n837), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n835), .A2(new_n842), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n673), .A2(new_n681), .B1(new_n753), .B2(new_n760), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n769), .A2(new_n657), .A3(new_n663), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n688), .A2(new_n727), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n846), .B1(new_n709), .B2(new_n680), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n844), .A2(KEYINPUT52), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n849), .B1(new_n844), .B2(new_n847), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n843), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT52), .B1(new_n844), .B2(new_n847), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n843), .B(KEYINPUT53), .C1(new_n848), .C2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n828), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT111), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n855), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n847), .A2(new_n682), .A3(new_n761), .ZN(new_n860));
  INV_X1    g674(.A(new_n849), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n844), .A2(KEYINPUT52), .A3(new_n847), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT53), .B1(new_n864), .B2(new_n843), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT54), .B1(new_n859), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT111), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n843), .B1(new_n848), .B2(new_n854), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(new_n852), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n843), .B(KEYINPUT53), .C1(new_n848), .C2(new_n850), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(new_n828), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n490), .B1(new_n791), .B2(new_n793), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n789), .A2(new_n718), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n781), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT48), .Z(new_n876));
  NOR2_X1   g690(.A1(new_n632), .A2(new_n490), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n789), .A2(new_n688), .A3(new_n877), .A4(new_n718), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n630), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n744), .A2(new_n872), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n880), .A2(new_n752), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n879), .A2(new_n488), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n876), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n627), .A2(new_n628), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n878), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n749), .A2(new_n750), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n873), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT51), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT50), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n718), .A2(new_n188), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n691), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT112), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n744), .B(new_n872), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n826), .A2(new_n188), .A3(new_n718), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n895), .A2(KEYINPUT112), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n890), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n880), .B1(new_n895), .B2(KEYINPUT112), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n892), .A2(new_n893), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n898), .A2(KEYINPUT50), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n889), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n728), .A2(new_n667), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n902), .B1(new_n811), .B2(new_n813), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT114), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n880), .A2(new_n815), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT114), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n906), .B(new_n902), .C1(new_n811), .C2(new_n813), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n883), .B1(new_n901), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT113), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n894), .A2(new_n896), .A3(new_n890), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT50), .B1(new_n898), .B2(new_n899), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n903), .A2(new_n905), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n897), .A2(new_n900), .A3(KEYINPUT113), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n913), .A2(new_n914), .A3(new_n888), .A4(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT51), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n909), .A2(new_n918), .ZN(new_n919));
  AND4_X1   g733(.A1(new_n858), .A2(new_n867), .A3(new_n871), .A4(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(G952), .A2(G953), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n827), .B1(new_n920), .B2(new_n921), .ZN(G75));
  NOR2_X1   g736(.A1(new_n216), .A2(G952), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n310), .B1(new_n869), .B2(new_n870), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT56), .B1(new_n925), .B2(G210), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n313), .A2(new_n314), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(new_n218), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT115), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT55), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n924), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n925), .A2(G210), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT56), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n932), .A2(new_n933), .A3(new_n930), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT116), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n926), .A2(KEYINPUT116), .A3(new_n930), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n931), .B1(new_n936), .B2(new_n937), .ZN(G51));
  XNOR2_X1  g752(.A(new_n321), .B(KEYINPUT57), .ZN(new_n939));
  INV_X1    g753(.A(new_n871), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n828), .B1(new_n869), .B2(new_n870), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n713), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n800), .A2(new_n801), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT117), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n925), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n923), .B1(new_n943), .B2(new_n946), .ZN(G54));
  NAND3_X1  g761(.A1(new_n925), .A2(KEYINPUT58), .A3(G475), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n948), .A2(new_n434), .A3(new_n445), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n925), .A2(KEYINPUT58), .A3(G475), .A4(new_n446), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n949), .A2(new_n924), .A3(new_n950), .ZN(G60));
  NAND2_X1  g765(.A1(new_n620), .A2(new_n621), .ZN(new_n952));
  NAND2_X1  g766(.A1(G478), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT59), .Z(new_n954));
  NOR2_X1   g768(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(new_n940), .B2(new_n941), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n924), .ZN(new_n957));
  INV_X1    g771(.A(new_n954), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n871), .B1(new_n856), .B2(new_n857), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n866), .A2(KEYINPUT111), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n957), .B1(new_n961), .B2(new_n952), .ZN(G63));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT60), .Z(new_n964));
  INV_X1    g778(.A(new_n870), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT52), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n860), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n863), .ZN(new_n968));
  AOI21_X1  g782(.A(KEYINPUT53), .B1(new_n968), .B2(new_n843), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n964), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n532), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n923), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n869), .A2(new_n870), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT118), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n973), .A2(new_n974), .A3(new_n656), .A4(new_n964), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n656), .B(new_n964), .C1(new_n965), .C2(new_n969), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(KEYINPUT118), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n972), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT61), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n923), .A2(new_n979), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n970), .A2(KEYINPUT119), .A3(new_n971), .ZN(new_n982));
  AOI21_X1  g796(.A(KEYINPUT119), .B1(new_n970), .B2(new_n971), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n976), .B(new_n981), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n980), .A2(new_n984), .ZN(G66));
  NAND2_X1  g799(.A1(new_n842), .A2(new_n216), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT120), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n216), .B1(new_n495), .B2(G224), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT121), .Z(new_n989));
  NAND2_X1  g803(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n927), .B1(G898), .B2(new_n216), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(G69));
  NAND3_X1  g806(.A1(new_n546), .A2(new_n549), .A3(new_n554), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n440), .A2(new_n441), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n993), .B(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n844), .A2(new_n710), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n704), .A2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT62), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n818), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(new_n996), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n700), .A2(new_n703), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n1000), .B(new_n998), .C1(new_n1001), .C2(new_n693), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(KEYINPUT122), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT122), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n997), .A2(new_n1004), .A3(new_n998), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n999), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n839), .B(KEYINPUT123), .ZN(new_n1007));
  NOR3_X1   g821(.A1(new_n1007), .A2(new_n613), .A3(new_n815), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1008), .A2(new_n697), .A3(new_n702), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n1006), .A2(new_n216), .A3(new_n808), .A4(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n995), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n323), .A2(KEYINPUT124), .A3(G900), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n1013), .B(G953), .C1(KEYINPUT124), .C2(G900), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n995), .A2(new_n1014), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n808), .A2(new_n818), .ZN(new_n1016));
  NOR3_X1   g830(.A1(new_n806), .A2(new_n727), .A3(new_n874), .ZN(new_n1017));
  INV_X1    g831(.A(new_n787), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AND2_X1   g833(.A1(new_n1019), .A2(new_n785), .ZN(new_n1020));
  AND3_X1   g834(.A1(new_n1016), .A2(new_n1000), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1015), .B1(new_n1021), .B2(new_n216), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1012), .A2(new_n1022), .ZN(G72));
  XNOR2_X1  g837(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n583), .A2(new_n310), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1024), .B(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(new_n568), .ZN(new_n1027));
  OR2_X1    g841(.A1(new_n596), .A2(new_n595), .ZN(new_n1028));
  OAI221_X1 g842(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .C1(new_n859), .C2(new_n865), .ZN(new_n1029));
  INV_X1    g843(.A(new_n1026), .ZN(new_n1030));
  INV_X1    g844(.A(new_n842), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1030), .B1(new_n1021), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n570), .A2(new_n556), .A3(new_n562), .ZN(new_n1033));
  OAI211_X1 g847(.A(new_n924), .B(new_n1029), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  AND3_X1   g848(.A1(new_n808), .A2(new_n1031), .A3(new_n1009), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1030), .B1(new_n1006), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g850(.A(KEYINPUT126), .B1(new_n1036), .B2(new_n685), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1038));
  INV_X1    g852(.A(new_n999), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n1038), .A2(new_n1039), .A3(new_n1035), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1040), .A2(new_n1026), .ZN(new_n1041));
  INV_X1    g855(.A(KEYINPUT126), .ZN(new_n1042));
  INV_X1    g856(.A(new_n685), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1034), .B1(new_n1037), .B2(new_n1044), .ZN(G57));
endmodule


