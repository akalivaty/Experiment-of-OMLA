

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X2 U554 ( .A(G2104), .ZN(n527) );
  XNOR2_X2 U555 ( .A(n533), .B(KEYINPUT64), .ZN(G160) );
  NOR2_X1 U556 ( .A1(n696), .A2(n695), .ZN(n705) );
  AND2_X1 U557 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U558 ( .A1(G8), .A2(n661), .ZN(n703) );
  INV_X1 U559 ( .A(n661), .ZN(n642) );
  AND2_X2 U560 ( .A1(n527), .A2(G2105), .ZN(n880) );
  NOR2_X1 U561 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U562 ( .A(KEYINPUT1), .B(n544), .Z(n784) );
  XOR2_X1 U563 ( .A(KEYINPUT74), .B(n602), .Z(n521) );
  NOR2_X1 U564 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U565 ( .A(n606), .B(KEYINPUT15), .ZN(n928) );
  NOR2_X1 U566 ( .A1(G651), .A2(n548), .ZN(n789) );
  NOR2_X1 U567 ( .A1(G651), .A2(G543), .ZN(n788) );
  AND2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n881) );
  NAND2_X1 U569 ( .A1(G113), .A2(n881), .ZN(n524) );
  NOR2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XOR2_X1 U571 ( .A(KEYINPUT17), .B(n522), .Z(n534) );
  NAND2_X1 U572 ( .A1(G137), .A2(n534), .ZN(n523) );
  NAND2_X1 U573 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U574 ( .A(n525), .B(KEYINPUT66), .ZN(n532) );
  NAND2_X1 U575 ( .A1(G125), .A2(n880), .ZN(n526) );
  XOR2_X1 U576 ( .A(KEYINPUT65), .B(n526), .Z(n530) );
  NOR2_X4 U577 ( .A1(G2105), .A2(n527), .ZN(n876) );
  NAND2_X1 U578 ( .A1(G101), .A2(n876), .ZN(n528) );
  XOR2_X1 U579 ( .A(KEYINPUT23), .B(n528), .Z(n529) );
  NAND2_X1 U580 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U581 ( .A1(n532), .A2(n531), .ZN(n533) );
  BUF_X1 U582 ( .A(n534), .Z(n875) );
  NAND2_X1 U583 ( .A1(G138), .A2(n875), .ZN(n536) );
  NAND2_X1 U584 ( .A1(G102), .A2(n876), .ZN(n535) );
  NAND2_X1 U585 ( .A1(n536), .A2(n535), .ZN(n541) );
  NAND2_X1 U586 ( .A1(G126), .A2(n880), .ZN(n538) );
  NAND2_X1 U587 ( .A1(G114), .A2(n881), .ZN(n537) );
  NAND2_X1 U588 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U589 ( .A(KEYINPUT87), .B(n539), .Z(n540) );
  NOR2_X1 U590 ( .A1(n541), .A2(n540), .ZN(G164) );
  NAND2_X1 U591 ( .A1(G91), .A2(n788), .ZN(n543) );
  XOR2_X1 U592 ( .A(KEYINPUT0), .B(G543), .Z(n548) );
  NAND2_X1 U593 ( .A1(G53), .A2(n789), .ZN(n542) );
  NAND2_X1 U594 ( .A1(n543), .A2(n542), .ZN(n547) );
  INV_X1 U595 ( .A(G651), .ZN(n549) );
  NOR2_X1 U596 ( .A1(G543), .A2(n549), .ZN(n544) );
  NAND2_X1 U597 ( .A1(G65), .A2(n784), .ZN(n545) );
  XNOR2_X1 U598 ( .A(KEYINPUT71), .B(n545), .ZN(n546) );
  NOR2_X1 U599 ( .A1(n547), .A2(n546), .ZN(n552) );
  OR2_X1 U600 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X2 U601 ( .A(KEYINPUT67), .B(n550), .ZN(n785) );
  NAND2_X1 U602 ( .A1(n785), .A2(G78), .ZN(n551) );
  NAND2_X1 U603 ( .A1(n552), .A2(n551), .ZN(G299) );
  NAND2_X1 U604 ( .A1(G52), .A2(n789), .ZN(n553) );
  XOR2_X1 U605 ( .A(KEYINPUT68), .B(n553), .Z(n560) );
  NAND2_X1 U606 ( .A1(n788), .A2(G90), .ZN(n554) );
  XNOR2_X1 U607 ( .A(KEYINPUT69), .B(n554), .ZN(n557) );
  NAND2_X1 U608 ( .A1(n785), .A2(G77), .ZN(n555) );
  XOR2_X1 U609 ( .A(KEYINPUT70), .B(n555), .Z(n556) );
  NOR2_X1 U610 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U611 ( .A(n558), .B(KEYINPUT9), .ZN(n559) );
  NOR2_X1 U612 ( .A1(n560), .A2(n559), .ZN(n562) );
  NAND2_X1 U613 ( .A1(n784), .A2(G64), .ZN(n561) );
  NAND2_X1 U614 ( .A1(n562), .A2(n561), .ZN(G301) );
  NAND2_X1 U615 ( .A1(n788), .A2(G89), .ZN(n563) );
  XNOR2_X1 U616 ( .A(n563), .B(KEYINPUT4), .ZN(n565) );
  NAND2_X1 U617 ( .A1(G76), .A2(n785), .ZN(n564) );
  NAND2_X1 U618 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U619 ( .A(n566), .B(KEYINPUT5), .ZN(n572) );
  NAND2_X1 U620 ( .A1(n789), .A2(G51), .ZN(n567) );
  XNOR2_X1 U621 ( .A(n567), .B(KEYINPUT76), .ZN(n569) );
  NAND2_X1 U622 ( .A1(G63), .A2(n784), .ZN(n568) );
  NAND2_X1 U623 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U624 ( .A(KEYINPUT6), .B(n570), .Z(n571) );
  NAND2_X1 U625 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U626 ( .A(n573), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G62), .A2(n784), .ZN(n575) );
  NAND2_X1 U629 ( .A1(G50), .A2(n789), .ZN(n574) );
  NAND2_X1 U630 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U631 ( .A(KEYINPUT83), .B(n576), .ZN(n580) );
  NAND2_X1 U632 ( .A1(G75), .A2(n785), .ZN(n578) );
  NAND2_X1 U633 ( .A1(G88), .A2(n788), .ZN(n577) );
  AND2_X1 U634 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U635 ( .A1(n580), .A2(n579), .ZN(G303) );
  NAND2_X1 U636 ( .A1(G49), .A2(n789), .ZN(n582) );
  NAND2_X1 U637 ( .A1(G74), .A2(G651), .ZN(n581) );
  NAND2_X1 U638 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U639 ( .A1(n784), .A2(n583), .ZN(n585) );
  NAND2_X1 U640 ( .A1(n548), .A2(G87), .ZN(n584) );
  NAND2_X1 U641 ( .A1(n585), .A2(n584), .ZN(G288) );
  NAND2_X1 U642 ( .A1(G73), .A2(n785), .ZN(n586) );
  XNOR2_X1 U643 ( .A(n586), .B(KEYINPUT2), .ZN(n593) );
  NAND2_X1 U644 ( .A1(G61), .A2(n784), .ZN(n588) );
  NAND2_X1 U645 ( .A1(G86), .A2(n788), .ZN(n587) );
  NAND2_X1 U646 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U647 ( .A1(n789), .A2(G48), .ZN(n589) );
  XOR2_X1 U648 ( .A(KEYINPUT82), .B(n589), .Z(n590) );
  NOR2_X1 U649 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U650 ( .A1(n593), .A2(n592), .ZN(G305) );
  AND2_X1 U651 ( .A1(n785), .A2(G72), .ZN(n597) );
  NAND2_X1 U652 ( .A1(G60), .A2(n784), .ZN(n595) );
  NAND2_X1 U653 ( .A1(G47), .A2(n789), .ZN(n594) );
  NAND2_X1 U654 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U655 ( .A1(n597), .A2(n596), .ZN(n599) );
  NAND2_X1 U656 ( .A1(n788), .A2(G85), .ZN(n598) );
  NAND2_X1 U657 ( .A1(n599), .A2(n598), .ZN(G290) );
  NAND2_X1 U658 ( .A1(G54), .A2(n789), .ZN(n605) );
  NAND2_X1 U659 ( .A1(G66), .A2(n784), .ZN(n601) );
  NAND2_X1 U660 ( .A1(G92), .A2(n788), .ZN(n600) );
  NAND2_X1 U661 ( .A1(n601), .A2(n600), .ZN(n603) );
  NAND2_X1 U662 ( .A1(n785), .A2(G79), .ZN(n602) );
  NOR2_X1 U663 ( .A1(n603), .A2(n521), .ZN(n604) );
  NAND2_X1 U664 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U665 ( .A1(G56), .A2(n784), .ZN(n607) );
  XOR2_X1 U666 ( .A(KEYINPUT14), .B(n607), .Z(n614) );
  NAND2_X1 U667 ( .A1(n788), .A2(G81), .ZN(n608) );
  XOR2_X1 U668 ( .A(KEYINPUT12), .B(n608), .Z(n611) );
  NAND2_X1 U669 ( .A1(n785), .A2(G68), .ZN(n609) );
  XOR2_X1 U670 ( .A(KEYINPUT72), .B(n609), .Z(n610) );
  NOR2_X1 U671 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U672 ( .A(n612), .B(KEYINPUT13), .ZN(n613) );
  NOR2_X1 U673 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U674 ( .A1(n789), .A2(G43), .ZN(n615) );
  NAND2_X1 U675 ( .A1(n616), .A2(n615), .ZN(n927) );
  NOR2_X1 U676 ( .A1(G164), .A2(G1384), .ZN(n707) );
  NAND2_X1 U677 ( .A1(G40), .A2(G160), .ZN(n706) );
  INV_X1 U678 ( .A(n706), .ZN(n617) );
  NAND2_X1 U679 ( .A1(n707), .A2(n617), .ZN(n661) );
  NAND2_X1 U680 ( .A1(n642), .A2(G1996), .ZN(n619) );
  XOR2_X1 U681 ( .A(KEYINPUT26), .B(KEYINPUT93), .Z(n618) );
  XNOR2_X1 U682 ( .A(n619), .B(n618), .ZN(n621) );
  NAND2_X1 U683 ( .A1(n661), .A2(G1341), .ZN(n620) );
  NAND2_X1 U684 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U685 ( .A1(n927), .A2(n622), .ZN(n628) );
  NAND2_X1 U686 ( .A1(n928), .A2(n628), .ZN(n627) );
  AND2_X1 U687 ( .A1(n642), .A2(G2067), .ZN(n623) );
  XOR2_X1 U688 ( .A(n623), .B(KEYINPUT94), .Z(n625) );
  NAND2_X1 U689 ( .A1(n661), .A2(G1348), .ZN(n624) );
  NAND2_X1 U690 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U691 ( .A1(n627), .A2(n626), .ZN(n630) );
  OR2_X1 U692 ( .A1(n928), .A2(n628), .ZN(n629) );
  NAND2_X1 U693 ( .A1(n630), .A2(n629), .ZN(n636) );
  INV_X1 U694 ( .A(G299), .ZN(n797) );
  NAND2_X1 U695 ( .A1(n642), .A2(G2072), .ZN(n631) );
  XNOR2_X1 U696 ( .A(KEYINPUT27), .B(n631), .ZN(n634) );
  NAND2_X1 U697 ( .A1(G1956), .A2(n661), .ZN(n632) );
  XOR2_X1 U698 ( .A(KEYINPUT92), .B(n632), .Z(n633) );
  NOR2_X1 U699 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U700 ( .A1(n797), .A2(n637), .ZN(n635) );
  NAND2_X1 U701 ( .A1(n636), .A2(n635), .ZN(n640) );
  NOR2_X1 U702 ( .A1(n797), .A2(n637), .ZN(n638) );
  XOR2_X1 U703 ( .A(n638), .B(KEYINPUT28), .Z(n639) );
  NAND2_X1 U704 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U705 ( .A(n641), .B(KEYINPUT29), .ZN(n646) );
  XOR2_X1 U706 ( .A(G2078), .B(KEYINPUT25), .Z(n972) );
  NOR2_X1 U707 ( .A1(n972), .A2(n661), .ZN(n644) );
  NOR2_X1 U708 ( .A1(n642), .A2(G1961), .ZN(n643) );
  NOR2_X1 U709 ( .A1(n644), .A2(n643), .ZN(n654) );
  NOR2_X1 U710 ( .A1(G301), .A2(n654), .ZN(n645) );
  XNOR2_X1 U711 ( .A(n647), .B(KEYINPUT95), .ZN(n660) );
  NOR2_X1 U712 ( .A1(G1966), .A2(n703), .ZN(n673) );
  NOR2_X1 U713 ( .A1(G2084), .A2(n661), .ZN(n670) );
  INV_X1 U714 ( .A(G8), .ZN(n648) );
  OR2_X1 U715 ( .A1(n670), .A2(n648), .ZN(n649) );
  OR2_X1 U716 ( .A1(n673), .A2(n649), .ZN(n650) );
  XNOR2_X1 U717 ( .A(n650), .B(KEYINPUT97), .ZN(n652) );
  XOR2_X1 U718 ( .A(KEYINPUT30), .B(KEYINPUT96), .Z(n651) );
  XNOR2_X1 U719 ( .A(n652), .B(n651), .ZN(n653) );
  NOR2_X1 U720 ( .A1(n653), .A2(G168), .ZN(n656) );
  AND2_X1 U721 ( .A1(G301), .A2(n654), .ZN(n655) );
  XOR2_X1 U722 ( .A(n657), .B(KEYINPUT31), .Z(n658) );
  XNOR2_X1 U723 ( .A(n658), .B(KEYINPUT98), .ZN(n659) );
  NAND2_X1 U724 ( .A1(n660), .A2(n659), .ZN(n671) );
  NAND2_X1 U725 ( .A1(n671), .A2(G286), .ZN(n668) );
  NOR2_X1 U726 ( .A1(G1971), .A2(n703), .ZN(n663) );
  NOR2_X1 U727 ( .A1(G2090), .A2(n661), .ZN(n662) );
  NOR2_X1 U728 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U729 ( .A(KEYINPUT99), .B(n664), .Z(n665) );
  NAND2_X1 U730 ( .A1(n665), .A2(G303), .ZN(n666) );
  OR2_X1 U731 ( .A1(n648), .A2(n666), .ZN(n667) );
  XNOR2_X1 U732 ( .A(n669), .B(KEYINPUT32), .ZN(n697) );
  NAND2_X1 U733 ( .A1(G8), .A2(n670), .ZN(n675) );
  INV_X1 U734 ( .A(n671), .ZN(n672) );
  NOR2_X1 U735 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U736 ( .A1(n675), .A2(n674), .ZN(n698) );
  NAND2_X1 U737 ( .A1(G288), .A2(G1976), .ZN(n676) );
  XNOR2_X1 U738 ( .A(n676), .B(KEYINPUT100), .ZN(n918) );
  INV_X1 U739 ( .A(n918), .ZN(n677) );
  NOR2_X1 U740 ( .A1(n677), .A2(n703), .ZN(n678) );
  NOR2_X1 U741 ( .A1(KEYINPUT33), .A2(n678), .ZN(n681) );
  NOR2_X1 U742 ( .A1(G1976), .A2(G288), .ZN(n916) );
  NAND2_X1 U743 ( .A1(n916), .A2(KEYINPUT33), .ZN(n679) );
  NOR2_X1 U744 ( .A1(n679), .A2(n703), .ZN(n680) );
  NOR2_X1 U745 ( .A1(n681), .A2(n680), .ZN(n683) );
  AND2_X1 U746 ( .A1(n698), .A2(n683), .ZN(n682) );
  NAND2_X1 U747 ( .A1(n697), .A2(n682), .ZN(n690) );
  INV_X1 U748 ( .A(n683), .ZN(n688) );
  NOR2_X1 U749 ( .A1(G1971), .A2(G303), .ZN(n684) );
  NOR2_X1 U750 ( .A1(n916), .A2(n684), .ZN(n686) );
  INV_X1 U751 ( .A(KEYINPUT33), .ZN(n685) );
  AND2_X1 U752 ( .A1(n686), .A2(n685), .ZN(n687) );
  OR2_X1 U753 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U754 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U755 ( .A(G1981), .B(G305), .Z(n913) );
  NAND2_X1 U756 ( .A1(n691), .A2(n913), .ZN(n692) );
  XNOR2_X1 U757 ( .A(n692), .B(KEYINPUT101), .ZN(n696) );
  NOR2_X1 U758 ( .A1(G1981), .A2(G305), .ZN(n693) );
  XOR2_X1 U759 ( .A(n693), .B(KEYINPUT24), .Z(n694) );
  NOR2_X1 U760 ( .A1(n703), .A2(n694), .ZN(n695) );
  NAND2_X1 U761 ( .A1(n698), .A2(n697), .ZN(n701) );
  NOR2_X1 U762 ( .A1(G2090), .A2(G303), .ZN(n699) );
  NAND2_X1 U763 ( .A1(G8), .A2(n699), .ZN(n700) );
  NAND2_X1 U764 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U765 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U766 ( .A1(n705), .A2(n704), .ZN(n739) );
  NOR2_X1 U767 ( .A1(n707), .A2(n706), .ZN(n752) );
  NAND2_X1 U768 ( .A1(G129), .A2(n880), .ZN(n709) );
  NAND2_X1 U769 ( .A1(G117), .A2(n881), .ZN(n708) );
  NAND2_X1 U770 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U771 ( .A1(n876), .A2(G105), .ZN(n710) );
  XOR2_X1 U772 ( .A(KEYINPUT38), .B(n710), .Z(n711) );
  NOR2_X1 U773 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U774 ( .A(n713), .B(KEYINPUT90), .ZN(n715) );
  NAND2_X1 U775 ( .A1(G141), .A2(n875), .ZN(n714) );
  NAND2_X1 U776 ( .A1(n715), .A2(n714), .ZN(n872) );
  NAND2_X1 U777 ( .A1(n872), .A2(G1996), .ZN(n724) );
  NAND2_X1 U778 ( .A1(G119), .A2(n880), .ZN(n717) );
  NAND2_X1 U779 ( .A1(G107), .A2(n881), .ZN(n716) );
  NAND2_X1 U780 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U781 ( .A(KEYINPUT89), .B(n718), .ZN(n722) );
  NAND2_X1 U782 ( .A1(G131), .A2(n875), .ZN(n720) );
  NAND2_X1 U783 ( .A1(G95), .A2(n876), .ZN(n719) );
  AND2_X1 U784 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U785 ( .A1(n722), .A2(n721), .ZN(n859) );
  NAND2_X1 U786 ( .A1(G1991), .A2(n859), .ZN(n723) );
  NAND2_X1 U787 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U788 ( .A(n725), .B(KEYINPUT91), .ZN(n1003) );
  NAND2_X1 U789 ( .A1(G140), .A2(n875), .ZN(n727) );
  NAND2_X1 U790 ( .A1(G104), .A2(n876), .ZN(n726) );
  NAND2_X1 U791 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U792 ( .A(KEYINPUT34), .B(n728), .ZN(n733) );
  NAND2_X1 U793 ( .A1(G128), .A2(n880), .ZN(n730) );
  NAND2_X1 U794 ( .A1(G116), .A2(n881), .ZN(n729) );
  NAND2_X1 U795 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U796 ( .A(n731), .B(KEYINPUT35), .Z(n732) );
  NOR2_X1 U797 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U798 ( .A(KEYINPUT36), .B(n734), .Z(n735) );
  XOR2_X1 U799 ( .A(KEYINPUT88), .B(n735), .Z(n890) );
  XNOR2_X1 U800 ( .A(G2067), .B(KEYINPUT37), .ZN(n749) );
  NOR2_X1 U801 ( .A1(n890), .A2(n749), .ZN(n747) );
  XNOR2_X1 U802 ( .A(G1986), .B(G290), .ZN(n923) );
  NOR2_X1 U803 ( .A1(n747), .A2(n923), .ZN(n736) );
  NAND2_X1 U804 ( .A1(n1003), .A2(n736), .ZN(n737) );
  NAND2_X1 U805 ( .A1(n752), .A2(n737), .ZN(n738) );
  NAND2_X1 U806 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U807 ( .A(n740), .B(KEYINPUT102), .ZN(n755) );
  NOR2_X1 U808 ( .A1(G1996), .A2(n872), .ZN(n997) );
  INV_X1 U809 ( .A(n1003), .ZN(n744) );
  NOR2_X1 U810 ( .A1(G1991), .A2(n859), .ZN(n988) );
  NOR2_X1 U811 ( .A1(G1986), .A2(G290), .ZN(n741) );
  NOR2_X1 U812 ( .A1(n988), .A2(n741), .ZN(n742) );
  XOR2_X1 U813 ( .A(KEYINPUT103), .B(n742), .Z(n743) );
  NOR2_X1 U814 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U815 ( .A1(n997), .A2(n745), .ZN(n746) );
  XNOR2_X1 U816 ( .A(n746), .B(KEYINPUT39), .ZN(n748) );
  INV_X1 U817 ( .A(n747), .ZN(n993) );
  NAND2_X1 U818 ( .A1(n748), .A2(n993), .ZN(n750) );
  NAND2_X1 U819 ( .A1(n890), .A2(n749), .ZN(n1002) );
  NAND2_X1 U820 ( .A1(n750), .A2(n1002), .ZN(n751) );
  XNOR2_X1 U821 ( .A(KEYINPUT104), .B(n751), .ZN(n753) );
  NAND2_X1 U822 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U823 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U824 ( .A(n756), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U825 ( .A(G301), .ZN(G171) );
  AND2_X1 U826 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U827 ( .A(G132), .ZN(G219) );
  INV_X1 U828 ( .A(G82), .ZN(G220) );
  INV_X1 U829 ( .A(G57), .ZN(G237) );
  NAND2_X1 U830 ( .A1(G7), .A2(G661), .ZN(n757) );
  XNOR2_X1 U831 ( .A(n757), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U832 ( .A(G223), .ZN(n823) );
  NAND2_X1 U833 ( .A1(n823), .A2(G567), .ZN(n758) );
  XOR2_X1 U834 ( .A(KEYINPUT11), .B(n758), .Z(G234) );
  XNOR2_X1 U835 ( .A(G860), .B(KEYINPUT73), .ZN(n766) );
  OR2_X1 U836 ( .A1(n927), .A2(n766), .ZN(G153) );
  NAND2_X1 U837 ( .A1(G868), .A2(G171), .ZN(n760) );
  INV_X1 U838 ( .A(G868), .ZN(n806) );
  NAND2_X1 U839 ( .A1(n928), .A2(n806), .ZN(n759) );
  NAND2_X1 U840 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U841 ( .A(n761), .B(KEYINPUT75), .ZN(G284) );
  XNOR2_X1 U842 ( .A(KEYINPUT77), .B(G868), .ZN(n762) );
  NOR2_X1 U843 ( .A1(G286), .A2(n762), .ZN(n764) );
  NOR2_X1 U844 ( .A1(G868), .A2(G299), .ZN(n763) );
  NOR2_X1 U845 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U846 ( .A(KEYINPUT78), .B(n765), .ZN(G297) );
  NAND2_X1 U847 ( .A1(n766), .A2(G559), .ZN(n767) );
  NAND2_X1 U848 ( .A1(n767), .A2(n928), .ZN(n768) );
  XNOR2_X1 U849 ( .A(n768), .B(KEYINPUT16), .ZN(n769) );
  XOR2_X1 U850 ( .A(KEYINPUT79), .B(n769), .Z(G148) );
  NOR2_X1 U851 ( .A1(G868), .A2(n927), .ZN(n772) );
  NAND2_X1 U852 ( .A1(G868), .A2(n928), .ZN(n770) );
  NOR2_X1 U853 ( .A1(G559), .A2(n770), .ZN(n771) );
  NOR2_X1 U854 ( .A1(n772), .A2(n771), .ZN(G282) );
  XNOR2_X1 U855 ( .A(G2100), .B(KEYINPUT81), .ZN(n782) );
  NAND2_X1 U856 ( .A1(G123), .A2(n880), .ZN(n773) );
  XNOR2_X1 U857 ( .A(n773), .B(KEYINPUT18), .ZN(n774) );
  XNOR2_X1 U858 ( .A(n774), .B(KEYINPUT80), .ZN(n776) );
  NAND2_X1 U859 ( .A1(G111), .A2(n881), .ZN(n775) );
  NAND2_X1 U860 ( .A1(n776), .A2(n775), .ZN(n780) );
  NAND2_X1 U861 ( .A1(G135), .A2(n875), .ZN(n778) );
  NAND2_X1 U862 ( .A1(G99), .A2(n876), .ZN(n777) );
  NAND2_X1 U863 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U864 ( .A1(n780), .A2(n779), .ZN(n987) );
  XNOR2_X1 U865 ( .A(n987), .B(G2096), .ZN(n781) );
  NAND2_X1 U866 ( .A1(n782), .A2(n781), .ZN(G156) );
  NAND2_X1 U867 ( .A1(n928), .A2(G559), .ZN(n803) );
  XNOR2_X1 U868 ( .A(n927), .B(n803), .ZN(n783) );
  NOR2_X1 U869 ( .A1(n783), .A2(G860), .ZN(n794) );
  NAND2_X1 U870 ( .A1(G67), .A2(n784), .ZN(n787) );
  NAND2_X1 U871 ( .A1(G80), .A2(n785), .ZN(n786) );
  NAND2_X1 U872 ( .A1(n787), .A2(n786), .ZN(n793) );
  NAND2_X1 U873 ( .A1(G93), .A2(n788), .ZN(n791) );
  NAND2_X1 U874 ( .A1(G55), .A2(n789), .ZN(n790) );
  NAND2_X1 U875 ( .A1(n791), .A2(n790), .ZN(n792) );
  OR2_X1 U876 ( .A1(n793), .A2(n792), .ZN(n805) );
  XOR2_X1 U877 ( .A(n794), .B(n805), .Z(G145) );
  INV_X1 U878 ( .A(G303), .ZN(G166) );
  XOR2_X1 U879 ( .A(KEYINPUT84), .B(KEYINPUT19), .Z(n795) );
  XNOR2_X1 U880 ( .A(G288), .B(n795), .ZN(n796) );
  XNOR2_X1 U881 ( .A(G305), .B(n796), .ZN(n799) );
  XNOR2_X1 U882 ( .A(n797), .B(G166), .ZN(n798) );
  XNOR2_X1 U883 ( .A(n799), .B(n798), .ZN(n800) );
  XNOR2_X1 U884 ( .A(n805), .B(n800), .ZN(n801) );
  XNOR2_X1 U885 ( .A(G290), .B(n801), .ZN(n802) );
  XNOR2_X1 U886 ( .A(n802), .B(n927), .ZN(n894) );
  XNOR2_X1 U887 ( .A(n803), .B(n894), .ZN(n804) );
  NAND2_X1 U888 ( .A1(n804), .A2(G868), .ZN(n808) );
  NAND2_X1 U889 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U890 ( .A1(n808), .A2(n807), .ZN(G295) );
  NAND2_X1 U891 ( .A1(G2084), .A2(G2078), .ZN(n809) );
  XOR2_X1 U892 ( .A(KEYINPUT20), .B(n809), .Z(n810) );
  NAND2_X1 U893 ( .A1(G2090), .A2(n810), .ZN(n812) );
  XOR2_X1 U894 ( .A(KEYINPUT85), .B(KEYINPUT21), .Z(n811) );
  XNOR2_X1 U895 ( .A(n812), .B(n811), .ZN(n813) );
  NAND2_X1 U896 ( .A1(G2072), .A2(n813), .ZN(G158) );
  XNOR2_X1 U897 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U898 ( .A1(G69), .A2(G120), .ZN(n814) );
  NOR2_X1 U899 ( .A1(G237), .A2(n814), .ZN(n815) );
  NAND2_X1 U900 ( .A1(G108), .A2(n815), .ZN(n829) );
  NAND2_X1 U901 ( .A1(n829), .A2(G567), .ZN(n821) );
  NOR2_X1 U902 ( .A1(G220), .A2(G219), .ZN(n816) );
  XOR2_X1 U903 ( .A(KEYINPUT22), .B(n816), .Z(n817) );
  NOR2_X1 U904 ( .A1(G218), .A2(n817), .ZN(n818) );
  NAND2_X1 U905 ( .A1(G96), .A2(n818), .ZN(n828) );
  NAND2_X1 U906 ( .A1(G2106), .A2(n828), .ZN(n819) );
  XNOR2_X1 U907 ( .A(KEYINPUT86), .B(n819), .ZN(n820) );
  NAND2_X1 U908 ( .A1(n821), .A2(n820), .ZN(n830) );
  NAND2_X1 U909 ( .A1(G483), .A2(G661), .ZN(n822) );
  NOR2_X1 U910 ( .A1(n830), .A2(n822), .ZN(n827) );
  NAND2_X1 U911 ( .A1(n827), .A2(G36), .ZN(G176) );
  NAND2_X1 U912 ( .A1(G2106), .A2(n823), .ZN(G217) );
  NAND2_X1 U913 ( .A1(G15), .A2(G2), .ZN(n824) );
  XNOR2_X1 U914 ( .A(KEYINPUT105), .B(n824), .ZN(n825) );
  NAND2_X1 U915 ( .A1(n825), .A2(G661), .ZN(G259) );
  NAND2_X1 U916 ( .A1(G3), .A2(G1), .ZN(n826) );
  NAND2_X1 U917 ( .A1(n827), .A2(n826), .ZN(G188) );
  INV_X1 U919 ( .A(G120), .ZN(G236) );
  INV_X1 U920 ( .A(G96), .ZN(G221) );
  INV_X1 U921 ( .A(G69), .ZN(G235) );
  NOR2_X1 U922 ( .A1(n829), .A2(n828), .ZN(G325) );
  INV_X1 U923 ( .A(G325), .ZN(G261) );
  INV_X1 U924 ( .A(n830), .ZN(G319) );
  XOR2_X1 U925 ( .A(G2100), .B(G2678), .Z(n832) );
  XNOR2_X1 U926 ( .A(G2090), .B(KEYINPUT43), .ZN(n831) );
  XNOR2_X1 U927 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U928 ( .A(n833), .B(KEYINPUT42), .Z(n835) );
  XNOR2_X1 U929 ( .A(G2067), .B(G2072), .ZN(n834) );
  XNOR2_X1 U930 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U931 ( .A(KEYINPUT106), .B(G2096), .Z(n837) );
  XNOR2_X1 U932 ( .A(G2084), .B(G2078), .ZN(n836) );
  XNOR2_X1 U933 ( .A(n837), .B(n836), .ZN(n838) );
  XNOR2_X1 U934 ( .A(n839), .B(n838), .ZN(G227) );
  XOR2_X1 U935 ( .A(G1976), .B(G1956), .Z(n841) );
  XNOR2_X1 U936 ( .A(G1966), .B(G1961), .ZN(n840) );
  XNOR2_X1 U937 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U938 ( .A(G1971), .B(G1986), .Z(n843) );
  XNOR2_X1 U939 ( .A(G1996), .B(G1991), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U941 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U942 ( .A(KEYINPUT107), .B(G2474), .ZN(n846) );
  XNOR2_X1 U943 ( .A(n847), .B(n846), .ZN(n849) );
  XOR2_X1 U944 ( .A(G1981), .B(KEYINPUT41), .Z(n848) );
  XNOR2_X1 U945 ( .A(n849), .B(n848), .ZN(G229) );
  NAND2_X1 U946 ( .A1(n880), .A2(G124), .ZN(n850) );
  XNOR2_X1 U947 ( .A(n850), .B(KEYINPUT44), .ZN(n852) );
  NAND2_X1 U948 ( .A1(G112), .A2(n881), .ZN(n851) );
  NAND2_X1 U949 ( .A1(n852), .A2(n851), .ZN(n856) );
  NAND2_X1 U950 ( .A1(G136), .A2(n875), .ZN(n854) );
  NAND2_X1 U951 ( .A1(G100), .A2(n876), .ZN(n853) );
  NAND2_X1 U952 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U953 ( .A1(n856), .A2(n855), .ZN(G162) );
  XOR2_X1 U954 ( .A(KEYINPUT48), .B(KEYINPUT112), .Z(n858) );
  XNOR2_X1 U955 ( .A(KEYINPUT46), .B(KEYINPUT111), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(n862) );
  XNOR2_X1 U957 ( .A(n987), .B(G160), .ZN(n860) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U959 ( .A(n862), .B(n861), .ZN(n874) );
  NAND2_X1 U960 ( .A1(n880), .A2(G127), .ZN(n863) );
  XNOR2_X1 U961 ( .A(n863), .B(KEYINPUT110), .ZN(n865) );
  NAND2_X1 U962 ( .A1(G115), .A2(n881), .ZN(n864) );
  NAND2_X1 U963 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U964 ( .A(n866), .B(KEYINPUT47), .ZN(n868) );
  NAND2_X1 U965 ( .A1(G103), .A2(n876), .ZN(n867) );
  NAND2_X1 U966 ( .A1(n868), .A2(n867), .ZN(n871) );
  NAND2_X1 U967 ( .A1(G139), .A2(n875), .ZN(n869) );
  XNOR2_X1 U968 ( .A(KEYINPUT109), .B(n869), .ZN(n870) );
  NOR2_X1 U969 ( .A1(n871), .A2(n870), .ZN(n1007) );
  XNOR2_X1 U970 ( .A(n872), .B(n1007), .ZN(n873) );
  XNOR2_X1 U971 ( .A(n874), .B(n873), .ZN(n889) );
  NAND2_X1 U972 ( .A1(G142), .A2(n875), .ZN(n878) );
  NAND2_X1 U973 ( .A1(G106), .A2(n876), .ZN(n877) );
  NAND2_X1 U974 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U975 ( .A(n879), .B(KEYINPUT45), .ZN(n886) );
  NAND2_X1 U976 ( .A1(G130), .A2(n880), .ZN(n883) );
  NAND2_X1 U977 ( .A1(G118), .A2(n881), .ZN(n882) );
  NAND2_X1 U978 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U979 ( .A(KEYINPUT108), .B(n884), .Z(n885) );
  NAND2_X1 U980 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U981 ( .A(n887), .B(G162), .ZN(n888) );
  XOR2_X1 U982 ( .A(n889), .B(n888), .Z(n892) );
  XNOR2_X1 U983 ( .A(G164), .B(n890), .ZN(n891) );
  XNOR2_X1 U984 ( .A(n892), .B(n891), .ZN(n893) );
  NOR2_X1 U985 ( .A1(G37), .A2(n893), .ZN(G395) );
  XOR2_X1 U986 ( .A(n894), .B(G286), .Z(n896) );
  XNOR2_X1 U987 ( .A(G171), .B(n928), .ZN(n895) );
  XNOR2_X1 U988 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U989 ( .A1(G37), .A2(n897), .ZN(G397) );
  XOR2_X1 U990 ( .A(G2451), .B(G2430), .Z(n899) );
  XNOR2_X1 U991 ( .A(G2438), .B(G2443), .ZN(n898) );
  XNOR2_X1 U992 ( .A(n899), .B(n898), .ZN(n905) );
  XOR2_X1 U993 ( .A(G2435), .B(G2454), .Z(n901) );
  XNOR2_X1 U994 ( .A(G1341), .B(G1348), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n903) );
  XOR2_X1 U996 ( .A(G2446), .B(G2427), .Z(n902) );
  XNOR2_X1 U997 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U998 ( .A(n905), .B(n904), .Z(n906) );
  NAND2_X1 U999 ( .A1(G14), .A2(n906), .ZN(n912) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n912), .ZN(n909) );
  NOR2_X1 U1001 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(KEYINPUT49), .B(n907), .ZN(n908) );
  NOR2_X1 U1003 ( .A1(n909), .A2(n908), .ZN(n911) );
  NOR2_X1 U1004 ( .A1(G395), .A2(G397), .ZN(n910) );
  NAND2_X1 U1005 ( .A1(n911), .A2(n910), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(G108), .ZN(G238) );
  INV_X1 U1008 ( .A(n912), .ZN(G401) );
  XNOR2_X1 U1009 ( .A(G1966), .B(G168), .ZN(n914) );
  NAND2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n915), .B(KEYINPUT57), .ZN(n936) );
  INV_X1 U1012 ( .A(n916), .ZN(n917) );
  NAND2_X1 U1013 ( .A1(n918), .A2(n917), .ZN(n920) );
  XNOR2_X1 U1014 ( .A(G1956), .B(G299), .ZN(n919) );
  NOR2_X1 U1015 ( .A1(n920), .A2(n919), .ZN(n925) );
  XNOR2_X1 U1016 ( .A(G166), .B(G1971), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(n921), .B(KEYINPUT121), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1019 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1020 ( .A(KEYINPUT122), .B(n926), .ZN(n934) );
  XNOR2_X1 U1021 ( .A(G171), .B(G1961), .ZN(n932) );
  XNOR2_X1 U1022 ( .A(G1341), .B(n927), .ZN(n930) );
  XOR2_X1 U1023 ( .A(G1348), .B(n928), .Z(n929) );
  NOR2_X1 U1024 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1025 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1026 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1027 ( .A1(n936), .A2(n935), .ZN(n939) );
  XNOR2_X1 U1028 ( .A(G16), .B(KEYINPUT120), .ZN(n937) );
  XNOR2_X1 U1029 ( .A(n937), .B(KEYINPUT56), .ZN(n938) );
  NAND2_X1 U1030 ( .A1(n939), .A2(n938), .ZN(n1021) );
  XNOR2_X1 U1031 ( .A(G1971), .B(G22), .ZN(n941) );
  XNOR2_X1 U1032 ( .A(G1976), .B(G23), .ZN(n940) );
  NOR2_X1 U1033 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1034 ( .A(KEYINPUT126), .B(n942), .ZN(n945) );
  XNOR2_X1 U1035 ( .A(G1986), .B(KEYINPUT127), .ZN(n943) );
  XNOR2_X1 U1036 ( .A(n943), .B(G24), .ZN(n944) );
  NAND2_X1 U1037 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1038 ( .A(n946), .B(KEYINPUT58), .ZN(n963) );
  XNOR2_X1 U1039 ( .A(KEYINPUT123), .B(G1956), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(n947), .B(G20), .ZN(n953) );
  XNOR2_X1 U1041 ( .A(KEYINPUT59), .B(G4), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(n948), .B(KEYINPUT125), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(G1348), .B(n949), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(G1981), .B(G6), .ZN(n950) );
  NOR2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n956) );
  XNOR2_X1 U1047 ( .A(KEYINPUT124), .B(G1341), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(G19), .B(n954), .ZN(n955) );
  NOR2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(KEYINPUT60), .B(n957), .ZN(n961) );
  XNOR2_X1 U1051 ( .A(G1966), .B(G21), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(G5), .B(G1961), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(KEYINPUT61), .B(n964), .ZN(n966) );
  INV_X1 U1057 ( .A(G16), .ZN(n965) );
  NAND2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1059 ( .A1(n967), .A2(G11), .ZN(n1019) );
  XNOR2_X1 U1060 ( .A(G2084), .B(G34), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(n968), .B(KEYINPUT54), .ZN(n984) );
  XNOR2_X1 U1062 ( .A(G2090), .B(G35), .ZN(n981) );
  XOR2_X1 U1063 ( .A(G1991), .B(G25), .Z(n969) );
  NAND2_X1 U1064 ( .A1(n969), .A2(G28), .ZN(n978) );
  XNOR2_X1 U1065 ( .A(G1996), .B(G32), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(G33), .B(G2072), .ZN(n970) );
  NOR2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n976) );
  XNOR2_X1 U1068 ( .A(G2067), .B(G26), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(G27), .B(n972), .ZN(n973) );
  NOR2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(KEYINPUT53), .B(n979), .ZN(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(n982), .B(KEYINPUT119), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1077 ( .A1(G29), .A2(n985), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(n986), .B(KEYINPUT55), .ZN(n1017) );
  XNOR2_X1 U1079 ( .A(KEYINPUT52), .B(KEYINPUT118), .ZN(n1014) );
  XOR2_X1 U1080 ( .A(G160), .B(G2084), .Z(n991) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(KEYINPUT113), .B(n989), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1084 ( .A(KEYINPUT114), .B(n992), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1086 ( .A(n995), .B(KEYINPUT115), .ZN(n1001) );
  XOR2_X1 U1087 ( .A(G2090), .B(G162), .Z(n996) );
  XNOR2_X1 U1088 ( .A(KEYINPUT116), .B(n996), .ZN(n998) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1090 ( .A(KEYINPUT51), .B(n999), .Z(n1000) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1005) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1094 ( .A(KEYINPUT117), .B(n1006), .Z(n1012) );
  XOR2_X1 U1095 ( .A(G2072), .B(n1007), .Z(n1009) );
  XOR2_X1 U1096 ( .A(G164), .B(G2078), .Z(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(KEYINPUT50), .B(n1010), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(n1014), .B(n1013), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(G29), .A2(n1015), .ZN(n1016) );
  NAND2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1103 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1104 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1022), .Z(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

