//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 1 0 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  OR3_X1    g002(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT27), .ZN(new_n210));
  INV_X1    g009(.A(G183gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT68), .ZN(new_n213));
  NAND2_X1  g012(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n214));
  AND3_X1   g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n213), .B1(new_n212), .B2(new_n214), .ZN(new_n216));
  OAI211_X1 g015(.A(KEYINPUT28), .B(new_n209), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT27), .B1(new_n218), .B2(new_n211), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n210), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n209), .A3(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI211_X1 g022(.A(new_n203), .B(new_n208), .C1(new_n217), .C2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT25), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(KEYINPUT65), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n209), .ZN(new_n228));
  NAND3_X1  g027(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n225), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  OR3_X1    g031(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n233), .A2(new_n234), .B1(G169gat), .B2(G176gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(new_n230), .B2(new_n226), .ZN(new_n237));
  INV_X1    g036(.A(new_n226), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n238), .A2(new_n228), .A3(KEYINPUT64), .A4(new_n229), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n235), .A3(new_n239), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n232), .A2(new_n235), .B1(new_n240), .B2(new_n225), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT73), .B1(new_n224), .B2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n203), .B1(new_n217), .B2(new_n223), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n207), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n232), .A2(new_n235), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n240), .A2(new_n225), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT73), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n244), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(G226gat), .A2(G233gat), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n251), .A2(KEYINPUT29), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n242), .A2(new_n249), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n243), .A2(new_n254), .A3(new_n207), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n254), .B1(new_n243), .B2(new_n207), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n247), .B(new_n251), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G218gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT71), .B(KEYINPUT22), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT72), .B(G218gat), .ZN(new_n261));
  INV_X1    g060(.A(G211gat), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G197gat), .B(G204gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n259), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n267), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n269), .A2(G218gat), .A3(new_n265), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n258), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT74), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n250), .B1(new_n242), .B2(new_n249), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n247), .B1(new_n255), .B2(new_n256), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n275), .B1(new_n276), .B2(new_n252), .ZN(new_n277));
  INV_X1    g076(.A(new_n271), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n258), .A2(KEYINPUT74), .A3(new_n271), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n274), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G8gat), .B(G36gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT75), .ZN(new_n283));
  XOR2_X1   g082(.A(new_n283), .B(G64gat), .Z(new_n284));
  INV_X1    g083(.A(G92gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n274), .A2(new_n279), .A3(new_n280), .A4(new_n286), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(KEYINPUT30), .A3(new_n289), .ZN(new_n290));
  OR3_X1    g089(.A1(new_n281), .A2(KEYINPUT30), .A3(new_n287), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XOR2_X1   g091(.A(G141gat), .B(G148gat), .Z(new_n293));
  INV_X1    g092(.A(KEYINPUT2), .ZN(new_n294));
  AND2_X1   g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G155gat), .ZN(new_n297));
  INV_X1    g096(.A(G162gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n293), .A2(new_n294), .A3(new_n296), .A4(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT77), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT76), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT76), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(G155gat), .B2(G162gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n302), .B1(new_n306), .B2(new_n296), .ZN(new_n307));
  AOI211_X1 g106(.A(KEYINPUT77), .B(new_n295), .C1(new_n303), .C2(new_n305), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n301), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT70), .B(G120gat), .ZN(new_n312));
  INV_X1    g111(.A(G113gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(G127gat), .B(G134gat), .Z(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT1), .B1(new_n312), .B2(new_n313), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT1), .B1(G113gat), .B2(G120gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n319), .B1(G113gat), .B2(G120gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT4), .B1(new_n311), .B2(new_n322), .ZN(new_n323));
  NOR3_X1   g122(.A1(new_n304), .A2(G155gat), .A3(G162gat), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT76), .B1(new_n297), .B2(new_n298), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n296), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT77), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n306), .A2(new_n302), .A3(new_n296), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(new_n310), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n300), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT4), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n316), .A2(new_n317), .B1(new_n315), .B2(new_n320), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n323), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT5), .ZN(new_n335));
  NAND2_X1  g134(.A1(G225gat), .A2(G233gat), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT3), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n330), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n329), .A2(KEYINPUT3), .A3(new_n300), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n322), .A3(new_n339), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n334), .A2(new_n335), .A3(new_n336), .A4(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n332), .B1(new_n330), .B2(new_n337), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n323), .A2(new_n333), .B1(new_n344), .B2(new_n339), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n345), .A2(KEYINPUT78), .A3(new_n335), .A4(new_n336), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G1gat), .B(G29gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT0), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(G57gat), .ZN(new_n350));
  INV_X1    g149(.A(G85gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n330), .B(new_n332), .ZN(new_n353));
  INV_X1    g152(.A(new_n336), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n334), .A2(new_n340), .ZN(new_n356));
  OAI211_X1 g155(.A(KEYINPUT5), .B(new_n355), .C1(new_n356), .C2(new_n354), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n347), .A2(new_n352), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT6), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n359), .B1(new_n358), .B2(new_n360), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n352), .B1(new_n347), .B2(new_n357), .ZN(new_n363));
  NOR3_X1   g162(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(KEYINPUT6), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT80), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n363), .A2(KEYINPUT80), .A3(KEYINPUT6), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n292), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT29), .B1(new_n268), .B2(new_n270), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n311), .B1(new_n371), .B2(KEYINPUT3), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT81), .ZN(new_n373));
  NAND2_X1  g172(.A1(G228gat), .A2(G233gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(G78gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT31), .B(G50gat), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(G78gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n373), .A2(new_n379), .A3(new_n374), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n376), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n379), .B1(new_n373), .B2(new_n374), .ZN(new_n382));
  INV_X1    g181(.A(new_n374), .ZN(new_n383));
  AOI211_X1 g182(.A(G78gat), .B(new_n383), .C1(new_n372), .C2(KEYINPUT81), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n377), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G22gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n338), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n278), .B1(KEYINPUT29), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n387), .B1(new_n389), .B2(new_n372), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(G106gat), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n389), .A2(new_n372), .A3(new_n387), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n393), .ZN(new_n395));
  OAI21_X1  g194(.A(G106gat), .B1(new_n395), .B2(new_n390), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n386), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n381), .A2(new_n385), .A3(new_n396), .A4(new_n394), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G15gat), .B(G43gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(G71gat), .ZN(new_n402));
  INV_X1    g201(.A(G99gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n276), .A2(new_n332), .ZN(new_n405));
  INV_X1    g204(.A(G227gat), .ZN(new_n406));
  INV_X1    g205(.A(G233gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n322), .B(new_n247), .C1(new_n255), .C2(new_n256), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n405), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n404), .B1(new_n411), .B2(KEYINPUT33), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n408), .B1(new_n405), .B2(new_n409), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT34), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n415), .B1(new_n410), .B2(KEYINPUT32), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n410), .A2(KEYINPUT32), .A3(new_n415), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n414), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n418), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n420), .A2(new_n416), .A3(new_n413), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n412), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n413), .B1(new_n420), .B2(new_n416), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n417), .A2(new_n418), .A3(new_n414), .ZN(new_n424));
  INV_X1    g223(.A(new_n412), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n400), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT35), .B1(new_n370), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT84), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT83), .ZN(new_n430));
  INV_X1    g229(.A(new_n426), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n425), .B1(new_n423), .B2(new_n424), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n422), .A2(KEYINPUT83), .A3(new_n426), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n369), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n347), .A2(new_n357), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n352), .B(KEYINPUT82), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n439), .A2(new_n360), .A3(new_n358), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT35), .B1(new_n290), .B2(new_n291), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n435), .A2(new_n400), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT84), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n444), .B(KEYINPUT35), .C1(new_n370), .C2(new_n427), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n431), .A2(new_n432), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT36), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n356), .A2(new_n354), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n449), .A2(KEYINPUT39), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n450), .A2(new_n438), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n449), .B(KEYINPUT39), .C1(new_n354), .C2(new_n353), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OR2_X1    g252(.A1(new_n453), .A2(KEYINPUT40), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n453), .A2(KEYINPUT40), .B1(new_n437), .B2(new_n438), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n454), .A2(new_n455), .A3(new_n291), .A4(new_n290), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT37), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n274), .A2(new_n279), .A3(new_n457), .A4(new_n280), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n287), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n277), .A2(new_n271), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n258), .A2(new_n278), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n460), .A2(KEYINPUT37), .A3(new_n461), .ZN(new_n462));
  OR3_X1    g261(.A1(new_n459), .A2(KEYINPUT38), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n436), .A2(new_n440), .A3(new_n463), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n281), .A2(KEYINPUT37), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT38), .B1(new_n465), .B2(new_n459), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n289), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n400), .B(new_n456), .C1(new_n464), .C2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n400), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n370), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n448), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n446), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(G29gat), .A2(G36gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(KEYINPUT14), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G43gat), .B(G50gat), .ZN(new_n476));
  OR2_X1    g275(.A1(new_n476), .A2(KEYINPUT15), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(KEYINPUT15), .ZN(new_n478));
  NAND2_X1  g277(.A1(G29gat), .A2(G36gat), .ZN(new_n479));
  XOR2_X1   g278(.A(new_n479), .B(KEYINPUT85), .Z(new_n480));
  NAND4_X1  g279(.A1(new_n475), .A2(new_n477), .A3(new_n478), .A4(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n479), .ZN(new_n482));
  OAI211_X1 g281(.A(KEYINPUT15), .B(new_n476), .C1(new_n474), .C2(new_n482), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n481), .A2(new_n483), .A3(KEYINPUT17), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n483), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT86), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  XOR2_X1   g286(.A(KEYINPUT87), .B(KEYINPUT17), .Z(new_n488));
  AOI21_X1  g287(.A(new_n484), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G99gat), .A2(G106gat), .ZN(new_n490));
  AOI22_X1  g289(.A1(KEYINPUT8), .A2(new_n490), .B1(new_n351), .B2(new_n285), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(KEYINPUT94), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT7), .ZN(new_n493));
  OAI211_X1 g292(.A(KEYINPUT93), .B(new_n493), .C1(new_n351), .C2(new_n285), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n493), .A2(KEYINPUT93), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(KEYINPUT93), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n495), .A2(G85gat), .A3(G92gat), .A4(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n492), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  XOR2_X1   g297(.A(G99gat), .B(G106gat), .Z(new_n499));
  OR2_X1    g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n499), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n489), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n504));
  INV_X1    g303(.A(new_n487), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n503), .B(new_n504), .C1(new_n502), .C2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(G134gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(G190gat), .B(G218gat), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n507), .A2(new_n508), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(G162gat), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n513), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G71gat), .B(G78gat), .ZN(new_n517));
  XOR2_X1   g316(.A(G57gat), .B(G64gat), .Z(new_n518));
  OR2_X1    g317(.A1(new_n518), .A2(KEYINPUT90), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT9), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n520), .B1(new_n518), .B2(KEYINPUT90), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n517), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT91), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n524), .ZN(new_n526));
  AND4_X1   g325(.A1(new_n525), .A2(new_n518), .A3(new_n526), .A4(new_n517), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT21), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT92), .B(KEYINPUT21), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(new_n522), .B2(new_n527), .ZN(new_n531));
  XNOR2_X1  g330(.A(G15gat), .B(G22gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT16), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n532), .B1(new_n533), .B2(G1gat), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(G1gat), .B2(new_n532), .ZN(new_n535));
  INV_X1    g334(.A(G8gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n529), .A2(new_n531), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(new_n531), .B2(new_n537), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n540));
  XNOR2_X1  g339(.A(G155gat), .B(G183gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n539), .B(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G231gat), .A2(G233gat), .ZN(new_n544));
  INV_X1    g343(.A(G127gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(G211gat), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n543), .B(new_n547), .Z(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n516), .A2(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n472), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n537), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT88), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n552), .A2(KEYINPUT88), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n489), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n487), .A2(new_n552), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G229gat), .A2(G233gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT18), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n487), .B(new_n552), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n558), .B(KEYINPUT13), .Z(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n557), .A2(KEYINPUT18), .A3(new_n558), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n561), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G113gat), .B(G141gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G197gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT11), .ZN(new_n569));
  INV_X1    g368(.A(G169gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n571), .B(KEYINPUT12), .Z(new_n572));
  NAND2_X1  g371(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n572), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n561), .A2(new_n574), .A3(new_n564), .A4(new_n565), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT89), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n580));
  INV_X1    g379(.A(new_n499), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n528), .B1(KEYINPUT95), .B2(new_n581), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n502), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n502), .A2(new_n582), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n580), .B1(new_n585), .B2(KEYINPUT10), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT10), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n583), .A2(KEYINPUT96), .A3(new_n587), .A4(new_n584), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n500), .A2(KEYINPUT10), .A3(new_n528), .A4(new_n501), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G230gat), .A2(G233gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n592), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n585), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G120gat), .B(G148gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT97), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n598), .B(G176gat), .Z(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(G204gat), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n596), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n579), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n551), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n364), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(new_n436), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(G1gat), .ZN(G1324gat));
  INV_X1    g410(.A(new_n292), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n606), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n613), .B(KEYINPUT98), .Z(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(G8gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT16), .B(G8gat), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT42), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n614), .A2(new_n616), .ZN(new_n619));
  OAI221_X1 g418(.A(new_n615), .B1(new_n613), .B2(new_n618), .C1(new_n619), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g419(.A(new_n448), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n606), .A2(G15gat), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n435), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n605), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n622), .B1(G15gat), .B2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n625), .B(KEYINPUT99), .Z(G1326gat));
  NOR2_X1   g425(.A1(new_n605), .A2(new_n400), .ZN(new_n627));
  XOR2_X1   g426(.A(KEYINPUT43), .B(G22gat), .Z(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(G1327gat));
  INV_X1    g428(.A(new_n516), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n630), .B1(new_n446), .B2(new_n471), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n603), .A2(new_n548), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n632), .A2(new_n579), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(G29gat), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n635), .A2(new_n636), .A3(new_n609), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT45), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n472), .A2(KEYINPUT100), .A3(new_n516), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT44), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n631), .A2(KEYINPUT100), .A3(KEYINPUT44), .ZN(new_n642));
  INV_X1    g441(.A(new_n576), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n634), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n641), .A2(KEYINPUT101), .A3(new_n642), .A4(new_n644), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n608), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n638), .B1(new_n636), .B2(new_n649), .ZN(G1328gat));
  INV_X1    g449(.A(G36gat), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n651), .A3(new_n612), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n652), .B(KEYINPUT46), .Z(new_n653));
  AOI21_X1  g452(.A(new_n292), .B1(new_n647), .B2(new_n648), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n653), .B1(new_n651), .B2(new_n654), .ZN(G1329gat));
  OAI21_X1  g454(.A(G43gat), .B1(new_n645), .B2(new_n448), .ZN(new_n656));
  INV_X1    g455(.A(G43gat), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n635), .A2(new_n657), .A3(new_n435), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n656), .A2(KEYINPUT47), .A3(new_n658), .ZN(new_n659));
  AND4_X1   g458(.A1(KEYINPUT100), .A2(new_n472), .A3(KEYINPUT44), .A4(new_n516), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT44), .B1(new_n631), .B2(KEYINPUT100), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT101), .B1(new_n662), .B2(new_n644), .ZN(new_n663));
  INV_X1    g462(.A(new_n648), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n621), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(new_n666), .A3(G43gat), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n448), .B1(new_n647), .B2(new_n648), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT102), .B1(new_n668), .B2(new_n657), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n667), .A2(new_n658), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n659), .B1(new_n670), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g470(.A(G50gat), .B1(new_n645), .B2(new_n400), .ZN(new_n672));
  INV_X1    g471(.A(G50gat), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n635), .A2(new_n673), .A3(new_n469), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n672), .A2(KEYINPUT48), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n674), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n469), .B1(new_n663), .B2(new_n664), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n676), .B1(new_n677), .B2(G50gat), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n675), .B1(new_n678), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g478(.A1(new_n551), .A2(new_n603), .A3(new_n643), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n609), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g482(.A1(new_n680), .A2(new_n292), .ZN(new_n684));
  NOR2_X1   g483(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT49), .B(G64gat), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n686), .B1(new_n684), .B2(new_n687), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT103), .Z(G1333gat));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n681), .A2(KEYINPUT104), .A3(G71gat), .A4(new_n621), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n551), .A2(G71gat), .A3(new_n603), .A4(new_n643), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n692), .B1(new_n693), .B2(new_n448), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(G71gat), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(new_n680), .B2(new_n623), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n690), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n695), .A2(new_n690), .A3(new_n697), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT50), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n700), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT50), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n702), .A2(new_n703), .A3(new_n698), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n701), .A2(new_n704), .ZN(G1334gat));
  NOR2_X1   g504(.A1(new_n680), .A2(new_n400), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(new_n379), .ZN(G1335gat));
  NOR2_X1   g506(.A1(new_n576), .A2(new_n548), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n472), .A2(new_n516), .A3(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(KEYINPUT107), .B1(new_n710), .B2(KEYINPUT51), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(KEYINPUT51), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n713), .A2(new_n351), .A3(new_n609), .A4(new_n603), .ZN(new_n714));
  INV_X1    g513(.A(new_n708), .ZN(new_n715));
  INV_X1    g514(.A(new_n603), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n641), .A2(new_n642), .A3(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n641), .A2(KEYINPUT106), .A3(new_n642), .A4(new_n717), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n608), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n714), .B1(new_n351), .B2(new_n722), .ZN(G1336gat));
  NOR3_X1   g522(.A1(new_n716), .A2(G92gat), .A3(new_n292), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n713), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT52), .ZN(new_n726));
  OAI21_X1  g525(.A(G92gat), .B1(new_n718), .B2(new_n292), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT106), .B1(new_n662), .B2(new_n717), .ZN(new_n729));
  INV_X1    g528(.A(new_n721), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n612), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n709), .A2(KEYINPUT108), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT51), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n631), .A2(new_n734), .A3(new_n708), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n732), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n732), .A2(KEYINPUT109), .A3(new_n733), .A4(new_n735), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(new_n712), .A3(new_n739), .ZN(new_n740));
  AOI22_X1  g539(.A1(new_n731), .A2(G92gat), .B1(new_n724), .B2(new_n740), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n741), .A2(KEYINPUT110), .A3(new_n726), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n738), .A2(new_n712), .A3(new_n739), .ZN(new_n744));
  INV_X1    g543(.A(new_n724), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n292), .B1(new_n720), .B2(new_n721), .ZN(new_n746));
  OAI22_X1  g545(.A1(new_n744), .A2(new_n745), .B1(new_n746), .B2(new_n285), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n743), .B1(new_n747), .B2(KEYINPUT52), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n728), .B1(new_n742), .B2(new_n748), .ZN(G1337gat));
  NAND3_X1  g548(.A1(new_n435), .A2(new_n603), .A3(new_n403), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT111), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n713), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n448), .B1(new_n720), .B2(new_n721), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n403), .B2(new_n753), .ZN(G1338gat));
  NOR3_X1   g553(.A1(new_n716), .A2(G106gat), .A3(new_n400), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n713), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT53), .ZN(new_n757));
  OAI21_X1  g556(.A(G106gat), .B1(new_n718), .B2(new_n400), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n469), .B1(new_n729), .B2(new_n730), .ZN(new_n760));
  AOI22_X1  g559(.A1(new_n760), .A2(G106gat), .B1(new_n740), .B2(new_n755), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(new_n761), .B2(new_n757), .ZN(G1339gat));
  NOR2_X1   g561(.A1(new_n608), .A2(new_n612), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n589), .A2(new_n594), .A3(new_n590), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n593), .A2(KEYINPUT54), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n591), .A2(new_n592), .A3(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n766), .A2(KEYINPUT55), .A3(new_n600), .A4(new_n768), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n769), .A2(new_n601), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n766), .A2(new_n600), .A3(new_n768), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n770), .A2(KEYINPUT113), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n771), .A2(new_n772), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n769), .A2(new_n601), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n643), .B1(new_n774), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n557), .A2(new_n558), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n562), .A2(new_n563), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n571), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n575), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n716), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n630), .B1(new_n779), .B2(new_n784), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n783), .B(KEYINPUT114), .Z(new_n786));
  NOR2_X1   g585(.A1(new_n630), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n774), .A2(new_n778), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n549), .ZN(new_n791));
  NOR4_X1   g590(.A1(new_n516), .A2(new_n549), .A3(new_n603), .A4(new_n576), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n764), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n623), .A2(new_n469), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(G113gat), .B1(new_n796), .B2(new_n579), .ZN(new_n797));
  INV_X1    g596(.A(new_n427), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n576), .A2(new_n313), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n797), .B1(new_n799), .B2(new_n800), .ZN(G1340gat));
  OAI21_X1  g600(.A(G120gat), .B1(new_n796), .B2(new_n716), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n716), .A2(G120gat), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n799), .B2(new_n803), .ZN(G1341gat));
  NOR3_X1   g603(.A1(new_n796), .A2(new_n545), .A3(new_n549), .ZN(new_n805));
  INV_X1    g604(.A(new_n799), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n548), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n805), .B1(new_n545), .B2(new_n807), .ZN(G1342gat));
  OR3_X1    g607(.A1(new_n799), .A2(G134gat), .A3(new_n630), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n809), .A2(KEYINPUT56), .ZN(new_n810));
  OAI21_X1  g609(.A(G134gat), .B1(new_n796), .B2(new_n630), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(KEYINPUT56), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(G1343gat));
  INV_X1    g612(.A(G141gat), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n548), .B1(new_n785), .B2(new_n789), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n469), .B1(new_n815), .B2(new_n792), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n816), .A2(KEYINPUT57), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n621), .A2(new_n764), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n771), .B(new_n819), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n578), .B(new_n770), .C1(new_n820), .C2(KEYINPUT55), .ZN(new_n821));
  INV_X1    g620(.A(new_n784), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n516), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n548), .B1(new_n824), .B2(new_n789), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n469), .B1(new_n825), .B2(new_n792), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT57), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n817), .A2(new_n818), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n814), .B1(new_n829), .B2(new_n578), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n621), .A2(new_n400), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT116), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n794), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n832), .A2(KEYINPUT116), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n834), .A2(G141gat), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n578), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT58), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n817), .A2(new_n827), .A3(new_n576), .A4(new_n818), .ZN(new_n840));
  AOI22_X1  g639(.A1(G141gat), .A2(new_n840), .B1(new_n836), .B2(new_n578), .ZN(new_n841));
  OAI22_X1  g640(.A1(new_n830), .A2(new_n839), .B1(new_n841), .B2(new_n838), .ZN(G1344gat));
  NOR2_X1   g641(.A1(new_n834), .A2(new_n835), .ZN(new_n843));
  INV_X1    g642(.A(G148gat), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(new_n844), .A3(new_n603), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n816), .A2(KEYINPUT57), .ZN(new_n847));
  NOR4_X1   g646(.A1(new_n630), .A2(new_n777), .A3(new_n786), .A4(new_n776), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n549), .B1(new_n823), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n550), .A2(new_n716), .A3(new_n579), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT57), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n469), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n847), .A2(new_n852), .A3(new_n603), .A4(new_n818), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n844), .B1(new_n853), .B2(KEYINPUT117), .ZN(new_n854));
  AOI22_X1  g653(.A1(new_n816), .A2(KEYINPUT57), .B1(new_n851), .B2(new_n469), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n855), .A2(new_n856), .A3(new_n603), .A4(new_n818), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n846), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n817), .A2(new_n827), .A3(new_n603), .A4(new_n818), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n859), .A2(new_n846), .A3(G148gat), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n845), .B1(new_n858), .B2(new_n860), .ZN(G1345gat));
  NOR3_X1   g660(.A1(new_n828), .A2(new_n297), .A3(new_n549), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n834), .A2(new_n549), .A3(new_n835), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT118), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n862), .B1(new_n864), .B2(new_n297), .ZN(G1346gat));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n829), .A2(new_n866), .A3(new_n516), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT119), .B1(new_n828), .B2(new_n630), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(G162gat), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n843), .A2(new_n298), .A3(new_n516), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(G1347gat));
  OAI211_X1 g670(.A(new_n608), .B(new_n612), .C1(new_n815), .C2(new_n792), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n427), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n570), .A3(new_n576), .ZN(new_n874));
  INV_X1    g673(.A(new_n795), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n872), .A2(new_n875), .A3(new_n579), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n874), .B1(new_n570), .B2(new_n876), .ZN(G1348gat));
  INV_X1    g676(.A(new_n872), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n878), .A2(G176gat), .A3(new_n795), .A4(new_n603), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT121), .ZN(new_n880));
  AOI21_X1  g679(.A(G176gat), .B1(new_n873), .B2(new_n603), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n881), .A2(KEYINPUT120), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(KEYINPUT120), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(G1349gat));
  INV_X1    g683(.A(KEYINPUT60), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n609), .B1(new_n791), .B2(new_n793), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n215), .A2(new_n216), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n549), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n886), .A2(new_n612), .A3(new_n798), .A4(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT123), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n872), .A2(new_n549), .A3(new_n875), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n889), .B(new_n890), .C1(new_n891), .C2(new_n211), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n885), .B1(new_n893), .B2(KEYINPUT122), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n889), .B(KEYINPUT122), .C1(new_n891), .C2(new_n211), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n892), .A2(new_n896), .A3(KEYINPUT60), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n894), .A2(new_n895), .A3(new_n897), .ZN(G1350gat));
  NAND3_X1  g697(.A1(new_n873), .A2(new_n209), .A3(new_n516), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n886), .A2(new_n516), .A3(new_n612), .A4(new_n795), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n900), .A2(new_n901), .A3(G190gat), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n900), .B2(G190gat), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g705(.A(KEYINPUT124), .B(new_n899), .C1(new_n902), .C2(new_n903), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1351gat));
  NOR3_X1   g707(.A1(new_n621), .A2(new_n609), .A3(new_n292), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n847), .A2(new_n852), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(KEYINPUT127), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT127), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n855), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n909), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(G197gat), .B1(new_n914), .B2(new_n579), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT125), .B1(new_n831), .B2(new_n612), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n831), .A2(KEYINPUT125), .A3(new_n612), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n886), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n919), .A2(G197gat), .A3(new_n643), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT126), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n920), .B(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n915), .A2(new_n922), .ZN(G1352gat));
  OAI21_X1  g722(.A(G204gat), .B1(new_n914), .B2(new_n716), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n919), .A2(G204gat), .A3(new_n716), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT62), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1353gat));
  NAND2_X1  g726(.A1(new_n909), .A2(new_n548), .ZN(new_n928));
  OAI21_X1  g727(.A(G211gat), .B1(new_n910), .B2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT63), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n929), .B(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n919), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(new_n262), .A3(new_n548), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1354gat));
  AOI21_X1  g733(.A(G218gat), .B1(new_n932), .B2(new_n516), .ZN(new_n935));
  INV_X1    g734(.A(new_n914), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n630), .A2(new_n261), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(G1355gat));
endmodule


