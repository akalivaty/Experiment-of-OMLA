//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 1 0 1 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n553, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n569, new_n570, new_n571, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT65), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT66), .Z(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n457), .A2(G567), .ZN(new_n460));
  INV_X1    g035(.A(G2106), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n454), .B2(new_n461), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT67), .Z(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  XNOR2_X1  g042(.A(new_n466), .B(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G137), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n476), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n468), .B(new_n474), .C1(new_n475), .C2(new_n477), .ZN(new_n478));
  XOR2_X1   g053(.A(new_n478), .B(KEYINPUT69), .Z(G160));
  NAND2_X1  g054(.A1(new_n476), .A2(G2105), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT70), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n473), .A2(G136), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND4_X1  g062(.A1(new_n469), .A2(new_n471), .A3(G126), .A4(G2105), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n476), .A2(KEYINPUT71), .A3(G126), .A4(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(new_n475), .B2(G114), .ZN(new_n493));
  NOR2_X1   g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT72), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n476), .A2(G138), .A3(new_n475), .ZN(new_n500));
  XNOR2_X1  g075(.A(new_n500), .B(KEYINPUT4), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n492), .A2(KEYINPUT72), .A3(new_n496), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n499), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G62), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n505), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI211_X1 g095(.A(new_n507), .B(new_n509), .C1(new_n515), .C2(new_n516), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n523));
  OR3_X1    g098(.A1(new_n514), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n514), .B2(new_n522), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(G166));
  AOI22_X1  g101(.A1(new_n517), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n527), .A2(new_n510), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n515), .A2(new_n516), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n506), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G51), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n528), .A2(new_n531), .A3(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  OAI211_X1 g110(.A(G52), .B(G543), .C1(new_n515), .C2(new_n516), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n521), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n507), .A2(new_n509), .A3(G64), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n505), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n542));
  OR3_X1    g117(.A1(new_n538), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n538), .B2(new_n541), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(G171));
  AOI22_X1  g120(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n505), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT75), .B(G43), .Z(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n518), .A2(new_n548), .B1(new_n549), .B2(new_n521), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n553), .A2(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(new_n530), .A2(G53), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n521), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G91), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n563), .B2(new_n505), .ZN(new_n564));
  OR3_X1    g139(.A1(new_n560), .A2(KEYINPUT76), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT76), .B1(new_n560), .B2(new_n564), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  NOR2_X1   g143(.A1(G166), .A2(KEYINPUT77), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(new_n524), .B2(new_n525), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n569), .A2(new_n571), .ZN(G303));
  NAND2_X1  g147(.A1(new_n561), .A2(G87), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n530), .A2(G49), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT78), .ZN(new_n578));
  AND3_X1   g153(.A1(new_n507), .A2(new_n509), .A3(G61), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(G48), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n518), .A2(new_n583), .B1(new_n584), .B2(new_n521), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n505), .ZN(new_n589));
  XNOR2_X1  g164(.A(KEYINPUT80), .B(G47), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n518), .A2(new_n590), .B1(new_n591), .B2(new_n521), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n589), .A2(new_n592), .ZN(G290));
  INV_X1    g168(.A(G92), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n521), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT10), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n510), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(new_n530), .B2(G54), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n602), .B2(G171), .ZN(G284));
  XOR2_X1   g179(.A(G284), .B(KEYINPUT81), .Z(G321));
  NOR2_X1   g180(.A1(G286), .A2(new_n602), .ZN(new_n606));
  INV_X1    g181(.A(G299), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(new_n602), .ZN(G297));
  AOI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(new_n602), .ZN(G280));
  INV_X1    g184(.A(new_n601), .ZN(new_n610));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G860), .ZN(G148));
  NOR2_X1   g187(.A1(new_n601), .A2(G559), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT82), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n615), .B(KEYINPUT83), .C1(G868), .C2(new_n551), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(KEYINPUT83), .B2(new_n615), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT84), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n481), .A2(G123), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n473), .A2(G135), .ZN(new_n621));
  NOR2_X1   g196(.A1(G99), .A2(G2105), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(new_n475), .B2(G111), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n620), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2096), .Z(new_n625));
  NAND2_X1  g200(.A1(new_n476), .A2(new_n465), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT12), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n625), .A2(new_n630), .ZN(G156));
  XOR2_X1   g206(.A(KEYINPUT15), .B(G2435), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2438), .ZN(new_n633));
  XOR2_X1   g208(.A(G2427), .B(G2430), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT85), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n633), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(KEYINPUT14), .ZN(new_n637));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G1341), .B(G1348), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n642), .B(new_n643), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(G14), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(G401));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  XOR2_X1   g222(.A(G2067), .B(G2678), .Z(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n647), .B1(new_n651), .B2(KEYINPUT18), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2096), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(new_n629), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n649), .A2(new_n650), .ZN(new_n656));
  AOI21_X1  g231(.A(KEYINPUT18), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n654), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n659), .A2(new_n660), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n662), .A2(new_n664), .A3(new_n666), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n669), .B(new_n670), .C1(new_n668), .C2(new_n667), .ZN(new_n671));
  XOR2_X1   g246(.A(G1981), .B(G1986), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1991), .B(G1996), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT86), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(G229));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n679), .A2(KEYINPUT23), .A3(G20), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT23), .ZN(new_n681));
  INV_X1    g256(.A(G20), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n681), .B1(new_n682), .B2(G16), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n680), .B(new_n683), .C1(new_n607), .C2(new_n679), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(G1956), .Z(new_n685));
  NOR2_X1   g260(.A1(G16), .A2(G19), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n551), .B2(G16), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n687), .A2(G1341), .ZN(new_n688));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n481), .A2(G128), .ZN(new_n690));
  NOR2_X1   g265(.A1(G104), .A2(G2105), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT89), .ZN(new_n692));
  INV_X1    g267(.A(G116), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n464), .B1(new_n693), .B2(G2105), .ZN(new_n694));
  AOI22_X1  g269(.A1(G140), .A2(new_n473), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n689), .B1(new_n690), .B2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G26), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n697), .A2(G29), .ZN(new_n698));
  OAI21_X1  g273(.A(KEYINPUT28), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(KEYINPUT28), .B2(new_n698), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n688), .B1(new_n700), .B2(G2067), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n685), .B(new_n701), .C1(G1341), .C2(new_n687), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n465), .A2(G103), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT90), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(KEYINPUT25), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n703), .B(KEYINPUT90), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT25), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(G115), .A2(G2104), .ZN(new_n710));
  INV_X1    g285(.A(G127), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n472), .B2(new_n711), .ZN(new_n712));
  AOI22_X1  g287(.A1(new_n712), .A2(G2105), .B1(new_n473), .B2(G139), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n706), .A2(new_n709), .A3(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G29), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G29), .B2(G33), .ZN(new_n717));
  INV_X1    g292(.A(G2072), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT91), .ZN(new_n720));
  NOR2_X1   g295(.A1(G16), .A2(G21), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G168), .B2(G16), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n722), .A2(G1966), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT92), .Z(new_n724));
  OR2_X1    g299(.A1(KEYINPUT24), .A2(G34), .ZN(new_n725));
  NAND2_X1  g300(.A1(KEYINPUT24), .A2(G34), .ZN(new_n726));
  AOI21_X1  g301(.A(G29), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G160), .B2(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G2084), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n689), .A2(G27), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G164), .B2(new_n689), .ZN(new_n731));
  INV_X1    g306(.A(G2078), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n720), .A2(new_n724), .A3(new_n729), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n481), .A2(G129), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n465), .A2(G105), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n473), .A2(G141), .ZN(new_n737));
  NAND3_X1  g312(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT26), .Z(new_n739));
  NAND4_X1  g314(.A1(new_n735), .A2(new_n736), .A3(new_n737), .A4(new_n739), .ZN(new_n740));
  MUX2_X1   g315(.A(G32), .B(new_n740), .S(G29), .Z(new_n741));
  XOR2_X1   g316(.A(KEYINPUT27), .B(G1996), .Z(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT30), .B(G28), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n743), .B1(new_n689), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n722), .A2(G1966), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n624), .A2(new_n689), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n741), .A2(new_n742), .B1(new_n717), .B2(new_n718), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n745), .A2(new_n746), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n679), .A2(G5), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G171), .B2(new_n679), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n751), .A2(G1961), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(G1961), .ZN(new_n753));
  OAI221_X1 g328(.A(new_n752), .B1(KEYINPUT93), .B2(new_n753), .C1(new_n728), .C2(G2084), .ZN(new_n754));
  NOR3_X1   g329(.A1(new_n734), .A2(new_n749), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT31), .B(G11), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n753), .A2(KEYINPUT93), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n702), .B1(new_n758), .B2(KEYINPUT94), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT94), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n755), .A2(new_n760), .A3(new_n756), .A4(new_n757), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n679), .A2(G23), .ZN(new_n762));
  INV_X1    g337(.A(G288), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(new_n679), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT88), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT33), .B(G1976), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  MUX2_X1   g342(.A(G6), .B(G305), .S(G16), .Z(new_n768));
  XOR2_X1   g343(.A(KEYINPUT32), .B(G1981), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G16), .A2(G22), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G166), .B2(G16), .ZN(new_n772));
  INV_X1    g347(.A(G1971), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n767), .A2(new_n770), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT34), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n481), .A2(G119), .ZN(new_n777));
  NOR2_X1   g352(.A1(G95), .A2(G2105), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT87), .ZN(new_n779));
  INV_X1    g354(.A(G107), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n464), .B1(new_n780), .B2(G2105), .ZN(new_n781));
  AOI22_X1  g356(.A1(G131), .A2(new_n473), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n777), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n783), .A2(new_n689), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G25), .B2(new_n689), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT35), .B(G1991), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n785), .A2(new_n787), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n679), .A2(G24), .ZN(new_n790));
  INV_X1    g365(.A(G290), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(new_n679), .ZN(new_n792));
  INV_X1    g367(.A(G1986), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n788), .A2(new_n789), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n776), .A2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT36), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n776), .A2(KEYINPUT36), .A3(new_n795), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n759), .B(new_n761), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n700), .A2(G2067), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n679), .A2(G4), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n610), .B2(new_n679), .ZN(new_n803));
  INV_X1    g378(.A(G1348), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(G29), .A2(G35), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G162), .B2(G29), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT29), .ZN(new_n809));
  INV_X1    g384(.A(G2090), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  NOR4_X1   g387(.A1(new_n800), .A2(new_n801), .A3(new_n806), .A4(new_n812), .ZN(G311));
  NOR2_X1   g388(.A1(new_n800), .A2(new_n812), .ZN(new_n814));
  INV_X1    g389(.A(new_n801), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n814), .A2(new_n815), .A3(new_n805), .ZN(G150));
  NAND2_X1  g391(.A1(G80), .A2(G543), .ZN(new_n817));
  INV_X1    g392(.A(G67), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n510), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G651), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(KEYINPUT95), .ZN(new_n821));
  INV_X1    g396(.A(G55), .ZN(new_n822));
  INV_X1    g397(.A(G93), .ZN(new_n823));
  OAI22_X1  g398(.A1(new_n518), .A2(new_n822), .B1(new_n823), .B2(new_n521), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n820), .A2(KEYINPUT95), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n821), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G860), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT37), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n610), .A2(G559), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT38), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT39), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n821), .A2(new_n826), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT96), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n833), .A2(new_n551), .A3(new_n834), .A4(new_n825), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n551), .A2(new_n834), .ZN(new_n836));
  OAI21_X1  g411(.A(KEYINPUT96), .B1(new_n547), .B2(new_n550), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n836), .A2(new_n837), .A3(new_n827), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n832), .B(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n829), .B1(new_n841), .B2(G860), .ZN(G145));
  NAND2_X1  g417(.A1(new_n473), .A2(G142), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT99), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n481), .A2(G130), .ZN(new_n846));
  OR2_X1    g421(.A1(G106), .A2(G2105), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n847), .B(G2104), .C1(G118), .C2(new_n475), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(new_n783), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT100), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n777), .A2(new_n782), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n852), .A2(new_n846), .A3(new_n848), .A4(new_n845), .ZN(new_n853));
  AND3_X1   g428(.A1(new_n850), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n851), .B1(new_n850), .B2(new_n853), .ZN(new_n855));
  INV_X1    g430(.A(new_n627), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n850), .A2(new_n853), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(KEYINPUT100), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n850), .A2(new_n853), .A3(new_n851), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n627), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(KEYINPUT98), .B1(new_n492), .B2(new_n496), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n864));
  AOI211_X1 g439(.A(new_n864), .B(new_n495), .C1(new_n490), .C2(new_n491), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n501), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n690), .A2(new_n695), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n868), .A2(new_n740), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n740), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n714), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(new_n715), .A3(new_n870), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n862), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT101), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n862), .A2(new_n872), .A3(KEYINPUT101), .A4(new_n873), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n877), .B1(new_n876), .B2(new_n878), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n872), .A2(new_n873), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n881), .A2(new_n862), .ZN(new_n882));
  NOR3_X1   g457(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(G160), .B(KEYINPUT97), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n486), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n624), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT40), .ZN(new_n888));
  INV_X1    g463(.A(G37), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n862), .B1(new_n881), .B2(KEYINPUT103), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n890), .B1(KEYINPUT103), .B2(new_n881), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n876), .A2(new_n878), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(new_n886), .A3(new_n892), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n887), .A2(new_n888), .A3(new_n889), .A4(new_n893), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n889), .B(new_n893), .C1(new_n883), .C2(new_n886), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT40), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(G395));
  NAND2_X1  g472(.A1(new_n827), .A2(new_n602), .ZN(new_n898));
  XNOR2_X1  g473(.A(G166), .B(G290), .ZN(new_n899));
  XNOR2_X1  g474(.A(G305), .B(new_n763), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n899), .B(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  XOR2_X1   g477(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(new_n904), .B(KEYINPUT107), .Z(new_n905));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n905), .B1(new_n906), .B2(new_n902), .ZN(new_n907));
  INV_X1    g482(.A(new_n566), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n560), .A2(KEYINPUT76), .A3(new_n564), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n908), .A2(new_n909), .A3(new_n601), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n610), .B1(new_n565), .B2(new_n566), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n910), .B2(new_n911), .ZN(new_n914));
  NOR3_X1   g489(.A1(new_n910), .A2(new_n911), .A3(KEYINPUT41), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n914), .A2(new_n916), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n614), .B(new_n840), .ZN(new_n920));
  MUX2_X1   g495(.A(new_n912), .B(new_n919), .S(new_n920), .Z(new_n921));
  XNOR2_X1  g496(.A(new_n907), .B(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n898), .B1(new_n922), .B2(new_n602), .ZN(G295));
  OAI21_X1  g498(.A(new_n898), .B1(new_n922), .B2(new_n602), .ZN(G331));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n543), .A2(new_n544), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(G286), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT109), .ZN(new_n929));
  NAND2_X1  g504(.A1(G171), .A2(KEYINPUT108), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT109), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n927), .A2(G286), .A3(new_n931), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n930), .B1(new_n929), .B2(new_n932), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n839), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n932), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n931), .B1(new_n927), .B2(G286), .ZN(new_n937));
  OAI211_X1 g512(.A(KEYINPUT108), .B(G171), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n840), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT41), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(new_n910), .B2(new_n911), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n601), .B1(new_n908), .B2(new_n909), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n565), .A2(new_n566), .A3(new_n610), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(new_n944), .A3(new_n913), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n935), .A2(new_n940), .A3(new_n942), .A4(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n940), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n840), .B1(new_n938), .B2(new_n939), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n912), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n946), .A2(new_n947), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n902), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n949), .A2(new_n950), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n919), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(new_n901), .A3(new_n951), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(new_n957), .A3(new_n889), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT111), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n954), .A2(new_n957), .A3(new_n960), .A4(new_n889), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n925), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n956), .A2(new_n951), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n902), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(new_n889), .A3(new_n957), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n965), .A2(new_n925), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT44), .B1(new_n962), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n954), .A2(new_n957), .A3(new_n925), .A4(new_n889), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n967), .A2(new_n972), .ZN(G397));
  NAND2_X1  g548(.A1(new_n497), .A2(new_n864), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n492), .A2(KEYINPUT98), .A3(new_n496), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(G1384), .B1(new_n976), .B2(new_n501), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n977), .B(KEYINPUT112), .ZN(new_n978));
  XNOR2_X1  g553(.A(KEYINPUT113), .B(KEYINPUT45), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G40), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n478), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(G1996), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n984), .A2(KEYINPUT46), .ZN(new_n985));
  INV_X1    g560(.A(new_n983), .ZN(new_n986));
  INV_X1    g561(.A(G2067), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n867), .B(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n986), .B1(new_n740), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n984), .A2(KEYINPUT46), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n985), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT47), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n992), .B(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(G290), .A2(G1986), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n986), .A2(new_n995), .ZN(new_n996));
  XOR2_X1   g571(.A(new_n996), .B(KEYINPUT48), .Z(new_n997));
  XNOR2_X1  g572(.A(new_n740), .B(G1996), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n989), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n783), .A2(new_n787), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n852), .A2(new_n786), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n997), .B1(new_n986), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n867), .A2(G2067), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n1000), .B(KEYINPUT127), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1004), .B1(new_n999), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n983), .A2(new_n1006), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n994), .A2(new_n1003), .A3(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(G303), .A2(KEYINPUT114), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1009));
  OAI21_X1  g584(.A(G8), .B1(new_n569), .B2(new_n571), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1009), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1384), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n866), .A2(KEYINPUT45), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n982), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n979), .B1(new_n503), .B2(new_n1017), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n773), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n982), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n866), .A2(new_n1017), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1022), .B1(new_n1023), .B2(KEYINPUT50), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT72), .B1(new_n492), .B2(new_n496), .ZN(new_n1025));
  AOI211_X1 g600(.A(new_n498), .B(new_n495), .C1(new_n490), .C2(new_n491), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1384), .B1(new_n1027), .B2(new_n501), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n503), .A2(new_n1030), .A3(new_n1017), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT117), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1024), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1021), .B1(new_n1034), .B2(G2090), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT115), .B(G8), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1016), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(G305), .A2(G1981), .ZN(new_n1039));
  INV_X1    g614(.A(G1981), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n582), .A2(new_n1040), .A3(new_n586), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT49), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1036), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(new_n977), .B2(new_n982), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1039), .A2(KEYINPUT49), .A3(new_n1041), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1044), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n977), .A2(new_n982), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n763), .A2(G1976), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(new_n1036), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT52), .ZN(new_n1052));
  INV_X1    g627(.A(G1976), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(G288), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1046), .A2(new_n1050), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1048), .A2(new_n1052), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1048), .A2(new_n1052), .A3(KEYINPUT118), .A4(new_n1055), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n866), .A2(new_n1030), .A3(new_n1017), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1061), .B(new_n982), .C1(new_n1028), .C2(new_n1030), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1021), .B1(G2090), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1015), .A2(G8), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1061), .A2(new_n982), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1030), .B1(new_n503), .B2(new_n1017), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G2084), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n503), .A2(new_n1017), .A3(new_n979), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n982), .B(new_n1069), .C1(new_n977), .C2(KEYINPUT45), .ZN(new_n1070));
  INV_X1    g645(.A(G1966), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1067), .A2(new_n1068), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1072), .A2(G286), .A3(new_n1045), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1038), .A2(new_n1060), .A3(new_n1064), .A4(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT63), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1063), .A2(G8), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1056), .B1(new_n1016), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1078), .A2(new_n1064), .A3(new_n1073), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1076), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1048), .A2(new_n1053), .A3(new_n763), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n1041), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n1046), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n1064), .B2(new_n1056), .ZN(new_n1084));
  XNOR2_X1  g659(.A(new_n1084), .B(KEYINPUT116), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(G168), .A2(new_n1045), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1069), .A2(new_n982), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT45), .B1(new_n866), .B2(new_n1017), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1071), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n503), .A2(new_n1017), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT50), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1092), .A2(new_n1068), .A3(new_n982), .A4(new_n1061), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  AOI211_X1 g669(.A(KEYINPUT51), .B(new_n1087), .C1(new_n1094), .C2(new_n1036), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT126), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1087), .ZN(new_n1098));
  INV_X1    g673(.A(G8), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1098), .B1(new_n1072), .B2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT125), .B(KEYINPUT51), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1097), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1099), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1097), .B(new_n1102), .C1(new_n1104), .C2(new_n1087), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1096), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1072), .A2(new_n1098), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1107), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1087), .B1(new_n1094), .B2(G8), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT126), .B1(new_n1112), .B2(new_n1101), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1095), .B1(new_n1113), .B2(new_n1105), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT62), .B1(new_n1114), .B2(new_n1109), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT53), .B1(new_n1116), .B2(new_n732), .ZN(new_n1117));
  INV_X1    g692(.A(G1961), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1117), .B1(new_n1118), .B2(new_n1062), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n1120));
  OR3_X1    g695(.A1(new_n1070), .A2(new_n1120), .A3(G2078), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1111), .A2(new_n1115), .A3(G171), .A4(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(G171), .B(KEYINPUT54), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1124), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1125), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n560), .B2(new_n564), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n560), .A2(new_n564), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT57), .ZN(new_n1132));
  OAI211_X1 g707(.A(KEYINPUT121), .B(new_n1127), .C1(new_n560), .C2(new_n564), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1130), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT123), .ZN(new_n1135));
  XOR2_X1   g710(.A(KEYINPUT119), .B(G1956), .Z(new_n1136));
  AND2_X1   g711(.A1(new_n1034), .A2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(KEYINPUT56), .B(G2072), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1116), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g714(.A(KEYINPUT124), .B(new_n1135), .C1(new_n1137), .C2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1034), .A2(new_n1136), .B1(new_n1116), .B2(new_n1138), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1134), .B(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1141), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n804), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1146));
  AND4_X1   g721(.A1(new_n1017), .A2(new_n866), .A3(new_n982), .A4(new_n987), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1146), .A2(KEYINPUT122), .A3(new_n1148), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1151), .A2(new_n610), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1140), .A2(new_n1145), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1142), .A2(new_n1134), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AOI211_X1 g731(.A(new_n1150), .B(new_n1147), .C1(new_n1062), .C2(new_n804), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT122), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1157), .A2(new_n1158), .A3(KEYINPUT60), .ZN(new_n1159));
  OAI21_X1  g734(.A(KEYINPUT60), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n610), .ZN(new_n1161));
  OAI211_X1 g736(.A(KEYINPUT60), .B(new_n601), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1159), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n979), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1091), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(G1996), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1165), .A2(new_n1166), .A3(new_n982), .A4(new_n1018), .ZN(new_n1167));
  XOR2_X1   g742(.A(KEYINPUT58), .B(G1341), .Z(new_n1168));
  NAND2_X1  g743(.A1(new_n1049), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n551), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(KEYINPUT59), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT59), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1170), .A2(new_n1173), .A3(new_n551), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1155), .A2(KEYINPUT61), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1142), .A2(new_n1177), .A3(new_n1134), .ZN(new_n1178));
  OR2_X1    g753(.A1(new_n1142), .A2(new_n1134), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1175), .A2(new_n1176), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1156), .B1(new_n1163), .B2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g756(.A(KEYINPUT53), .B(new_n732), .C1(new_n978), .C2(new_n979), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1119), .B(new_n1124), .C1(new_n1019), .C2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1126), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1123), .A2(new_n1184), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1038), .A2(new_n1060), .A3(new_n1064), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1086), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n791), .A2(new_n793), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n1002), .A2(new_n995), .A3(new_n1188), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1189), .A2(new_n983), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1008), .B1(new_n1187), .B2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g766(.A(new_n462), .B1(new_n968), .B2(new_n969), .ZN(new_n1193));
  NOR2_X1   g767(.A1(G229), .A2(G227), .ZN(new_n1194));
  NAND4_X1  g768(.A1(new_n1193), .A2(new_n895), .A3(new_n645), .A4(new_n1194), .ZN(G225));
  INV_X1    g769(.A(G225), .ZN(G308));
endmodule


