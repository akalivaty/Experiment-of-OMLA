

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586;

  XOR2_X1 U326 ( .A(KEYINPUT28), .B(n466), .Z(n529) );
  INV_X1 U327 ( .A(KEYINPUT58), .ZN(n457) );
  XNOR2_X1 U328 ( .A(G120GAT), .B(KEYINPUT83), .ZN(n294) );
  XNOR2_X1 U329 ( .A(n294), .B(KEYINPUT84), .ZN(n295) );
  XOR2_X1 U330 ( .A(n295), .B(KEYINPUT0), .Z(n297) );
  XNOR2_X1 U331 ( .A(G113GAT), .B(G134GAT), .ZN(n296) );
  XNOR2_X1 U332 ( .A(n297), .B(n296), .ZN(n428) );
  XOR2_X1 U333 ( .A(KEYINPUT19), .B(KEYINPUT86), .Z(n299) );
  XNOR2_X1 U334 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n298) );
  XNOR2_X1 U335 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U336 ( .A(G169GAT), .B(n300), .Z(n322) );
  XNOR2_X1 U337 ( .A(n428), .B(n322), .ZN(n313) );
  XOR2_X1 U338 ( .A(G176GAT), .B(G190GAT), .Z(n302) );
  XNOR2_X1 U339 ( .A(G43GAT), .B(G99GAT), .ZN(n301) );
  XNOR2_X1 U340 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U341 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n304) );
  XNOR2_X1 U342 ( .A(G183GAT), .B(G71GAT), .ZN(n303) );
  XNOR2_X1 U343 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U344 ( .A(n306), .B(n305), .Z(n311) );
  XOR2_X1 U345 ( .A(G15GAT), .B(G127GAT), .Z(n371) );
  XOR2_X1 U346 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n308) );
  NAND2_X1 U347 ( .A1(G227GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U348 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U349 ( .A(n371), .B(n309), .ZN(n310) );
  XNOR2_X1 U350 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U351 ( .A(n313), .B(n312), .ZN(n555) );
  XOR2_X1 U352 ( .A(G211GAT), .B(KEYINPUT78), .Z(n315) );
  XNOR2_X1 U353 ( .A(G8GAT), .B(G183GAT), .ZN(n314) );
  XNOR2_X1 U354 ( .A(n315), .B(n314), .ZN(n362) );
  XOR2_X1 U355 ( .A(G197GAT), .B(KEYINPUT21), .Z(n445) );
  XOR2_X1 U356 ( .A(n362), .B(n445), .Z(n317) );
  NAND2_X1 U357 ( .A1(G226GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U358 ( .A(n317), .B(n316), .ZN(n320) );
  XOR2_X1 U359 ( .A(G64GAT), .B(G204GAT), .Z(n319) );
  XNOR2_X1 U360 ( .A(G176GAT), .B(G92GAT), .ZN(n318) );
  XNOR2_X1 U361 ( .A(n319), .B(n318), .ZN(n326) );
  XOR2_X1 U362 ( .A(n320), .B(n326), .Z(n324) );
  XNOR2_X1 U363 ( .A(G36GAT), .B(G190GAT), .ZN(n321) );
  XNOR2_X1 U364 ( .A(n321), .B(G218GAT), .ZN(n351) );
  XNOR2_X1 U365 ( .A(n322), .B(n351), .ZN(n323) );
  XNOR2_X1 U366 ( .A(n324), .B(n323), .ZN(n515) );
  XOR2_X1 U367 ( .A(G99GAT), .B(G85GAT), .Z(n325) );
  XNOR2_X1 U368 ( .A(KEYINPUT74), .B(n325), .ZN(n349) );
  XNOR2_X1 U369 ( .A(n326), .B(n349), .ZN(n339) );
  XOR2_X1 U370 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n328) );
  XNOR2_X1 U371 ( .A(KEYINPUT73), .B(KEYINPUT31), .ZN(n327) );
  XNOR2_X1 U372 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U373 ( .A(KEYINPUT32), .B(G120GAT), .Z(n330) );
  NAND2_X1 U374 ( .A1(G230GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U375 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U376 ( .A(n332), .B(n331), .Z(n337) );
  XOR2_X1 U377 ( .A(KEYINPUT13), .B(KEYINPUT72), .Z(n334) );
  XNOR2_X1 U378 ( .A(G71GAT), .B(G57GAT), .ZN(n333) );
  XNOR2_X1 U379 ( .A(n334), .B(n333), .ZN(n370) );
  XNOR2_X1 U380 ( .A(G148GAT), .B(G106GAT), .ZN(n335) );
  XNOR2_X1 U381 ( .A(n335), .B(G78GAT), .ZN(n444) );
  XNOR2_X1 U382 ( .A(n370), .B(n444), .ZN(n336) );
  XNOR2_X1 U383 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U384 ( .A(n339), .B(n338), .ZN(n575) );
  INV_X1 U385 ( .A(KEYINPUT45), .ZN(n377) );
  XOR2_X1 U386 ( .A(G50GAT), .B(G162GAT), .Z(n442) );
  XOR2_X1 U387 ( .A(KEYINPUT9), .B(G106GAT), .Z(n341) );
  XNOR2_X1 U388 ( .A(G134GAT), .B(G92GAT), .ZN(n340) );
  XNOR2_X1 U389 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U390 ( .A(n442), .B(n342), .ZN(n344) );
  AND2_X1 U391 ( .A1(G232GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U392 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U393 ( .A(KEYINPUT10), .B(KEYINPUT77), .Z(n346) );
  XNOR2_X1 U394 ( .A(KEYINPUT11), .B(KEYINPUT76), .ZN(n345) );
  XOR2_X1 U395 ( .A(n346), .B(n345), .Z(n347) );
  XNOR2_X1 U396 ( .A(n348), .B(n347), .ZN(n353) );
  INV_X1 U397 ( .A(n349), .ZN(n350) );
  XNOR2_X1 U398 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U399 ( .A(n353), .B(n352), .ZN(n358) );
  XOR2_X1 U400 ( .A(KEYINPUT7), .B(KEYINPUT71), .Z(n355) );
  XNOR2_X1 U401 ( .A(G43GAT), .B(G29GAT), .ZN(n354) );
  XNOR2_X1 U402 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U403 ( .A(KEYINPUT8), .B(n356), .Z(n392) );
  INV_X1 U404 ( .A(n392), .ZN(n357) );
  XNOR2_X1 U405 ( .A(n358), .B(n357), .ZN(n472) );
  XNOR2_X1 U406 ( .A(n472), .B(KEYINPUT101), .ZN(n359) );
  XNOR2_X1 U407 ( .A(n359), .B(KEYINPUT36), .ZN(n584) );
  XOR2_X1 U408 ( .A(KEYINPUT79), .B(G78GAT), .Z(n361) );
  XNOR2_X1 U409 ( .A(G1GAT), .B(G64GAT), .ZN(n360) );
  XNOR2_X1 U410 ( .A(n361), .B(n360), .ZN(n366) );
  XOR2_X1 U411 ( .A(n362), .B(KEYINPUT15), .Z(n364) );
  NAND2_X1 U412 ( .A1(G231GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U413 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U414 ( .A(n366), .B(n365), .ZN(n375) );
  XOR2_X1 U415 ( .A(G22GAT), .B(G155GAT), .Z(n439) );
  XOR2_X1 U416 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n368) );
  XNOR2_X1 U417 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n367) );
  XNOR2_X1 U418 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U419 ( .A(n439), .B(n369), .Z(n373) );
  XNOR2_X1 U420 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U421 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U422 ( .A(n375), .B(n374), .ZN(n548) );
  NOR2_X1 U423 ( .A1(n584), .A2(n548), .ZN(n376) );
  XNOR2_X1 U424 ( .A(n377), .B(n376), .ZN(n378) );
  NOR2_X1 U425 ( .A1(n575), .A2(n378), .ZN(n399) );
  XOR2_X1 U426 ( .A(G197GAT), .B(G113GAT), .Z(n380) );
  XNOR2_X1 U427 ( .A(G1GAT), .B(G141GAT), .ZN(n379) );
  XNOR2_X1 U428 ( .A(n380), .B(n379), .ZN(n382) );
  XOR2_X1 U429 ( .A(G36GAT), .B(G50GAT), .Z(n381) );
  XNOR2_X1 U430 ( .A(n382), .B(n381), .ZN(n396) );
  XOR2_X1 U431 ( .A(G22GAT), .B(G15GAT), .Z(n384) );
  XNOR2_X1 U432 ( .A(G169GAT), .B(G8GAT), .ZN(n383) );
  XNOR2_X1 U433 ( .A(n384), .B(n383), .ZN(n388) );
  XOR2_X1 U434 ( .A(KEYINPUT70), .B(KEYINPUT67), .Z(n386) );
  XNOR2_X1 U435 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n385) );
  XNOR2_X1 U436 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U437 ( .A(n388), .B(n387), .Z(n394) );
  XOR2_X1 U438 ( .A(KEYINPUT66), .B(KEYINPUT65), .Z(n390) );
  XNOR2_X1 U439 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n389) );
  XNOR2_X1 U440 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U441 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U442 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U443 ( .A(n396), .B(n395), .ZN(n398) );
  NAND2_X1 U444 ( .A1(G229GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X2 U445 ( .A(n398), .B(n397), .ZN(n571) );
  NAND2_X1 U446 ( .A1(n399), .A2(n571), .ZN(n406) );
  XOR2_X1 U447 ( .A(KEYINPUT47), .B(KEYINPUT112), .Z(n404) );
  XNOR2_X1 U448 ( .A(KEYINPUT41), .B(n575), .ZN(n557) );
  NOR2_X1 U449 ( .A1(n571), .A2(n557), .ZN(n400) );
  XNOR2_X1 U450 ( .A(n400), .B(KEYINPUT46), .ZN(n401) );
  NOR2_X1 U451 ( .A1(n472), .A2(n401), .ZN(n402) );
  INV_X1 U452 ( .A(n548), .ZN(n579) );
  XNOR2_X1 U453 ( .A(KEYINPUT111), .B(n579), .ZN(n564) );
  NAND2_X1 U454 ( .A1(n402), .A2(n564), .ZN(n403) );
  XNOR2_X1 U455 ( .A(n404), .B(n403), .ZN(n405) );
  NAND2_X1 U456 ( .A1(n406), .A2(n405), .ZN(n407) );
  XNOR2_X1 U457 ( .A(n407), .B(KEYINPUT48), .ZN(n408) );
  XNOR2_X1 U458 ( .A(KEYINPUT113), .B(n408), .ZN(n523) );
  NOR2_X1 U459 ( .A1(n515), .A2(n523), .ZN(n409) );
  XNOR2_X1 U460 ( .A(KEYINPUT54), .B(n409), .ZN(n431) );
  XOR2_X1 U461 ( .A(G148GAT), .B(KEYINPUT94), .Z(n411) );
  XNOR2_X1 U462 ( .A(G57GAT), .B(KEYINPUT4), .ZN(n410) );
  XNOR2_X1 U463 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U464 ( .A(G127GAT), .B(n412), .Z(n414) );
  NAND2_X1 U465 ( .A1(G225GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U466 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U467 ( .A(n415), .B(KEYINPUT95), .Z(n420) );
  XOR2_X1 U468 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n417) );
  XNOR2_X1 U469 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n416) );
  XNOR2_X1 U470 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U471 ( .A(G141GAT), .B(n418), .Z(n451) );
  XNOR2_X1 U472 ( .A(n451), .B(KEYINPUT5), .ZN(n419) );
  XNOR2_X1 U473 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U474 ( .A(G162GAT), .B(G85GAT), .Z(n422) );
  XNOR2_X1 U475 ( .A(G29GAT), .B(G1GAT), .ZN(n421) );
  XNOR2_X1 U476 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U477 ( .A(n424), .B(n423), .Z(n430) );
  XOR2_X1 U478 ( .A(KEYINPUT96), .B(KEYINPUT6), .Z(n426) );
  XNOR2_X1 U479 ( .A(G155GAT), .B(KEYINPUT1), .ZN(n425) );
  XNOR2_X1 U480 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U481 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U482 ( .A(n430), .B(n429), .Z(n524) );
  AND2_X1 U483 ( .A1(n431), .A2(n524), .ZN(n432) );
  XOR2_X1 U484 ( .A(n432), .B(KEYINPUT64), .Z(n569) );
  XOR2_X1 U485 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n434) );
  NAND2_X1 U486 ( .A1(G228GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U488 ( .A(KEYINPUT22), .B(n435), .ZN(n449) );
  XOR2_X1 U489 ( .A(KEYINPUT24), .B(KEYINPUT93), .Z(n437) );
  XNOR2_X1 U490 ( .A(G218GAT), .B(G204GAT), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U492 ( .A(n438), .B(KEYINPUT23), .Z(n441) );
  XNOR2_X1 U493 ( .A(G211GAT), .B(n439), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n443) );
  XOR2_X1 U495 ( .A(n443), .B(n442), .Z(n447) );
  XNOR2_X1 U496 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U497 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U498 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U499 ( .A(n451), .B(n450), .ZN(n466) );
  NOR2_X1 U500 ( .A1(n569), .A2(n466), .ZN(n453) );
  XNOR2_X1 U501 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n452) );
  XNOR2_X1 U502 ( .A(n453), .B(n452), .ZN(n554) );
  AND2_X1 U503 ( .A1(n554), .A2(n472), .ZN(n454) );
  AND2_X1 U504 ( .A1(n555), .A2(n454), .ZN(n455) );
  XNOR2_X1 U505 ( .A(G190GAT), .B(n455), .ZN(n456) );
  XNOR2_X1 U506 ( .A(n457), .B(n456), .ZN(G1351GAT) );
  NOR2_X1 U507 ( .A1(n571), .A2(n575), .ZN(n487) );
  XNOR2_X1 U508 ( .A(n515), .B(KEYINPUT97), .ZN(n458) );
  XNOR2_X1 U509 ( .A(n458), .B(KEYINPUT27), .ZN(n525) );
  NAND2_X1 U510 ( .A1(n525), .A2(n529), .ZN(n459) );
  NOR2_X1 U511 ( .A1(n555), .A2(n459), .ZN(n460) );
  NOR2_X1 U512 ( .A1(n524), .A2(n460), .ZN(n471) );
  INV_X1 U513 ( .A(n555), .ZN(n527) );
  NAND2_X1 U514 ( .A1(n466), .A2(n527), .ZN(n461) );
  XNOR2_X1 U515 ( .A(n461), .B(KEYINPUT26), .ZN(n462) );
  XNOR2_X1 U516 ( .A(KEYINPUT98), .B(n462), .ZN(n568) );
  INV_X1 U517 ( .A(n525), .ZN(n463) );
  NOR2_X1 U518 ( .A1(n568), .A2(n463), .ZN(n541) );
  NOR2_X1 U519 ( .A1(n515), .A2(n527), .ZN(n464) );
  XOR2_X1 U520 ( .A(KEYINPUT99), .B(n464), .Z(n465) );
  NOR2_X1 U521 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U522 ( .A(n467), .B(KEYINPUT25), .ZN(n468) );
  NAND2_X1 U523 ( .A1(n468), .A2(n524), .ZN(n469) );
  NOR2_X1 U524 ( .A1(n541), .A2(n469), .ZN(n470) );
  NOR2_X1 U525 ( .A1(n471), .A2(n470), .ZN(n485) );
  XOR2_X1 U526 ( .A(KEYINPUT16), .B(KEYINPUT82), .Z(n474) );
  INV_X1 U527 ( .A(n472), .ZN(n551) );
  NAND2_X1 U528 ( .A1(n579), .A2(n551), .ZN(n473) );
  XNOR2_X1 U529 ( .A(n474), .B(n473), .ZN(n475) );
  AND2_X1 U530 ( .A1(n485), .A2(n475), .ZN(n498) );
  NAND2_X1 U531 ( .A1(n487), .A2(n498), .ZN(n482) );
  NOR2_X1 U532 ( .A1(n524), .A2(n482), .ZN(n476) );
  XOR2_X1 U533 ( .A(G1GAT), .B(n476), .Z(n477) );
  XNOR2_X1 U534 ( .A(KEYINPUT34), .B(n477), .ZN(G1324GAT) );
  NOR2_X1 U535 ( .A1(n515), .A2(n482), .ZN(n478) );
  XOR2_X1 U536 ( .A(G8GAT), .B(n478), .Z(G1325GAT) );
  NOR2_X1 U537 ( .A1(n527), .A2(n482), .ZN(n480) );
  XNOR2_X1 U538 ( .A(KEYINPUT100), .B(KEYINPUT35), .ZN(n479) );
  XNOR2_X1 U539 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U540 ( .A(G15GAT), .B(n481), .ZN(G1326GAT) );
  NOR2_X1 U541 ( .A1(n529), .A2(n482), .ZN(n483) );
  XOR2_X1 U542 ( .A(G22GAT), .B(n483), .Z(G1327GAT) );
  NOR2_X1 U543 ( .A1(n584), .A2(n579), .ZN(n484) );
  NAND2_X1 U544 ( .A1(n485), .A2(n484), .ZN(n486) );
  XNOR2_X1 U545 ( .A(KEYINPUT37), .B(n486), .ZN(n513) );
  NAND2_X1 U546 ( .A1(n513), .A2(n487), .ZN(n488) );
  XNOR2_X1 U547 ( .A(KEYINPUT38), .B(n488), .ZN(n495) );
  NOR2_X1 U548 ( .A1(n495), .A2(n524), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n489), .B(KEYINPUT39), .ZN(n490) );
  XNOR2_X1 U550 ( .A(G29GAT), .B(n490), .ZN(G1328GAT) );
  NOR2_X1 U551 ( .A1(n515), .A2(n495), .ZN(n491) );
  XOR2_X1 U552 ( .A(KEYINPUT102), .B(n491), .Z(n492) );
  XNOR2_X1 U553 ( .A(G36GAT), .B(n492), .ZN(G1329GAT) );
  NOR2_X1 U554 ( .A1(n495), .A2(n527), .ZN(n493) );
  XOR2_X1 U555 ( .A(KEYINPUT40), .B(n493), .Z(n494) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  NOR2_X1 U557 ( .A1(n495), .A2(n529), .ZN(n496) );
  XOR2_X1 U558 ( .A(G50GAT), .B(n496), .Z(G1331GAT) );
  INV_X1 U559 ( .A(n571), .ZN(n497) );
  NOR2_X1 U560 ( .A1(n557), .A2(n497), .ZN(n512) );
  NAND2_X1 U561 ( .A1(n512), .A2(n498), .ZN(n506) );
  NOR2_X1 U562 ( .A1(n524), .A2(n506), .ZN(n500) );
  XNOR2_X1 U563 ( .A(KEYINPUT103), .B(KEYINPUT42), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(n501), .ZN(G1332GAT) );
  NOR2_X1 U566 ( .A1(n515), .A2(n506), .ZN(n502) );
  XOR2_X1 U567 ( .A(KEYINPUT104), .B(n502), .Z(n503) );
  XNOR2_X1 U568 ( .A(G64GAT), .B(n503), .ZN(G1333GAT) );
  NOR2_X1 U569 ( .A1(n527), .A2(n506), .ZN(n505) );
  XNOR2_X1 U570 ( .A(G71GAT), .B(KEYINPUT105), .ZN(n504) );
  XNOR2_X1 U571 ( .A(n505), .B(n504), .ZN(G1334GAT) );
  NOR2_X1 U572 ( .A1(n529), .A2(n506), .ZN(n511) );
  XOR2_X1 U573 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n508) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U576 ( .A(KEYINPUT106), .B(n509), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  NAND2_X1 U578 ( .A1(n513), .A2(n512), .ZN(n520) );
  NOR2_X1 U579 ( .A1(n524), .A2(n520), .ZN(n514) );
  XOR2_X1 U580 ( .A(G85GAT), .B(n514), .Z(G1336GAT) );
  NOR2_X1 U581 ( .A1(n515), .A2(n520), .ZN(n516) );
  XOR2_X1 U582 ( .A(G92GAT), .B(n516), .Z(G1337GAT) );
  NOR2_X1 U583 ( .A1(n527), .A2(n520), .ZN(n517) );
  XOR2_X1 U584 ( .A(G99GAT), .B(n517), .Z(G1338GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n519) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n518) );
  XNOR2_X1 U587 ( .A(n519), .B(n518), .ZN(n522) );
  NOR2_X1 U588 ( .A1(n529), .A2(n520), .ZN(n521) );
  XOR2_X1 U589 ( .A(n522), .B(n521), .Z(G1339GAT) );
  NOR2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n542) );
  NAND2_X1 U591 ( .A1(n525), .A2(n542), .ZN(n526) );
  NOR2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n528), .B(KEYINPUT114), .ZN(n530) );
  NAND2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n537) );
  NOR2_X1 U595 ( .A1(n571), .A2(n537), .ZN(n532) );
  XNOR2_X1 U596 ( .A(G113GAT), .B(KEYINPUT115), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(G1340GAT) );
  NOR2_X1 U598 ( .A1(n557), .A2(n537), .ZN(n534) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(G1341GAT) );
  NOR2_X1 U601 ( .A1(n564), .A2(n537), .ZN(n535) );
  XOR2_X1 U602 ( .A(KEYINPUT50), .B(n535), .Z(n536) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  NOR2_X1 U604 ( .A1(n551), .A2(n537), .ZN(n539) );
  XNOR2_X1 U605 ( .A(KEYINPUT116), .B(KEYINPUT51), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U607 ( .A(G134GAT), .B(n540), .ZN(G1343GAT) );
  NAND2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n550) );
  NOR2_X1 U609 ( .A1(n571), .A2(n550), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(G1344GAT) );
  NOR2_X1 U612 ( .A1(n557), .A2(n550), .ZN(n546) );
  XNOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(n547), .ZN(G1345GAT) );
  NOR2_X1 U616 ( .A1(n548), .A2(n550), .ZN(n549) );
  XOR2_X1 U617 ( .A(G155GAT), .B(n549), .Z(G1346GAT) );
  NOR2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U619 ( .A(KEYINPUT118), .B(n552), .Z(n553) );
  XNOR2_X1 U620 ( .A(G162GAT), .B(n553), .ZN(G1347GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n563) );
  NOR2_X1 U622 ( .A1(n563), .A2(n571), .ZN(n556) );
  XOR2_X1 U623 ( .A(G169GAT), .B(n556), .Z(G1348GAT) );
  NOR2_X1 U624 ( .A1(n557), .A2(n563), .ZN(n562) );
  XOR2_X1 U625 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n559) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U628 ( .A(KEYINPUT56), .B(n560), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1349GAT) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n566) );
  XNOR2_X1 U631 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n573) );
  OR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(KEYINPUT124), .ZN(n583) );
  NOR2_X1 U637 ( .A1(n571), .A2(n583), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n577) );
  INV_X1 U641 ( .A(n583), .ZN(n580) );
  NAND2_X1 U642 ( .A1(n580), .A2(n575), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XOR2_X1 U644 ( .A(G204GAT), .B(n578), .Z(G1353GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(KEYINPUT126), .ZN(n582) );
  XNOR2_X1 U647 ( .A(G211GAT), .B(n582), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(n585), .Z(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

