//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n591, new_n592, new_n593, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n630,
    new_n633, new_n635, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1174, new_n1175, new_n1176;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT67), .Z(G319));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT68), .B(G2105), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n462), .A2(G137), .A3(new_n464), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n465), .A2(new_n469), .ZN(G160));
  NAND2_X1  g045(.A1(new_n459), .A2(new_n461), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(new_n464), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n471), .A2(G2105), .ZN(new_n473));
  AOI22_X1  g048(.A1(G124), .A2(new_n472), .B1(new_n473), .B2(G136), .ZN(new_n474));
  NOR2_X1   g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT69), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G162));
  NAND3_X1  g054(.A1(new_n462), .A2(G138), .A3(new_n464), .ZN(new_n480));
  NAND2_X1  g055(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n462), .A2(new_n464), .A3(G138), .A4(new_n481), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT70), .B1(new_n467), .B2(G114), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n487), .A2(new_n488), .A3(G2105), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n486), .A2(new_n489), .A3(G2104), .A4(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n459), .A2(new_n461), .A3(G126), .A4(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n491), .A2(new_n492), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT71), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n485), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT73), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT73), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT75), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT75), .A3(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G62), .ZN(new_n511));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n504), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT74), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n500), .A2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT73), .B(G651), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  OAI211_X1 g093(.A(G543), .B(new_n516), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n514), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n515), .B1(new_n504), .B2(KEYINPUT6), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n522), .A2(KEYINPUT74), .A3(G50), .A4(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n518), .B1(new_n501), .B2(new_n503), .ZN(new_n525));
  NOR3_X1   g100(.A1(new_n525), .A2(new_n509), .A3(new_n515), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G88), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT76), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT76), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n524), .A2(new_n530), .A3(new_n527), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n513), .B1(new_n529), .B2(new_n531), .ZN(G166));
  INV_X1    g107(.A(KEYINPUT77), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n509), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT77), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n536), .A2(G63), .A3(G651), .ZN(new_n537));
  INV_X1    g112(.A(new_n519), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G51), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n526), .A2(G89), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT7), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n537), .A2(new_n539), .A3(new_n540), .A4(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  AOI22_X1  g119(.A1(new_n536), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n504), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n526), .A2(G90), .ZN(new_n547));
  INV_X1    g122(.A(G52), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n548), .B2(new_n519), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(G171));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n551), .B1(new_n534), .B2(new_n535), .ZN(new_n552));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT78), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT78), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT77), .ZN(new_n557));
  AOI21_X1  g132(.A(KEYINPUT77), .B1(new_n506), .B2(new_n508), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g134(.A(new_n556), .B(new_n553), .C1(new_n559), .C2(new_n551), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n555), .A2(new_n560), .A3(new_n517), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT79), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT79), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n555), .A2(new_n560), .A3(new_n563), .A4(new_n517), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g140(.A(KEYINPUT80), .B(G43), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n538), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n526), .A2(G81), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G860), .ZN(G153));
  AND3_X1   g146(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G36), .ZN(G176));
  NAND2_X1  g148(.A1(G1), .A2(G3), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT8), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n572), .A2(new_n575), .ZN(G188));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  INV_X1    g152(.A(G53), .ZN(new_n578));
  OAI211_X1 g153(.A(KEYINPUT81), .B(new_n577), .C1(new_n519), .C2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n526), .A2(G91), .ZN(new_n580));
  NAND2_X1  g155(.A1(G78), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G65), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n509), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G651), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n579), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  OR3_X1    g160(.A1(new_n519), .A2(KEYINPUT81), .A3(new_n578), .ZN(new_n586));
  OAI21_X1  g161(.A(KEYINPUT81), .B1(new_n519), .B2(new_n578), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n586), .A2(KEYINPUT9), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n585), .A2(new_n588), .ZN(G299));
  INV_X1    g164(.A(G171), .ZN(G301));
  INV_X1    g165(.A(new_n513), .ZN(new_n591));
  AOI221_X4 g166(.A(KEYINPUT76), .B1(new_n526), .B2(G88), .C1(new_n521), .C2(new_n523), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n530), .B1(new_n524), .B2(new_n527), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(G303));
  OAI21_X1  g169(.A(G651), .B1(new_n536), .B2(G74), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n538), .A2(G49), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n526), .A2(G87), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G288));
  INV_X1    g173(.A(G543), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n522), .A2(G48), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n517), .A2(G73), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n522), .A2(G86), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n517), .A2(G61), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n509), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n602), .A2(new_n605), .ZN(G305));
  AOI22_X1  g181(.A1(new_n536), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(new_n504), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n526), .A2(G85), .ZN(new_n609));
  INV_X1    g184(.A(G47), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n519), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(G290));
  NAND2_X1  g188(.A1(G301), .A2(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n526), .A2(G92), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n538), .A2(G54), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT82), .B(G66), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n509), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G651), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n617), .A2(new_n618), .A3(new_n622), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n623), .A2(KEYINPUT83), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(KEYINPUT83), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n614), .B1(new_n626), .B2(G868), .ZN(G284));
  XNOR2_X1  g202(.A(G284), .B(KEYINPUT84), .ZN(G321));
  NAND2_X1  g203(.A1(G286), .A2(G868), .ZN(new_n629));
  AND2_X1   g204(.A1(new_n585), .A2(new_n588), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G868), .ZN(G297));
  OAI21_X1  g206(.A(new_n629), .B1(new_n630), .B2(G868), .ZN(G280));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n626), .B1(new_n633), .B2(G860), .ZN(G148));
  INV_X1    g209(.A(G868), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n569), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(G559), .B1(new_n624), .B2(new_n625), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n636), .B1(new_n637), .B2(new_n635), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(KEYINPUT85), .A2(G2100), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT12), .Z(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT13), .Z(new_n643));
  NOR2_X1   g218(.A1(KEYINPUT85), .A2(G2100), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n640), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n472), .A2(G123), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n473), .A2(G135), .ZN(new_n647));
  OAI221_X1 g222(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n464), .C2(G111), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT86), .B(G2096), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n645), .B(new_n651), .C1(new_n643), .C2(new_n640), .ZN(G156));
  XNOR2_X1  g227(.A(G2427), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2430), .ZN(new_n654));
  XOR2_X1   g229(.A(KEYINPUT15), .B(G2435), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT14), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2446), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT16), .B(G2443), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n658), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT87), .B(G1341), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(G14), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT88), .ZN(G401));
  XOR2_X1   g242(.A(G2067), .B(G2678), .Z(new_n668));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT89), .B(KEYINPUT17), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  AND2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n672), .B1(new_n668), .B2(new_n669), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n668), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n671), .A2(new_n674), .ZN(new_n676));
  INV_X1    g251(.A(new_n668), .ZN(new_n677));
  INV_X1    g252(.A(new_n669), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n677), .A2(new_n678), .A3(new_n672), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT18), .Z(new_n680));
  NAND3_X1  g255(.A1(new_n675), .A2(new_n676), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G2096), .B(G2100), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G227));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n687), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n692));
  AOI21_X1  g267(.A(new_n689), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n685), .A2(new_n688), .A3(new_n690), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n693), .B(new_n694), .C1(new_n691), .C2(new_n692), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT92), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT91), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n698));
  XNOR2_X1  g273(.A(G1981), .B(G1986), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(G1991), .B(G1996), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n697), .B(new_n702), .ZN(G229));
  INV_X1    g278(.A(KEYINPUT34), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G6), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n602), .A2(new_n605), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(new_n705), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT32), .B(G1981), .Z(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n709), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n711), .B(new_n706), .C1(new_n707), .C2(new_n705), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n705), .A2(G22), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G303), .B2(G16), .ZN(new_n716));
  INV_X1    g291(.A(G1971), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n713), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n717), .B(new_n714), .C1(G166), .C2(new_n705), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(KEYINPUT94), .B1(G16), .B2(G23), .ZN(new_n722));
  OR3_X1    g297(.A1(KEYINPUT94), .A2(G16), .A3(G23), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n722), .B(new_n723), .C1(G288), .C2(new_n705), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT95), .B(KEYINPUT33), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1976), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n724), .B(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(KEYINPUT96), .B1(new_n721), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n714), .B1(G166), .B2(new_n705), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G1971), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n730), .A2(new_n727), .A3(new_n719), .A4(new_n713), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT96), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n704), .B1(new_n728), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n705), .A2(G24), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n612), .B2(new_n705), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(G1986), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n731), .A2(new_n732), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n729), .A2(G1971), .B1(new_n710), .B2(new_n712), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n739), .A2(KEYINPUT96), .A3(new_n727), .A4(new_n719), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n738), .A2(KEYINPUT34), .A3(new_n740), .ZN(new_n741));
  AOI22_X1  g316(.A1(G119), .A2(new_n472), .B1(new_n473), .B2(G131), .ZN(new_n742));
  OAI221_X1 g317(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n464), .C2(G107), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  MUX2_X1   g319(.A(G25), .B(new_n744), .S(G29), .Z(new_n745));
  XOR2_X1   g320(.A(KEYINPUT35), .B(G1991), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT93), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n745), .B(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n736), .B2(G1986), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n734), .A2(new_n737), .A3(new_n741), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(KEYINPUT36), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n741), .A2(new_n749), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT36), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n752), .A2(new_n753), .A3(new_n737), .A4(new_n734), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G29), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n756), .A2(G33), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT25), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G139), .B2(new_n473), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n464), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n757), .B1(new_n762), .B2(G29), .ZN(new_n763));
  INV_X1    g338(.A(G2072), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n756), .A2(G35), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G162), .B2(new_n756), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n767), .A2(KEYINPUT29), .ZN(new_n768));
  INV_X1    g343(.A(G2090), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(KEYINPUT29), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT28), .ZN(new_n772));
  INV_X1    g347(.A(G26), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(G29), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(G29), .ZN(new_n775));
  AOI22_X1  g350(.A1(G128), .A2(new_n472), .B1(new_n473), .B2(G140), .ZN(new_n776));
  OAI221_X1 g351(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n464), .C2(G116), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n775), .B1(new_n778), .B2(G29), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n774), .B1(new_n779), .B2(new_n772), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(G2067), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n771), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n756), .A2(G32), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n472), .A2(G129), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n473), .A2(G141), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n467), .A2(G105), .A3(G2104), .ZN(new_n786));
  NAND3_X1  g361(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT26), .Z(new_n788));
  NAND4_X1  g363(.A1(new_n784), .A2(new_n785), .A3(new_n786), .A4(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n783), .B1(new_n790), .B2(new_n756), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT98), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT27), .B(G1996), .Z(new_n793));
  NOR2_X1   g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n780), .A2(G2067), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(G29), .B1(new_n465), .B2(new_n469), .ZN(new_n797));
  OR2_X1    g372(.A1(KEYINPUT24), .A2(G34), .ZN(new_n798));
  NAND2_X1  g373(.A1(KEYINPUT24), .A2(G34), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n798), .A2(new_n756), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n801), .A2(KEYINPUT97), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(KEYINPUT97), .ZN(new_n803));
  INV_X1    g378(.A(G2084), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NOR4_X1   g380(.A1(new_n782), .A2(new_n794), .A3(new_n796), .A4(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(G1961), .ZN(new_n807));
  NOR2_X1   g382(.A1(G301), .A2(new_n705), .ZN(new_n808));
  NOR2_X1   g383(.A1(G5), .A2(G16), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n792), .A2(new_n793), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n804), .B1(new_n802), .B2(new_n803), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(KEYINPUT101), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n756), .A2(G27), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G164), .B2(new_n756), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G2078), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n769), .B1(new_n768), .B2(new_n770), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n763), .A2(new_n764), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT101), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n810), .A2(new_n811), .A3(new_n821), .A4(new_n812), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n806), .A2(new_n814), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(G4), .A2(G16), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n626), .B2(G16), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1348), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n705), .A2(G20), .ZN(new_n828));
  OAI211_X1 g403(.A(KEYINPUT23), .B(new_n828), .C1(new_n630), .C2(new_n705), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(KEYINPUT23), .B2(new_n828), .ZN(new_n830));
  INV_X1    g405(.A(G1956), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(G16), .A2(G21), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(G168), .B2(G16), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT99), .B(G1966), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n649), .ZN(new_n837));
  INV_X1    g412(.A(G28), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n838), .A2(KEYINPUT30), .ZN(new_n839));
  AOI21_X1  g414(.A(G29), .B1(new_n838), .B2(KEYINPUT30), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n837), .A2(G29), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n836), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(KEYINPUT31), .B(G11), .ZN(new_n843));
  OR3_X1    g418(.A1(new_n808), .A2(new_n807), .A3(new_n809), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(KEYINPUT100), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n842), .A2(new_n847), .A3(new_n843), .A4(new_n844), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n832), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n705), .A2(G19), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n570), .B2(new_n705), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(G1341), .Z(new_n852));
  AND4_X1   g427(.A1(new_n765), .A2(new_n827), .A3(new_n849), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n755), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(G311));
  INV_X1    g430(.A(KEYINPUT102), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n755), .A2(new_n853), .A3(KEYINPUT102), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(G150));
  AOI22_X1  g434(.A1(new_n536), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(new_n504), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n538), .A2(G55), .ZN(new_n862));
  INV_X1    g437(.A(new_n526), .ZN(new_n863));
  INV_X1    g438(.A(G93), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(G860), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT37), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n569), .A2(new_n866), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n562), .A2(new_n564), .B1(G81), .B2(new_n526), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n871), .A2(new_n567), .A3(new_n867), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n873), .B(new_n874), .Z(new_n875));
  NAND2_X1  g450(.A1(new_n626), .A2(G559), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT39), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n875), .B(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n869), .B1(new_n878), .B2(G860), .ZN(G145));
  XNOR2_X1  g454(.A(G160), .B(new_n837), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n744), .B(new_n789), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(new_n882));
  AOI22_X1  g457(.A1(G130), .A2(new_n472), .B1(new_n473), .B2(G142), .ZN(new_n883));
  OAI21_X1  g458(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n884), .A2(KEYINPUT104), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(KEYINPUT104), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n885), .B(new_n886), .C1(G118), .C2(new_n464), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n478), .B(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n882), .B(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n762), .B(new_n778), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n485), .A2(new_n496), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n642), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n891), .B(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n890), .B(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(G37), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g473(.A1(new_n626), .A2(new_n633), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n873), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n637), .A2(new_n872), .A3(new_n870), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n623), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n630), .A2(KEYINPUT105), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n905));
  NAND2_X1  g480(.A1(G299), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n623), .A2(new_n905), .A3(G299), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT106), .B1(new_n902), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(KEYINPUT41), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n902), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT106), .ZN(new_n913));
  INV_X1    g488(.A(new_n909), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n900), .A2(new_n901), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n910), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT42), .ZN(new_n917));
  XNOR2_X1  g492(.A(G303), .B(G288), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(G305), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(G290), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n918), .A2(G305), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(G305), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n612), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n910), .A2(new_n925), .A3(new_n912), .A4(new_n915), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n917), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n924), .B1(new_n917), .B2(new_n926), .ZN(new_n928));
  OAI21_X1  g503(.A(G868), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n867), .A2(new_n635), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(G295));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n930), .ZN(G331));
  INV_X1    g507(.A(new_n923), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n612), .B1(new_n921), .B2(new_n922), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AND4_X1   g510(.A1(new_n567), .A2(new_n565), .A3(new_n568), .A4(new_n867), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n867), .B1(new_n871), .B2(new_n567), .ZN(new_n937));
  OAI21_X1  g512(.A(G171), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n870), .A2(G301), .A3(new_n872), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n938), .A2(G168), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(G168), .B1(new_n938), .B2(new_n939), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n940), .A2(new_n941), .A3(new_n909), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT41), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n909), .B(new_n943), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n936), .A2(new_n937), .A3(G171), .ZN(new_n945));
  AOI21_X1  g520(.A(G301), .B1(new_n870), .B2(new_n872), .ZN(new_n946));
  OAI21_X1  g521(.A(G286), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n938), .A2(G168), .A3(new_n939), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n935), .B1(new_n942), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n911), .B1(new_n940), .B2(new_n941), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n947), .A2(new_n914), .A3(new_n948), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n924), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(new_n896), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n950), .A2(new_n896), .A3(new_n955), .A4(new_n953), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(KEYINPUT44), .A3(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n954), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n950), .A2(KEYINPUT43), .A3(new_n896), .A4(new_n953), .ZN(new_n962));
  XOR2_X1   g537(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n959), .A2(new_n964), .ZN(G397));
  AOI21_X1  g540(.A(new_n493), .B1(new_n483), .B2(new_n484), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n966), .A2(G1384), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n967), .A2(KEYINPUT45), .ZN(new_n968));
  NAND2_X1  g543(.A1(G160), .A2(G40), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n971), .B(KEYINPUT110), .Z(new_n972));
  INV_X1    g547(.A(G2067), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n778), .B(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G1996), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n974), .B1(new_n975), .B2(new_n790), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n971), .A2(G1996), .ZN(new_n977));
  AOI22_X1  g552(.A1(new_n972), .A2(new_n976), .B1(new_n790), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n972), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n744), .B(new_n747), .Z(new_n980));
  OAI21_X1  g555(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OR3_X1    g556(.A1(new_n971), .A2(G290), .A3(G1986), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n968), .A2(G1986), .A3(new_n970), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n982), .B1(new_n612), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT109), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT53), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n966), .A2(new_n988), .A3(G1384), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n493), .B(KEYINPUT71), .ZN(new_n991));
  AOI21_X1  g566(.A(G1384), .B1(new_n991), .B2(new_n485), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n990), .B(new_n970), .C1(KEYINPUT45), .C2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n987), .B1(new_n993), .B2(G2078), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT50), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT111), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n969), .B1(new_n995), .B2(new_n967), .ZN(new_n997));
  INV_X1    g572(.A(G1384), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n498), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(new_n1000), .A3(KEYINPUT50), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n996), .A2(new_n997), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n807), .ZN(new_n1003));
  INV_X1    g578(.A(G2078), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n990), .A2(KEYINPUT53), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n970), .B1(KEYINPUT45), .B2(new_n967), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n994), .A2(new_n1003), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(G171), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n999), .A2(new_n988), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1011), .A2(KEYINPUT53), .A3(new_n1004), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1012), .A2(new_n1003), .A3(new_n994), .A4(G301), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1009), .A2(KEYINPUT54), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT126), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT126), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1009), .A2(new_n1016), .A3(KEYINPUT54), .A4(new_n1013), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n993), .A2(new_n717), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT112), .B(G2090), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n996), .A2(new_n997), .A3(new_n1001), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G303), .A2(G8), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1019), .A2(new_n1022), .A3(KEYINPUT113), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1025), .A2(new_n1028), .A3(G8), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n892), .A2(new_n998), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(new_n969), .ZN(new_n1032));
  INV_X1    g607(.A(G8), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G305), .A2(G1981), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n602), .A2(new_n605), .A3(G1981), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n1037), .A3(KEYINPUT49), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT49), .ZN(new_n1039));
  INV_X1    g614(.A(G1981), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n707), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1039), .B1(new_n1041), .B2(new_n1036), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1034), .A2(new_n1038), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G288), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1045), .A2(G1976), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1046), .B(G8), .C1(new_n1031), .C2(new_n969), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1045), .A2(G1976), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1049), .A2(KEYINPUT114), .A3(new_n1034), .A4(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1034), .A2(KEYINPUT114), .A3(new_n1050), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1052), .A2(new_n1048), .A3(new_n1047), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1044), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1026), .B(KEYINPUT55), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n498), .A2(new_n995), .A3(new_n998), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n970), .B(new_n1056), .C1(new_n995), .C2(new_n967), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1058), .A2(new_n1021), .B1(new_n993), .B2(new_n717), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1055), .B1(new_n1059), .B2(new_n1033), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1030), .A2(new_n1054), .A3(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1012), .A2(new_n994), .A3(new_n1003), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(G171), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n994), .A2(new_n1003), .A3(new_n1007), .A4(G301), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT54), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1061), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n835), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n996), .A2(new_n997), .A3(new_n1001), .A4(new_n804), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1033), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT51), .B1(new_n1069), .B2(KEYINPUT125), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1067), .A2(new_n1068), .A3(G168), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1071), .A2(G8), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(G8), .ZN(new_n1074));
  AOI21_X1  g649(.A(G168), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1073), .B1(new_n1076), .B2(new_n1070), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1018), .A2(new_n1066), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G1348), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1002), .A2(new_n1079), .B1(new_n973), .B2(new_n1032), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT60), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT124), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(new_n1082), .A3(new_n623), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1080), .A2(KEYINPUT60), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n903), .A2(KEYINPUT124), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n623), .A2(new_n1082), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1080), .A2(KEYINPUT60), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1083), .A2(new_n1084), .A3(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n630), .A2(KEYINPUT116), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT117), .B1(G299), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(G299), .A2(new_n1092), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT57), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT45), .B1(new_n498), .B2(new_n998), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1098), .A2(new_n969), .A3(new_n989), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n1100), .B(KEYINPUT118), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1099), .A2(new_n1101), .B1(new_n1057), .B2(new_n831), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1091), .A2(KEYINPUT57), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1097), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1102), .B1(new_n1097), .B2(new_n1103), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1089), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n1088), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1097), .A2(new_n1103), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1102), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1111), .A2(KEYINPUT61), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1104), .A2(KEYINPUT122), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1097), .A2(new_n1102), .A3(new_n1114), .A4(new_n1103), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1112), .A2(new_n1113), .A3(KEYINPUT123), .A4(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1113), .A2(new_n1111), .A3(KEYINPUT61), .A4(new_n1115), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT58), .B(G1341), .ZN(new_n1120));
  OAI22_X1  g695(.A1(new_n993), .A2(G1996), .B1(new_n1032), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n570), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1123), .A2(KEYINPUT120), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1122), .B(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1108), .A2(new_n1116), .A3(new_n1119), .A4(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1111), .B1(new_n623), .B2(new_n1080), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1127), .A2(new_n1128), .A3(new_n1104), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1128), .B1(new_n1127), .B2(new_n1104), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1078), .B1(new_n1126), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(G1976), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1043), .A2(new_n1134), .A3(new_n1045), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1037), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT115), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT115), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1135), .A2(new_n1138), .A3(new_n1037), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1137), .A2(new_n1034), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1054), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1140), .B1(new_n1141), .B2(new_n1030), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT63), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1069), .A2(G168), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1143), .B1(new_n1061), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1025), .A2(G8), .A3(new_n1029), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1143), .B1(new_n1146), .B2(new_n1055), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1144), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1147), .A2(new_n1030), .A3(new_n1054), .A4(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1142), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1077), .A2(KEYINPUT62), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1061), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1063), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1073), .B(new_n1154), .C1(new_n1076), .C2(new_n1070), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .A4(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1150), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n986), .B1(new_n1133), .B2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n778), .A2(G2067), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n744), .A2(new_n747), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1159), .B1(new_n978), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1161), .A2(new_n979), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1162), .B(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n977), .B(KEYINPUT46), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n974), .A2(new_n790), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1165), .B1(new_n972), .B2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT47), .ZN(new_n1168));
  XOR2_X1   g743(.A(new_n982), .B(KEYINPUT48), .Z(new_n1169));
  NOR2_X1   g744(.A1(new_n981), .A2(new_n1169), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1164), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1158), .A2(new_n1171), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g747(.A1(G229), .A2(G227), .ZN(new_n1174));
  NOR2_X1   g748(.A1(G401), .A2(new_n1174), .ZN(new_n1175));
  AND2_X1   g749(.A1(new_n897), .A2(new_n456), .ZN(new_n1176));
  NAND4_X1  g750(.A1(new_n961), .A2(new_n1175), .A3(new_n962), .A4(new_n1176), .ZN(G225));
  INV_X1    g751(.A(G225), .ZN(G308));
endmodule


