//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n444, new_n445, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  XNOR2_X1  g012(.A(KEYINPUT67), .B(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XNOR2_X1  g015(.A(KEYINPUT68), .B(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  INV_X1    g017(.A(G2072), .ZN(new_n443));
  INV_X1    g018(.A(G2078), .ZN(new_n444));
  NOR2_X1   g019(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g020(.A1(new_n445), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT69), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(G113), .A3(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(G2105), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  AND3_X1   g051(.A1(new_n476), .A2(G101), .A3(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G137), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n478), .A2(G136), .ZN(new_n485));
  XOR2_X1   g060(.A(new_n485), .B(KEYINPUT70), .Z(new_n486));
  AOI21_X1  g061(.A(new_n476), .B1(new_n467), .B2(new_n468), .ZN(new_n487));
  AOI211_X1 g062(.A(new_n484), .B(new_n486), .C1(G124), .C2(new_n487), .ZN(G162));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G114), .C2(new_n476), .ZN(new_n490));
  AND2_X1   g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  NOR2_X1   g066(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n492));
  OAI211_X1 g067(.A(G126), .B(G2105), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n476), .C1(new_n491), .C2(new_n492), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT3), .B(G2104), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n497), .A2(new_n498), .A3(G138), .A4(new_n476), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(new_n496), .B2(new_n499), .ZN(G164));
  NAND2_X1  g075(.A1(G75), .A2(G543), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G62), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n508), .A2(new_n509), .B1(new_n502), .B2(new_n503), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G88), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n516), .A2(new_n517), .A3(G50), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n517), .B1(new_n516), .B2(G50), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n507), .B(new_n512), .C1(new_n518), .C2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n514), .A2(new_n515), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G543), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT72), .B(G51), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n524), .A2(G89), .ZN(new_n528));
  NAND2_X1  g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n504), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OR3_X1    g105(.A1(new_n527), .A2(new_n530), .A3(KEYINPUT73), .ZN(new_n531));
  OAI21_X1  g106(.A(KEYINPUT73), .B1(new_n527), .B2(new_n530), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(G168));
  XNOR2_X1  g108(.A(KEYINPUT5), .B(G543), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n534), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G651), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n511), .A2(G90), .B1(G52), .B2(new_n516), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT74), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(G171));
  AOI22_X1  g118(.A1(new_n534), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n536), .ZN(new_n545));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n525), .A2(new_n546), .B1(new_n510), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n504), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  INV_X1    g133(.A(G91), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n516), .A2(G53), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(KEYINPUT9), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(new_n516), .B2(G53), .ZN(new_n563));
  OAI221_X1 g138(.A(new_n558), .B1(new_n559), .B2(new_n510), .C1(new_n561), .C2(new_n563), .ZN(G299));
  INV_X1    g139(.A(G171), .ZN(G301));
  INV_X1    g140(.A(G168), .ZN(G286));
  OR2_X1    g141(.A1(new_n534), .A2(G74), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n567), .A2(G651), .B1(new_n516), .B2(G49), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n511), .A2(G87), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(KEYINPUT75), .B1(new_n511), .B2(G87), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n568), .B1(new_n571), .B2(new_n572), .ZN(G288));
  OAI21_X1  g148(.A(G61), .B1(new_n502), .B2(new_n503), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n536), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT76), .ZN(new_n577));
  OAI211_X1 g152(.A(G48), .B(G543), .C1(new_n509), .C2(new_n508), .ZN(new_n578));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n510), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n534), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n536), .ZN(new_n584));
  INV_X1    g159(.A(G47), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n525), .A2(new_n585), .B1(new_n510), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G290));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n590));
  INV_X1    g165(.A(G92), .ZN(new_n591));
  OAI21_X1  g166(.A(KEYINPUT77), .B1(new_n510), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  NOR3_X1   g168(.A1(new_n510), .A2(KEYINPUT77), .A3(new_n591), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n590), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OR3_X1    g170(.A1(new_n510), .A2(KEYINPUT77), .A3(new_n591), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n596), .A2(KEYINPUT10), .A3(new_n592), .ZN(new_n597));
  INV_X1    g172(.A(G54), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n598), .B1(new_n525), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n516), .A2(KEYINPUT78), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n504), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n600), .A2(new_n601), .B1(G651), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n595), .A2(new_n597), .A3(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n607), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g183(.A(new_n607), .B1(G868), .B2(G171), .ZN(G321));
  NOR2_X1   g184(.A1(G299), .A2(G868), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g186(.A(new_n610), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g187(.A(G860), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n606), .B1(G559), .B2(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT79), .Z(G148));
  INV_X1    g190(.A(new_n549), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n606), .A2(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n617), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g196(.A1(new_n466), .A2(G2105), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n497), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2100), .ZN(new_n627));
  AOI22_X1  g202(.A1(G123), .A2(new_n487), .B1(new_n478), .B2(G135), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  INV_X1    g204(.A(G111), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n629), .A2(KEYINPUT81), .B1(new_n630), .B2(G2105), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(KEYINPUT81), .B2(new_n629), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(KEYINPUT82), .B(G2096), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n627), .A2(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT83), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2427), .B(G2430), .Z(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n643), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(new_n651), .A3(G14), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT84), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT85), .ZN(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  XNOR2_X1  g232(.A(G2084), .B(G2090), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT18), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n657), .B(KEYINPUT17), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n661), .B(new_n658), .C1(new_n656), .C2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n658), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n656), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n660), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2096), .B(G2100), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1956), .B(G2474), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1961), .B(G1966), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT20), .ZN(new_n676));
  INV_X1    g251(.A(new_n671), .ZN(new_n677));
  INV_X1    g252(.A(new_n674), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n672), .A2(new_n673), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n676), .B(new_n680), .C1(new_n677), .C2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT87), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT88), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n683), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G229));
  MUX2_X1   g265(.A(G6), .B(G305), .S(G16), .Z(new_n691));
  XOR2_X1   g266(.A(KEYINPUT32), .B(G1981), .Z(new_n692));
  XOR2_X1   g267(.A(new_n691), .B(new_n692), .Z(new_n693));
  MUX2_X1   g268(.A(G23), .B(G288), .S(G16), .Z(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT33), .B(G1976), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n694), .B(new_n695), .Z(new_n696));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G22), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT91), .Z(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G166), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G1971), .ZN(new_n701));
  NOR3_X1   g276(.A1(new_n693), .A2(new_n696), .A3(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT34), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G25), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT89), .Z(new_n708));
  OR2_X1    g283(.A1(G95), .A2(G2105), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n709), .B(G2104), .C1(G107), .C2(new_n476), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT90), .ZN(new_n711));
  AOI22_X1  g286(.A1(G119), .A2(new_n487), .B1(new_n478), .B2(G131), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n708), .B1(new_n713), .B2(G29), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT35), .B(G1991), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n697), .A2(G24), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(new_n588), .B2(new_n697), .ZN(new_n718));
  INV_X1    g293(.A(G1986), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n704), .A2(new_n705), .A3(new_n716), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n706), .A2(G35), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G162), .B2(new_n706), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT29), .B(G2090), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT95), .B(KEYINPUT24), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G34), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(new_n706), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n480), .B2(new_n706), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G2084), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT100), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT30), .B(G28), .ZN(new_n736));
  OR2_X1    g311(.A1(KEYINPUT31), .A2(G11), .ZN(new_n737));
  NAND2_X1  g312(.A1(KEYINPUT31), .A2(G11), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n736), .A2(new_n706), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n633), .B2(new_n706), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT25), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n478), .A2(G139), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n497), .A2(G127), .ZN(new_n745));
  NAND2_X1  g320(.A1(G115), .A2(G2104), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n476), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(new_n706), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n706), .B2(G33), .ZN(new_n750));
  OAI221_X1 g325(.A(new_n734), .B1(new_n735), .B2(new_n740), .C1(new_n750), .C2(new_n443), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n443), .ZN(new_n752));
  NOR2_X1   g327(.A1(G164), .A2(new_n706), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G27), .B2(new_n706), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(new_n444), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n754), .A2(new_n444), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n740), .A2(new_n735), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n752), .A2(new_n755), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  NOR3_X1   g333(.A1(new_n729), .A2(new_n751), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n706), .A2(G26), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT28), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n478), .A2(G140), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n487), .A2(G128), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n476), .A2(G116), .ZN(new_n764));
  OAI21_X1  g339(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n762), .B(new_n763), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT94), .Z(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n761), .B1(new_n768), .B2(G29), .ZN(new_n769));
  INV_X1    g344(.A(G2067), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(G16), .A2(G19), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n549), .B2(G16), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT93), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G1341), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G4), .A2(G16), .ZN(new_n777));
  INV_X1    g352(.A(new_n606), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(G16), .ZN(new_n779));
  INV_X1    g354(.A(G1348), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n697), .A2(G5), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G171), .B2(new_n697), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1961), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n697), .A2(G20), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT23), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n563), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n558), .B1(new_n559), .B2(new_n510), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n786), .B1(new_n789), .B2(new_n697), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1956), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n784), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n759), .A2(new_n776), .A3(new_n781), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n706), .A2(G32), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n478), .A2(G141), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT96), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n487), .A2(G129), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT97), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT26), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n803), .A2(new_n804), .B1(G105), .B2(new_n622), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n797), .A2(new_n800), .A3(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT98), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n806), .A2(new_n807), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n794), .B1(new_n811), .B2(new_n706), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT27), .B(G1996), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  AND3_X1   g389(.A1(G168), .A2(KEYINPUT99), .A3(G16), .ZN(new_n815));
  AOI21_X1  g390(.A(KEYINPUT99), .B1(G168), .B2(G16), .ZN(new_n816));
  OAI22_X1  g391(.A1(new_n815), .A2(new_n816), .B1(G16), .B2(G21), .ZN(new_n817));
  INV_X1    g392(.A(G1966), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n793), .A2(new_n814), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n723), .A2(new_n725), .A3(new_n820), .ZN(G150));
  INV_X1    g396(.A(G150), .ZN(G311));
  NAND2_X1  g397(.A1(new_n778), .A2(G559), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT38), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n534), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(new_n536), .ZN(new_n826));
  INV_X1    g401(.A(G55), .ZN(new_n827));
  INV_X1    g402(.A(G93), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n525), .A2(new_n827), .B1(new_n510), .B2(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n616), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n826), .A2(new_n829), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n549), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n824), .B(new_n834), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n836), .A2(new_n613), .A3(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n832), .A2(new_n613), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT37), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n840), .ZN(G145));
  OAI21_X1  g416(.A(new_n768), .B1(new_n809), .B2(new_n810), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n806), .A2(new_n807), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n843), .A2(new_n808), .A3(new_n767), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n496), .A2(new_n499), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n490), .A2(new_n493), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AND3_X1   g422(.A1(new_n842), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n847), .B1(new_n842), .B2(new_n844), .ZN(new_n849));
  OAI22_X1  g424(.A1(new_n848), .A2(new_n849), .B1(new_n747), .B2(new_n744), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n842), .A2(new_n844), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(G164), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n842), .A2(new_n844), .A3(new_n847), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n852), .A2(new_n748), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n487), .A2(G130), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n476), .A2(G118), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n858), .B1(G142), .B2(new_n478), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(new_n713), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n625), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n850), .A2(new_n854), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT101), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n850), .A2(new_n854), .ZN(new_n864));
  INV_X1    g439(.A(new_n861), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n864), .A2(KEYINPUT101), .A3(new_n865), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n633), .B(new_n480), .ZN(new_n870));
  XOR2_X1   g445(.A(G162), .B(new_n870), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n871), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n862), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(G37), .B1(new_n874), .B2(new_n866), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n872), .A2(KEYINPUT40), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT40), .B1(new_n872), .B2(new_n875), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(G395));
  NAND2_X1  g453(.A1(G305), .A2(G166), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n577), .A2(G303), .A3(new_n581), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n569), .B(new_n570), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n882), .A2(G290), .A3(new_n568), .ZN(new_n883));
  NAND2_X1  g458(.A1(G288), .A2(new_n588), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n881), .A2(new_n885), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(KEYINPUT106), .B2(KEYINPUT42), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n889), .B(KEYINPUT107), .Z(new_n890));
  NAND2_X1  g465(.A1(new_n606), .A2(new_n789), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n778), .A2(G299), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n606), .A2(KEYINPUT103), .A3(new_n789), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n606), .A2(new_n789), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n900), .A2(new_n897), .ZN(new_n901));
  AOI22_X1  g476(.A1(new_n898), .A2(new_n899), .B1(new_n891), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n896), .A2(KEYINPUT104), .A3(new_n897), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n834), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n905), .B1(new_n831), .B2(new_n833), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n619), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n831), .A2(new_n833), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n910), .A2(KEYINPUT102), .ZN(new_n911));
  INV_X1    g486(.A(new_n619), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n911), .A2(new_n912), .A3(new_n907), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n904), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n891), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n918), .A2(new_n900), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT105), .B1(new_n914), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n920), .B1(new_n914), .B2(new_n904), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n890), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n889), .B(KEYINPUT107), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n904), .A2(new_n914), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n923), .B(new_n916), .C1(new_n924), .C2(new_n920), .ZN(new_n925));
  AND2_X1   g500(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n922), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n926), .B1(new_n922), .B2(new_n925), .ZN(new_n928));
  OAI21_X1  g503(.A(G868), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n830), .A2(new_n617), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(G295));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n930), .ZN(G331));
  NAND2_X1  g507(.A1(G171), .A2(G168), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n541), .A2(new_n531), .A3(new_n532), .A4(new_n542), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n910), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n834), .A2(new_n933), .A3(new_n934), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n938), .A2(new_n919), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(new_n940), .A3(new_n937), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n834), .A2(new_n933), .A3(KEYINPUT108), .A4(new_n934), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n939), .B1(new_n904), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT109), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT109), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n943), .B1(new_n902), .B2(new_n903), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n947), .B1(new_n948), .B2(new_n939), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT110), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n888), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n886), .A2(KEYINPUT110), .A3(new_n887), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n946), .A2(new_n949), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(G37), .B1(new_n945), .B2(new_n888), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT43), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n919), .B1(new_n941), .B2(new_n942), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n901), .A2(new_n893), .A3(new_n895), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n897), .B1(new_n918), .B2(new_n900), .ZN(new_n959));
  AOI22_X1  g534(.A1(new_n958), .A2(new_n959), .B1(new_n936), .B2(new_n937), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n953), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT111), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n953), .B(new_n963), .C1(new_n957), .C2(new_n960), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n955), .A2(new_n965), .A3(KEYINPUT43), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT44), .B1(new_n956), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n969), .B1(new_n954), .B2(new_n955), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n955), .A2(new_n965), .A3(new_n969), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n968), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n967), .A2(new_n972), .ZN(G397));
  XNOR2_X1  g548(.A(new_n767), .B(G2067), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n475), .A2(new_n479), .A3(G40), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT112), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n475), .A2(new_n479), .A3(KEYINPUT112), .A4(G40), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(G164), .B2(G1384), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  OR3_X1    g558(.A1(new_n974), .A2(KEYINPUT114), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n811), .A2(G1996), .ZN(new_n985));
  INV_X1    g560(.A(G1996), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n986), .B1(new_n809), .B2(new_n810), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n985), .A2(new_n982), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT114), .B1(new_n974), .B2(new_n983), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n984), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  XOR2_X1   g565(.A(new_n713), .B(new_n715), .Z(new_n991));
  OAI21_X1  g566(.A(new_n990), .B1(new_n983), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n982), .A2(G1986), .A3(G290), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n982), .A2(new_n719), .A3(new_n588), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  XOR2_X1   g570(.A(new_n995), .B(KEYINPUT113), .Z(new_n996));
  NOR2_X1   g571(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT126), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n999));
  INV_X1    g574(.A(G8), .ZN(new_n1000));
  NOR3_X1   g575(.A1(G166), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  INV_X1    g579(.A(G1384), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1004), .B1(new_n847), .B2(new_n1005), .ZN(new_n1006));
  AOI211_X1 g581(.A(KEYINPUT50), .B(G1384), .C1(new_n845), .C2(new_n846), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n979), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(KEYINPUT115), .B(G2090), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n847), .A2(KEYINPUT45), .A3(new_n1005), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n981), .A2(new_n1010), .A3(new_n977), .A4(new_n978), .ZN(new_n1011));
  INV_X1    g586(.A(G1971), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n1008), .A2(new_n1009), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1003), .B1(new_n1013), .B2(new_n1000), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1016));
  AOI21_X1  g591(.A(G1384), .B1(new_n845), .B2(new_n846), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n1004), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1018), .A2(new_n1019), .A3(new_n977), .A4(new_n978), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1009), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1015), .B(G8), .C1(new_n1016), .C2(new_n1022), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n1014), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1976), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT52), .B1(G288), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n977), .A2(new_n1017), .A3(new_n978), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n882), .A2(G1976), .A3(new_n568), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1026), .A2(G8), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(G8), .ZN(new_n1030));
  NOR2_X1   g605(.A1(G288), .A2(new_n1025), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT52), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G1981), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n576), .A2(KEYINPUT76), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT76), .ZN(new_n1036));
  AOI211_X1 g611(.A(new_n1036), .B(new_n536), .C1(new_n574), .C2(new_n575), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1034), .B(new_n581), .C1(new_n1035), .C2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(G1981), .B1(new_n580), .B2(new_n576), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT116), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1041), .B(G1981), .C1(new_n580), .C2(new_n576), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1038), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT49), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT117), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1043), .A2(new_n1047), .A3(new_n1044), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1030), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n524), .A2(new_n534), .A3(G86), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n534), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1050), .B(new_n578), .C1(new_n1051), .C2(new_n536), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1041), .B1(new_n1052), .B2(G1981), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1042), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1055), .A2(KEYINPUT118), .A3(KEYINPUT49), .A4(new_n1038), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1033), .B1(new_n1049), .B2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n1011), .B2(G2078), .ZN(new_n1062));
  INV_X1    g637(.A(G1961), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1020), .A2(new_n1063), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1010), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n977), .B(new_n978), .C1(KEYINPUT45), .C2(new_n1017), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n981), .A2(KEYINPUT119), .A3(new_n977), .A4(new_n978), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n444), .A2(KEYINPUT53), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1065), .A2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1024), .A2(G171), .A3(new_n1060), .A4(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(G1966), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1020), .A2(G2084), .ZN(new_n1076));
  OAI21_X1  g651(.A(G286), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT45), .B1(new_n847), .B2(new_n1005), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1068), .B1(new_n979), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1079), .A2(new_n1070), .A3(new_n1010), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n818), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1076), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(G168), .A3(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1077), .A2(new_n1083), .A3(G8), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT51), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1076), .B1(new_n1080), .B2(new_n818), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1000), .B1(new_n1086), .B2(G168), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT51), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1074), .B1(new_n1090), .B2(KEYINPUT62), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1085), .A2(new_n1092), .A3(new_n1089), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n998), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1088), .B1(new_n1087), .B2(new_n1077), .ZN(new_n1095));
  AOI211_X1 g670(.A(KEYINPUT51), .B(new_n1000), .C1(new_n1086), .C2(G168), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT62), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1074), .ZN(new_n1098));
  AND4_X1   g673(.A1(new_n998), .A2(new_n1097), .A3(new_n1093), .A4(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1094), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1101), .A2(KEYINPUT57), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(KEYINPUT57), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n789), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(G299), .A2(new_n1101), .A3(KEYINPUT57), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  XOR2_X1   g682(.A(KEYINPUT56), .B(G2072), .Z(new_n1108));
  OR2_X1    g683(.A1(new_n1011), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G1956), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1020), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1107), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1027), .A2(G2067), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1113), .B1(new_n780), .B2(new_n1020), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1114), .A2(new_n606), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1107), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1112), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT61), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1116), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1118), .B1(new_n1119), .B2(new_n1112), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n1106), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1122), .A2(KEYINPUT61), .A3(new_n1116), .ZN(new_n1123));
  AOI211_X1 g698(.A(new_n778), .B(new_n1113), .C1(new_n780), .C2(new_n1020), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT60), .B1(new_n1115), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT60), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1114), .A2(new_n1126), .A3(new_n778), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1120), .A2(new_n1123), .A3(new_n1125), .A4(new_n1127), .ZN(new_n1128));
  XOR2_X1   g703(.A(KEYINPUT58), .B(G1341), .Z(new_n1129));
  NAND2_X1  g704(.A1(new_n1027), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT122), .B(G1996), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1132), .B1(new_n1011), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n549), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1136), .B(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1117), .B1(new_n1128), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1073), .A2(G171), .ZN(new_n1140));
  INV_X1    g715(.A(new_n975), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n981), .A2(new_n1010), .A3(new_n1141), .A4(new_n1071), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1065), .A2(G301), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT54), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1030), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1145), .A2(new_n1059), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1033), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1147), .A2(new_n1014), .A3(new_n1023), .A4(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1144), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1065), .A2(G301), .A3(new_n1072), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1062), .A2(new_n1064), .A3(new_n1142), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(G171), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1151), .A2(KEYINPUT54), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1151), .A2(KEYINPUT125), .A3(KEYINPUT54), .A4(new_n1153), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1139), .A2(new_n1090), .A3(new_n1150), .A4(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT63), .ZN(new_n1160));
  OAI211_X1 g735(.A(G8), .B(G168), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1160), .B1(new_n1149), .B2(new_n1161), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1086), .A2(new_n1000), .A3(G286), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1024), .A2(KEYINPUT63), .A3(new_n1060), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(G288), .A2(G1976), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1147), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n1038), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1023), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1168), .A2(new_n1146), .B1(new_n1060), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT120), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1165), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1171), .B1(new_n1165), .B2(new_n1170), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1159), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n997), .B1(new_n1100), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n983), .B1(new_n974), .B2(new_n811), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT46), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n982), .A2(new_n986), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1176), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1179), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1180));
  XOR2_X1   g755(.A(new_n1180), .B(KEYINPUT47), .Z(new_n1181));
  NOR2_X1   g756(.A1(new_n713), .A2(new_n715), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n990), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n767), .A2(new_n770), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n983), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  XOR2_X1   g760(.A(new_n994), .B(KEYINPUT48), .Z(new_n1186));
  NOR2_X1   g761(.A1(new_n992), .A2(new_n1186), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1181), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1175), .A2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g764(.A1(new_n970), .A2(new_n971), .ZN(new_n1191));
  NOR2_X1   g765(.A1(G227), .A2(new_n462), .ZN(new_n1192));
  XNOR2_X1  g766(.A(new_n1192), .B(KEYINPUT127), .ZN(new_n1193));
  NOR3_X1   g767(.A1(G401), .A2(new_n1193), .A3(G229), .ZN(new_n1194));
  INV_X1    g768(.A(new_n875), .ZN(new_n1195));
  AOI21_X1  g769(.A(new_n873), .B1(new_n867), .B2(new_n868), .ZN(new_n1196));
  OAI21_X1  g770(.A(new_n1194), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g771(.A1(new_n1191), .A2(new_n1197), .ZN(G308));
  OAI221_X1 g772(.A(new_n1194), .B1(new_n1195), .B2(new_n1196), .C1(new_n970), .C2(new_n971), .ZN(G225));
endmodule


