//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n204));
  INV_X1    g003(.A(G29gat), .ZN(new_n205));
  INV_X1    g004(.A(G36gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NOR3_X1   g006(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT94), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI211_X1 g011(.A(KEYINPUT94), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI211_X1 g013(.A(new_n203), .B(new_n207), .C1(new_n209), .C2(new_n214), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n214), .A2(KEYINPUT95), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n214), .A2(KEYINPUT95), .B1(G29gat), .B2(G36gat), .ZN(new_n217));
  AOI211_X1 g016(.A(new_n208), .B(new_n204), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(KEYINPUT17), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT96), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT97), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n225), .A2(G1gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(G1gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT16), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G8gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT98), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n230), .B(G8gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT98), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n219), .A2(KEYINPUT17), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n234), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n235), .B1(new_n215), .B2(new_n218), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G229gat), .A2(G233gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(KEYINPUT18), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n232), .A2(new_n219), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  XOR2_X1   g044(.A(new_n242), .B(KEYINPUT13), .Z(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n239), .A2(new_n242), .A3(new_n240), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT18), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n243), .A2(new_n247), .A3(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G113gat), .B(G141gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(G197gat), .ZN(new_n253));
  XOR2_X1   g052(.A(KEYINPUT11), .B(G169gat), .Z(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT93), .B(KEYINPUT12), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n255), .B(new_n256), .Z(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n251), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n243), .A2(new_n257), .A3(new_n247), .A4(new_n250), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G190gat), .B(G218gat), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n220), .B(KEYINPUT96), .ZN(new_n264));
  NAND2_X1  g063(.A1(G85gat), .A2(G92gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT7), .ZN(new_n266));
  NAND2_X1  g065(.A1(G99gat), .A2(G106gat), .ZN(new_n267));
  INV_X1    g066(.A(G85gat), .ZN(new_n268));
  INV_X1    g067(.A(G92gat), .ZN(new_n269));
  AOI22_X1  g068(.A1(KEYINPUT8), .A2(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(G99gat), .B(G106gat), .Z(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n237), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n264), .A2(new_n274), .ZN(new_n275));
  AND2_X1   g074(.A1(G232gat), .A2(G233gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT41), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n277), .B1(new_n219), .B2(new_n273), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n263), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n278), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n280), .B(new_n262), .C1(new_n264), .C2(new_n274), .ZN(new_n281));
  XOR2_X1   g080(.A(G134gat), .B(G162gat), .Z(new_n282));
  NOR2_X1   g081(.A1(new_n276), .A2(KEYINPUT41), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT100), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n279), .A2(new_n281), .A3(KEYINPUT101), .A4(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n279), .A2(new_n281), .A3(new_n285), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT101), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n284), .B1(new_n279), .B2(new_n281), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n286), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT21), .ZN(new_n292));
  XNOR2_X1  g091(.A(G57gat), .B(G64gat), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G71gat), .B(G78gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n232), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n292), .ZN(new_n299));
  XNOR2_X1  g098(.A(G127gat), .B(G155gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n298), .B(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G231gat), .A2(G233gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT99), .ZN(new_n304));
  XOR2_X1   g103(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G183gat), .B(G211gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n302), .A2(new_n308), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G230gat), .ZN(new_n312));
  INV_X1    g111(.A(G233gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(new_n273), .B(new_n297), .Z(new_n315));
  INV_X1    g114(.A(KEYINPUT10), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OR3_X1    g116(.A1(new_n273), .A2(new_n316), .A3(new_n297), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n314), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NOR3_X1   g118(.A1(new_n315), .A2(new_n312), .A3(new_n313), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(G120gat), .B(G148gat), .Z(new_n322));
  XNOR2_X1  g121(.A(new_n322), .B(KEYINPUT102), .ZN(new_n323));
  XNOR2_X1  g122(.A(G176gat), .B(G204gat), .ZN(new_n324));
  XOR2_X1   g123(.A(new_n323), .B(new_n324), .Z(new_n325));
  OR2_X1    g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n321), .A2(new_n325), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n291), .A2(new_n311), .A3(new_n329), .ZN(new_n330));
  XOR2_X1   g129(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n331));
  INV_X1    g130(.A(KEYINPUT27), .ZN(new_n332));
  INV_X1    g131(.A(G183gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n332), .B1(new_n333), .B2(KEYINPUT67), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT67), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n335), .A2(KEYINPUT66), .A3(KEYINPUT27), .A4(G183gat), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n334), .B(new_n336), .C1(KEYINPUT66), .C2(G183gat), .ZN(new_n337));
  INV_X1    g136(.A(G190gat), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n331), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT27), .B(G183gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n340), .A2(KEYINPUT28), .A3(new_n338), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(KEYINPUT69), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT69), .ZN(new_n344));
  NOR2_X1   g143(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n335), .A2(G183gat), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n345), .B1(new_n346), .B2(new_n332), .ZN(new_n347));
  AOI21_X1  g146(.A(G190gat), .B1(new_n347), .B2(new_n336), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n344), .B(new_n341), .C1(new_n348), .C2(new_n331), .ZN(new_n349));
  NAND2_X1  g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G169gat), .ZN(new_n352));
  INV_X1    g151(.A(G176gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n351), .B1(KEYINPUT26), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n355), .B1(KEYINPUT26), .B2(new_n354), .ZN(new_n356));
  NAND2_X1  g155(.A1(G183gat), .A2(G190gat), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n343), .A2(new_n349), .A3(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(KEYINPUT64), .B(G176gat), .Z(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(KEYINPUT23), .A3(new_n352), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n357), .A2(KEYINPUT24), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT24), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(G183gat), .A3(G190gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n365), .B1(G183gat), .B2(G190gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT23), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n351), .B1(new_n367), .B2(new_n354), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n361), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT25), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n350), .B1(new_n354), .B2(new_n367), .ZN(new_n372));
  OR2_X1    g171(.A1(new_n372), .A2(KEYINPUT65), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT66), .B(G183gat), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n365), .B1(new_n374), .B2(G190gat), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n370), .B1(new_n354), .B2(new_n367), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n372), .A2(KEYINPUT65), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n373), .A2(new_n375), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n371), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n359), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT29), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(G226gat), .A2(G233gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(KEYINPUT78), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n356), .A2(new_n357), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n341), .B1(new_n348), .B2(new_n331), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n387), .B1(new_n388), .B2(KEYINPUT69), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n389), .A2(new_n349), .B1(new_n371), .B2(new_n378), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT79), .B1(new_n390), .B2(new_n385), .ZN(new_n391));
  XOR2_X1   g190(.A(G197gat), .B(G204gat), .Z(new_n392));
  XNOR2_X1  g191(.A(KEYINPUT76), .B(G211gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT77), .B(G218gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT22), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n392), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G211gat), .B(G218gat), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n397), .A2(new_n398), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n385), .B1(new_n359), .B2(new_n379), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT79), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n386), .A2(new_n391), .A3(new_n402), .A4(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n384), .B1(new_n380), .B2(new_n381), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n401), .B1(new_n407), .B2(new_n403), .ZN(new_n408));
  XNOR2_X1  g207(.A(G8gat), .B(G36gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(G64gat), .B(G92gat), .ZN(new_n410));
  XOR2_X1   g209(.A(new_n409), .B(new_n410), .Z(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT30), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n406), .A2(new_n408), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n404), .B1(new_n380), .B2(new_n384), .ZN(new_n416));
  AOI211_X1 g215(.A(KEYINPUT79), .B(new_n385), .C1(new_n359), .C2(new_n379), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT29), .B1(new_n359), .B2(new_n379), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n402), .B1(new_n419), .B2(new_n384), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n380), .A2(new_n384), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n422), .B1(new_n384), .B2(new_n419), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n418), .A2(new_n421), .B1(new_n423), .B2(new_n401), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n415), .B1(new_n424), .B2(new_n411), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT30), .B1(new_n424), .B2(new_n411), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n428));
  INV_X1    g227(.A(G113gat), .ZN(new_n429));
  INV_X1    g228(.A(G120gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G113gat), .A2(G120gat), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(KEYINPUT72), .A3(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT1), .ZN(new_n434));
  INV_X1    g233(.A(G134gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(G127gat), .ZN(new_n436));
  INV_X1    g235(.A(G127gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(G134gat), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n433), .A2(new_n434), .A3(new_n436), .A4(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT72), .B1(new_n431), .B2(new_n432), .ZN(new_n440));
  OR2_X1    g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT71), .ZN(new_n442));
  INV_X1    g241(.A(new_n432), .ZN(new_n443));
  NOR2_X1   g242(.A1(G113gat), .A2(G120gat), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n443), .A2(new_n444), .A3(KEYINPUT1), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT70), .B1(new_n436), .B2(new_n438), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n436), .A2(new_n438), .A3(KEYINPUT70), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n442), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT70), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n437), .A2(G134gat), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n435), .A2(G127gat), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n431), .A2(new_n434), .A3(new_n432), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n453), .A2(new_n442), .A3(new_n448), .A4(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n441), .B1(new_n449), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(G155gat), .A2(G162gat), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(G155gat), .A2(G162gat), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n458), .A2(KEYINPUT2), .ZN(new_n462));
  XNOR2_X1  g261(.A(G141gat), .B(G148gat), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n462), .B1(new_n463), .B2(KEYINPUT80), .ZN(new_n464));
  INV_X1    g263(.A(G148gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(G141gat), .ZN(new_n466));
  INV_X1    g265(.A(G141gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(G148gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT80), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n461), .B1(new_n464), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(KEYINPUT81), .B(G141gat), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n466), .B1(new_n473), .B2(new_n465), .ZN(new_n474));
  INV_X1    g273(.A(G155gat), .ZN(new_n475));
  INV_X1    g274(.A(G162gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n477), .A2(KEYINPUT82), .A3(new_n458), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT82), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n479), .B1(new_n459), .B2(new_n460), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n474), .A2(new_n462), .A3(new_n478), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n472), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n457), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n439), .A2(new_n440), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n453), .A2(new_n448), .A3(new_n454), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT71), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n484), .B1(new_n486), .B2(new_n455), .ZN(new_n487));
  INV_X1    g286(.A(new_n461), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n469), .A2(new_n470), .B1(KEYINPUT2), .B2(new_n458), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n463), .A2(KEYINPUT80), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n480), .A2(new_n478), .A3(new_n462), .ZN(new_n492));
  INV_X1    g291(.A(new_n466), .ZN(new_n493));
  AND2_X1   g292(.A1(KEYINPUT81), .A2(G141gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(KEYINPUT81), .A2(G141gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n493), .B1(new_n496), .B2(G148gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n491), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n487), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G225gat), .A2(G233gat), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n428), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT4), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(new_n457), .B2(new_n482), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT3), .B1(new_n491), .B2(new_n498), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT3), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n472), .A2(new_n481), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n457), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n487), .A2(new_n499), .A3(KEYINPUT4), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n506), .A2(new_n510), .A3(new_n511), .A4(new_n502), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n504), .A2(new_n512), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n457), .A2(new_n505), .A3(new_n482), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT4), .B1(new_n487), .B2(new_n499), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n428), .A2(new_n502), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n491), .A2(new_n498), .A3(KEYINPUT3), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n518), .A2(new_n487), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n517), .B1(new_n519), .B2(new_n507), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT84), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n517), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n506), .A2(new_n510), .A3(new_n511), .A4(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT84), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n513), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G1gat), .B(G29gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(KEYINPUT0), .ZN(new_n528));
  XNOR2_X1  g327(.A(G57gat), .B(G85gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n516), .A2(new_n520), .A3(KEYINPUT84), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n523), .A2(new_n524), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n530), .B1(new_n504), .B2(new_n512), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT6), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n531), .A2(KEYINPUT90), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n530), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n538), .B1(new_n534), .B2(new_n513), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT6), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT90), .B1(new_n531), .B2(new_n536), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n427), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT92), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G228gat), .A2(G233gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n509), .A2(new_n381), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n401), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n381), .B1(new_n399), .B2(new_n400), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n499), .B1(new_n550), .B2(new_n508), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n546), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT87), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n546), .B1(new_n548), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n401), .A2(new_n547), .A3(KEYINPUT87), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n550), .A2(KEYINPUT86), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT3), .B1(new_n550), .B2(KEYINPUT86), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n499), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n552), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(KEYINPUT31), .B(G50gat), .Z(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G78gat), .B(G106gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(G22gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n561), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n565), .B(new_n552), .C1(new_n556), .C2(new_n559), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n562), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n564), .B1(new_n562), .B2(new_n566), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G227gat), .A2(G233gat), .ZN(new_n570));
  AND3_X1   g369(.A1(new_n359), .A2(new_n457), .A3(new_n379), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n457), .B1(new_n359), .B2(new_n379), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n570), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT34), .B1(new_n574), .B2(KEYINPUT75), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n573), .B(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n380), .A2(new_n487), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n359), .A2(new_n457), .A3(new_n379), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n578), .A2(new_n574), .A3(new_n579), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n580), .A2(KEYINPUT32), .ZN(new_n581));
  XNOR2_X1  g380(.A(G15gat), .B(G43gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(G71gat), .B(G99gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT33), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n584), .B1(new_n580), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n581), .B1(KEYINPUT73), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT33), .B1(new_n584), .B2(KEYINPUT74), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n588), .B1(KEYINPUT74), .B2(new_n584), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n580), .A2(KEYINPUT32), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT73), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n590), .B1(new_n586), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n577), .B1(new_n587), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n584), .ZN(new_n594));
  NOR3_X1   g393(.A1(new_n571), .A2(new_n572), .A3(new_n570), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n591), .B(new_n594), .C1(new_n595), .C2(KEYINPUT33), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(new_n581), .A3(new_n589), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n580), .A2(KEYINPUT32), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n594), .B1(new_n595), .B2(KEYINPUT33), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n598), .B1(new_n599), .B2(new_n591), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n573), .B(new_n575), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n597), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n593), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT35), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n569), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  OAI211_X1 g404(.A(KEYINPUT92), .B(new_n427), .C1(new_n541), .C2(new_n542), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n545), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n534), .A2(new_n535), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT6), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT85), .B1(new_n610), .B2(new_n539), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT85), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n531), .A2(new_n612), .A3(new_n536), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(new_n613), .A3(new_n540), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n427), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n569), .A2(new_n603), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT35), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n607), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT89), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT40), .ZN(new_n620));
  OAI21_X1  g419(.A(KEYINPUT39), .B1(new_n501), .B2(new_n503), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT88), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI211_X1 g422(.A(KEYINPUT88), .B(KEYINPUT39), .C1(new_n501), .C2(new_n503), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n506), .A2(new_n511), .A3(new_n510), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n503), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n538), .B1(new_n626), .B2(KEYINPUT39), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n620), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n626), .A2(KEYINPUT39), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n630), .A2(new_n631), .A3(KEYINPUT40), .A4(new_n538), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n629), .A2(new_n531), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n619), .B1(new_n633), .B2(new_n427), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n632), .A2(new_n531), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n391), .A2(new_n405), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n408), .B1(new_n636), .B2(new_n420), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n413), .B1(new_n637), .B2(new_n412), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n411), .B1(new_n406), .B2(new_n408), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(new_n640), .A3(new_n415), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n635), .A2(new_n641), .A3(KEYINPUT89), .A4(new_n629), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n634), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n537), .A2(new_n540), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT91), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT37), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n411), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n637), .B2(new_n412), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT38), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n403), .B1(new_n382), .B2(new_n385), .ZN(new_n650));
  OAI21_X1  g449(.A(KEYINPUT37), .B1(new_n650), .B2(new_n401), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n401), .B1(new_n419), .B2(new_n384), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n649), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n645), .B1(new_n648), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n646), .B1(new_n423), .B2(new_n402), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n386), .A2(new_n391), .A3(new_n401), .A4(new_n405), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT38), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n658), .B(KEYINPUT91), .C1(new_n639), .C2(new_n647), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  OAI22_X1  g459(.A1(new_n639), .A2(new_n647), .B1(new_n424), .B2(new_n646), .ZN(new_n661));
  AOI22_X1  g460(.A1(new_n661), .A2(KEYINPUT38), .B1(new_n424), .B2(new_n411), .ZN(new_n662));
  INV_X1    g461(.A(new_n542), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n644), .A2(new_n660), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n643), .A2(new_n664), .A3(new_n569), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n569), .B1(new_n614), .B2(new_n427), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT36), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n587), .A2(new_n592), .A3(new_n577), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n601), .B1(new_n597), .B2(new_n600), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n593), .A2(new_n602), .A3(KEYINPUT36), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n665), .A2(new_n673), .ZN(new_n674));
  AOI211_X1 g473(.A(new_n261), .B(new_n330), .C1(new_n618), .C2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n614), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT104), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT103), .B(G1gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1324gat));
  XOR2_X1   g479(.A(KEYINPUT16), .B(G8gat), .Z(new_n681));
  AND3_X1   g480(.A1(new_n675), .A2(new_n641), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n231), .B1(new_n675), .B2(new_n641), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT42), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(KEYINPUT42), .B2(new_n682), .ZN(G1325gat));
  AOI21_X1  g484(.A(G15gat), .B1(new_n675), .B2(new_n603), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n672), .A2(G15gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT105), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n686), .B1(new_n675), .B2(new_n688), .ZN(G1326gat));
  INV_X1    g488(.A(new_n569), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT43), .B(G22gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  AOI21_X1  g492(.A(new_n291), .B1(new_n618), .B2(new_n674), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n261), .A2(new_n311), .A3(new_n328), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n697), .A2(new_n205), .A3(new_n676), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT106), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT45), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n618), .A2(new_n674), .ZN(new_n704));
  INV_X1    g503(.A(new_n291), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n291), .A2(new_n707), .ZN(new_n708));
  OAI211_X1 g507(.A(KEYINPUT107), .B(new_n286), .C1(new_n289), .C2(new_n290), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(new_n703), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n710), .B1(new_n674), .B2(new_n618), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n695), .B1(new_n706), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  OAI211_X1 g514(.A(KEYINPUT108), .B(new_n695), .C1(new_n706), .C2(new_n711), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n715), .A2(new_n614), .A3(new_n717), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n701), .B(new_n702), .C1(new_n718), .C2(new_n205), .ZN(G1328gat));
  NOR3_X1   g518(.A1(new_n696), .A2(G36gat), .A3(new_n427), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT46), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n715), .A2(new_n427), .A3(new_n717), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n722), .B2(new_n206), .ZN(G1329gat));
  AOI21_X1  g522(.A(G43gat), .B1(new_n593), .B2(new_n602), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n697), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT47), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n706), .A2(new_n711), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(new_n672), .A3(new_n695), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n726), .B1(new_n728), .B2(G43gat), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n729), .A2(KEYINPUT110), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(KEYINPUT110), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n672), .A3(new_n716), .ZN(new_n732));
  AOI22_X1  g531(.A1(new_n732), .A2(G43gat), .B1(new_n697), .B2(new_n724), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n734));
  OAI211_X1 g533(.A(new_n730), .B(new_n731), .C1(new_n733), .C2(new_n734), .ZN(G1330gat));
  OAI21_X1  g534(.A(G50gat), .B1(new_n712), .B2(new_n569), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n696), .A2(G50gat), .A3(new_n569), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT48), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n714), .A2(new_n690), .A3(new_n716), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n741), .A2(KEYINPUT111), .A3(G50gat), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT111), .B1(new_n741), .B2(G50gat), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n742), .A2(new_n743), .A3(new_n737), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n740), .B1(new_n744), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g544(.A1(new_n259), .A2(new_n260), .ZN(new_n746));
  INV_X1    g545(.A(new_n311), .ZN(new_n747));
  NOR4_X1   g546(.A1(new_n705), .A2(new_n746), .A3(new_n747), .A4(new_n329), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n704), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n749), .A2(new_n614), .ZN(new_n750));
  XNOR2_X1  g549(.A(KEYINPUT112), .B(G57gat), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1332gat));
  NOR2_X1   g551(.A1(new_n749), .A2(new_n427), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT49), .B(G64gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT113), .ZN(G1333gat));
  INV_X1    g557(.A(new_n672), .ZN(new_n759));
  OAI21_X1  g558(.A(G71gat), .B1(new_n749), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(G71gat), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n603), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(new_n749), .B2(new_n762), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g563(.A1(new_n749), .A2(new_n569), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(G78gat), .Z(G1335gat));
  NAND2_X1  g565(.A1(new_n261), .A2(new_n747), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT114), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n727), .A2(new_n328), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G85gat), .B1(new_n770), .B2(new_n614), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n694), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n772), .A2(KEYINPUT115), .A3(new_n773), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n774), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n676), .A2(new_n268), .A3(new_n328), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n771), .B1(new_n780), .B2(new_n781), .ZN(G1336gat));
  AOI21_X1  g581(.A(new_n269), .B1(new_n769), .B2(new_n641), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n783), .A2(KEYINPUT52), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n329), .A2(G92gat), .A3(new_n427), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n779), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n774), .A2(KEYINPUT116), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n774), .A2(KEYINPUT116), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n788), .B(new_n789), .C1(new_n777), .C2(new_n778), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n783), .B1(new_n790), .B2(new_n785), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n787), .B1(new_n791), .B2(new_n792), .ZN(G1337gat));
  XOR2_X1   g592(.A(KEYINPUT118), .B(G99gat), .Z(new_n794));
  AND2_X1   g593(.A1(new_n328), .A2(new_n603), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n779), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT117), .B1(new_n770), .B2(new_n759), .ZN(new_n797));
  INV_X1    g596(.A(new_n794), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n770), .A2(KEYINPUT117), .A3(new_n759), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n796), .B1(new_n799), .B2(new_n800), .ZN(G1338gat));
  NAND2_X1  g600(.A1(new_n769), .A2(new_n690), .ZN(new_n802));
  XNOR2_X1  g601(.A(KEYINPUT119), .B(G106gat), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT53), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n329), .A2(G106gat), .A3(new_n569), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n780), .B2(new_n806), .ZN(new_n807));
  AOI22_X1  g606(.A1(new_n790), .A2(new_n805), .B1(new_n802), .B2(new_n803), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(G1339gat));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n319), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n317), .A2(new_n318), .A3(new_n314), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n325), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n319), .B2(new_n811), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n814), .A2(KEYINPUT55), .A3(new_n816), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(new_n326), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n746), .A2(new_n822), .ZN(new_n823));
  OAI22_X1  g622(.A1(new_n241), .A2(new_n242), .B1(new_n245), .B2(new_n246), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n255), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n260), .A2(new_n825), .A3(new_n328), .ZN(new_n826));
  AOI22_X1  g625(.A1(new_n823), .A2(new_n826), .B1(new_n708), .B2(new_n709), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n260), .A2(new_n825), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(new_n821), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n829), .A2(new_n708), .A3(new_n709), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n747), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n330), .A2(new_n746), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n569), .A3(new_n603), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n614), .A2(new_n641), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT120), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(new_n429), .A3(new_n746), .ZN(new_n840));
  INV_X1    g639(.A(new_n838), .ZN(new_n841));
  OAI21_X1  g640(.A(G113gat), .B1(new_n841), .B2(new_n261), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(G1340gat));
  NAND3_X1  g642(.A1(new_n839), .A2(new_n430), .A3(new_n328), .ZN(new_n844));
  OAI21_X1  g643(.A(G120gat), .B1(new_n841), .B2(new_n329), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(G1341gat));
  NAND2_X1  g645(.A1(new_n838), .A2(new_n311), .ZN(new_n847));
  XOR2_X1   g646(.A(KEYINPUT121), .B(G127gat), .Z(new_n848));
  XNOR2_X1  g647(.A(new_n847), .B(new_n848), .ZN(G1342gat));
  INV_X1    g648(.A(new_n835), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n291), .A2(new_n641), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n676), .A3(new_n851), .ZN(new_n852));
  OR3_X1    g651(.A1(new_n852), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT56), .B1(new_n852), .B2(G134gat), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(KEYINPUT122), .A3(G134gat), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT122), .B1(new_n852), .B2(G134gat), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n853), .B(new_n854), .C1(new_n856), .C2(new_n857), .ZN(G1343gat));
  INV_X1    g657(.A(KEYINPUT124), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT58), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n837), .A2(new_n672), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n834), .A2(new_n690), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n261), .A2(G141gat), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n860), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT57), .B1(new_n834), .B2(new_n690), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n690), .A2(KEYINPUT57), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT123), .ZN(new_n869));
  AOI22_X1  g668(.A1(new_n746), .A2(new_n822), .B1(new_n826), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n826), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT123), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n705), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n747), .B1(new_n873), .B2(new_n830), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n868), .B1(new_n874), .B2(new_n833), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n746), .B(new_n861), .C1(new_n866), .C2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n865), .B1(new_n876), .B2(new_n473), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n859), .A2(KEYINPUT58), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n877), .B(new_n878), .ZN(G1344gat));
  INV_X1    g678(.A(new_n862), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n465), .A3(new_n328), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(G148gat), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n866), .A2(new_n875), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n884), .A2(new_n672), .A3(new_n837), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n883), .B1(new_n885), .B2(new_n328), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n291), .A2(new_n828), .A3(new_n821), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n747), .B1(new_n873), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n833), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT57), .B1(new_n889), .B2(new_n690), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n829), .A2(new_n708), .A3(new_n709), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n871), .B1(new_n746), .B2(new_n822), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n708), .A2(new_n709), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n832), .B1(new_n894), .B2(new_n747), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n868), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n328), .B(new_n861), .C1(new_n890), .C2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n882), .B1(new_n897), .B2(G148gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n881), .B1(new_n886), .B2(new_n898), .ZN(G1345gat));
  NAND3_X1  g698(.A1(new_n880), .A2(new_n475), .A3(new_n311), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n885), .A2(new_n311), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(new_n475), .ZN(G1346gat));
  AND2_X1   g701(.A1(new_n885), .A2(new_n893), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n834), .A2(new_n690), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n851), .A2(new_n476), .A3(new_n676), .A4(new_n759), .ZN(new_n905));
  OAI22_X1  g704(.A1(new_n903), .A2(new_n476), .B1(new_n904), .B2(new_n905), .ZN(G1347gat));
  NAND2_X1  g705(.A1(new_n614), .A2(new_n641), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT126), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n835), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n911), .A2(new_n352), .A3(new_n261), .ZN(new_n912));
  OAI21_X1  g711(.A(KEYINPUT125), .B1(new_n895), .B2(new_n676), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n834), .A2(new_n914), .A3(new_n614), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n616), .A2(new_n427), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n916), .A2(new_n746), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n912), .B1(new_n352), .B2(new_n918), .ZN(G1348gat));
  NAND2_X1  g718(.A1(new_n916), .A2(new_n917), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n353), .B1(new_n920), .B2(new_n329), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n895), .A2(new_n690), .ZN(new_n922));
  INV_X1    g721(.A(new_n360), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n922), .A2(new_n923), .A3(new_n795), .A4(new_n908), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n921), .A2(new_n924), .ZN(G1349gat));
  INV_X1    g724(.A(new_n374), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n926), .B1(new_n910), .B2(new_n311), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n311), .A2(new_n340), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n928), .B(new_n929), .C1(new_n920), .C2(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n920), .A2(new_n930), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT60), .B1(new_n932), .B2(new_n927), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1350gat));
  INV_X1    g733(.A(KEYINPUT61), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n910), .A2(new_n705), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n936), .B2(G190gat), .ZN(new_n937));
  AOI211_X1 g736(.A(KEYINPUT61), .B(new_n338), .C1(new_n910), .C2(new_n705), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n893), .A2(new_n338), .ZN(new_n939));
  OAI22_X1  g738(.A1(new_n937), .A2(new_n938), .B1(new_n920), .B2(new_n939), .ZN(G1351gat));
  NAND3_X1  g739(.A1(new_n759), .A2(new_n690), .A3(new_n641), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n941), .B1(new_n913), .B2(new_n915), .ZN(new_n942));
  AOI21_X1  g741(.A(G197gat), .B1(new_n942), .B2(new_n746), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n944), .B1(new_n890), .B2(new_n896), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n569), .B1(new_n888), .B2(new_n833), .ZN(new_n946));
  OAI221_X1 g745(.A(KEYINPUT127), .B1(new_n895), .B2(new_n868), .C1(new_n946), .C2(KEYINPUT57), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n909), .A2(new_n672), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n949), .A2(G197gat), .A3(new_n746), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n943), .B1(new_n948), .B2(new_n950), .ZN(G1352gat));
  NOR2_X1   g750(.A1(new_n329), .A2(G204gat), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n942), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n955));
  INV_X1    g754(.A(new_n949), .ZN(new_n956));
  AOI211_X1 g755(.A(new_n329), .B(new_n956), .C1(new_n945), .C2(new_n947), .ZN(new_n957));
  INV_X1    g756(.A(G204gat), .ZN(new_n958));
  OAI211_X1 g757(.A(new_n954), .B(new_n955), .C1(new_n957), .C2(new_n958), .ZN(G1353gat));
  INV_X1    g758(.A(new_n393), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n942), .A2(new_n960), .A3(new_n311), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n311), .B(new_n949), .C1(new_n890), .C2(new_n896), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n962), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT63), .B1(new_n962), .B2(G211gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1354gat));
  AOI21_X1  g764(.A(G218gat), .B1(new_n942), .B2(new_n893), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n956), .B1(new_n945), .B2(new_n947), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n705), .A2(new_n394), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n966), .B1(new_n967), .B2(new_n969), .ZN(G1355gat));
endmodule


