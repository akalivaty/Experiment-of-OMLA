//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G77), .ZN(new_n211));
  INV_X1    g0011(.A(G244), .ZN(new_n212));
  INV_X1    g0012(.A(G107), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n209), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  OR2_X1    g0019(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n209), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT0), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n220), .A2(new_n221), .A3(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G50), .ZN(new_n226));
  INV_X1    g0026(.A(new_n206), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n226), .B1(new_n227), .B2(KEYINPUT67), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n228), .B1(KEYINPUT67), .B2(new_n227), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT68), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(KEYINPUT65), .ZN(new_n232));
  INV_X1    g0032(.A(KEYINPUT65), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n233), .A2(G1), .A3(G13), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AND2_X1   g0036(.A1(KEYINPUT66), .A2(G20), .ZN(new_n237));
  NOR2_X1   g0037(.A1(KEYINPUT66), .A2(G20), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g0039(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g0040(.A(new_n225), .B1(new_n230), .B2(new_n240), .ZN(G361));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  INV_X1    g0042(.A(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT2), .B(G226), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G250), .B(G257), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G264), .B(G270), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G358));
  XNOR2_X1  g0050(.A(G50), .B(G68), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G58), .B(G77), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n251), .B(new_n252), .Z(new_n253));
  XOR2_X1   g0053(.A(G87), .B(G97), .Z(new_n254));
  XNOR2_X1  g0054(.A(G107), .B(G116), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n253), .B(new_n256), .ZN(G351));
  INV_X1    g0057(.A(KEYINPUT70), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT10), .ZN(new_n259));
  OR2_X1    g0059(.A1(new_n258), .A2(KEYINPUT10), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n232), .B(new_n234), .C1(new_n261), .C2(new_n209), .ZN(new_n262));
  INV_X1    g0062(.A(G20), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n263), .B1(new_n227), .B2(new_n226), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n239), .A2(G33), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT8), .B(G58), .ZN(new_n266));
  INV_X1    g0066(.A(G150), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  OAI22_X1  g0069(.A1(new_n265), .A2(new_n266), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n262), .B1(new_n264), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G13), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G1), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G20), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n226), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n262), .A2(new_n275), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G1), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G20), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G50), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n271), .B(new_n276), .C1(new_n278), .C2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT9), .ZN(new_n283));
  XNOR2_X1  g0083(.A(new_n282), .B(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G1), .A3(G13), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G274), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n279), .B1(G41), .B2(G45), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(new_n288), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n291), .A2(G226), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT3), .B(G33), .ZN(new_n293));
  INV_X1    g0093(.A(G1698), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(G222), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(G1698), .ZN(new_n296));
  INV_X1    g0096(.A(G223), .ZN(new_n297));
  OAI221_X1 g0097(.A(new_n295), .B1(new_n211), .B2(new_n293), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n235), .A2(new_n285), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  AOI211_X1 g0100(.A(new_n289), .B(new_n292), .C1(new_n298), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G190), .ZN(new_n302));
  INV_X1    g0102(.A(G200), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n302), .B1(new_n303), .B2(new_n301), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n259), .B(new_n260), .C1(new_n284), .C2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n304), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n282), .B(KEYINPUT9), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n306), .A2(new_n307), .A3(new_n258), .A4(KEYINPUT10), .ZN(new_n308));
  INV_X1    g0108(.A(G179), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n301), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n310), .B(new_n282), .C1(G169), .C2(new_n301), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n305), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n275), .A2(new_n202), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT12), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n277), .A2(G68), .A3(new_n280), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n268), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n265), .B2(new_n211), .ZN(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT11), .B1(new_n318), .B2(new_n262), .ZN(new_n319));
  AND3_X1   g0119(.A1(new_n318), .A2(KEYINPUT11), .A3(new_n262), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n316), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT14), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT71), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n286), .A2(new_n324), .A3(new_n288), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n325), .A2(G238), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n290), .A2(KEYINPUT71), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n289), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT13), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT3), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G33), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n330), .A2(new_n332), .A3(G232), .A4(G1698), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n330), .A2(new_n332), .A3(G226), .A4(new_n294), .ZN(new_n334));
  INV_X1    g0134(.A(G97), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n333), .B(new_n334), .C1(new_n261), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n300), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n328), .A2(new_n329), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n329), .B1(new_n328), .B2(new_n337), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n323), .B(G169), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n326), .A2(new_n327), .ZN(new_n341));
  INV_X1    g0141(.A(new_n287), .ZN(new_n342));
  INV_X1    g0142(.A(new_n288), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n341), .A2(new_n337), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT13), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n328), .A2(new_n329), .A3(new_n337), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(G179), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n340), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n346), .A2(new_n347), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n323), .B1(new_n350), .B2(G169), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n322), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(G200), .ZN(new_n353));
  INV_X1    g0153(.A(G190), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n353), .B(new_n321), .C1(new_n354), .C2(new_n350), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  OR2_X1    g0156(.A1(KEYINPUT66), .A2(G20), .ZN(new_n357));
  NAND2_X1  g0157(.A1(KEYINPUT66), .A2(G20), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G77), .ZN(new_n360));
  XNOR2_X1  g0160(.A(KEYINPUT15), .B(G87), .ZN(new_n361));
  OAI221_X1 g0161(.A(new_n360), .B1(new_n269), .B2(new_n266), .C1(new_n265), .C2(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n362), .A2(new_n262), .B1(new_n211), .B2(new_n275), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n277), .A2(G77), .A3(new_n280), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT69), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n365), .B(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G238), .ZN(new_n368));
  OAI22_X1  g0168(.A1(new_n296), .A2(new_n368), .B1(new_n213), .B2(new_n293), .ZN(new_n369));
  INV_X1    g0169(.A(new_n293), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n370), .A2(new_n243), .A3(G1698), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n300), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n372), .B(new_n344), .C1(new_n212), .C2(new_n290), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G200), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n354), .B2(new_n373), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n367), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n373), .A2(G179), .ZN(new_n377));
  INV_X1    g0177(.A(G169), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n377), .B1(new_n378), .B2(new_n373), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n367), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NOR4_X1   g0181(.A1(new_n312), .A2(new_n356), .A3(new_n376), .A4(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT16), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n331), .A2(KEYINPUT72), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT72), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT3), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n384), .A2(new_n386), .A3(new_n261), .ZN(new_n387));
  NAND2_X1  g0187(.A1(KEYINPUT3), .A2(G33), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n357), .A2(KEYINPUT7), .A3(new_n358), .A4(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT74), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n384), .A2(new_n386), .A3(new_n261), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT74), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(KEYINPUT3), .B2(G33), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n391), .A2(new_n392), .A3(new_n239), .A4(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT73), .ZN(new_n397));
  AOI21_X1  g0197(.A(G20), .B1(new_n330), .B2(new_n332), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n397), .B1(new_n398), .B2(KEYINPUT7), .ZN(new_n399));
  OAI211_X1 g0199(.A(KEYINPUT73), .B(new_n393), .C1(new_n293), .C2(G20), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n202), .B1(new_n396), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G58), .A2(G68), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n203), .A2(new_n205), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G20), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n268), .A2(G159), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n383), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n262), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n384), .A2(new_n386), .A3(G33), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n330), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n359), .A2(KEYINPUT7), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n202), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n330), .ZN(new_n414));
  XNOR2_X1  g0214(.A(KEYINPUT72), .B(KEYINPUT3), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(G33), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT7), .B1(new_n416), .B2(G20), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n407), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n409), .B1(new_n418), .B2(KEYINPUT16), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n408), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n266), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n280), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n278), .A2(new_n422), .B1(new_n274), .B2(new_n421), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  MUX2_X1   g0224(.A(G223), .B(G226), .S(G1698), .Z(new_n425));
  NAND2_X1  g0225(.A1(new_n416), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G87), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n427), .B(KEYINPUT75), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n299), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n344), .B1(new_n243), .B2(new_n290), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n303), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n289), .B1(G232), .B2(new_n291), .ZN(new_n433));
  XNOR2_X1  g0233(.A(KEYINPUT77), .B(G190), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n428), .B1(new_n416), .B2(new_n425), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n433), .B(new_n434), .C1(new_n299), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  AND4_X1   g0237(.A1(KEYINPUT78), .A2(new_n420), .A3(new_n424), .A4(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n423), .B1(new_n408), .B2(new_n419), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT78), .B1(new_n439), .B2(new_n437), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT17), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  AOI221_X4 g0241(.A(new_n423), .B1(new_n432), .B2(new_n436), .C1(new_n408), .C2(new_n419), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n442), .A2(KEYINPUT17), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n420), .A2(new_n424), .ZN(new_n445));
  OAI21_X1  g0245(.A(G169), .B1(new_n430), .B2(new_n431), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n433), .B(G179), .C1(new_n299), .C2(new_n435), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n445), .A2(KEYINPUT76), .A3(KEYINPUT18), .A4(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT18), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n439), .B2(new_n448), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n448), .B1(new_n420), .B2(new_n424), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT76), .B1(new_n454), .B2(KEYINPUT18), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n441), .B(new_n444), .C1(new_n453), .C2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n382), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT83), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n239), .A2(G33), .A3(G97), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT19), .ZN(new_n461));
  NAND3_X1  g0261(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n239), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(G97), .A2(G107), .ZN(new_n464));
  INV_X1    g0264(.A(G87), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n460), .A2(new_n461), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n410), .A2(G68), .A3(new_n239), .A4(new_n330), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n409), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n361), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(new_n274), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n459), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n460), .A2(new_n461), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n463), .A2(new_n466), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(new_n468), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n262), .ZN(new_n476));
  INV_X1    g0276(.A(new_n471), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(KEYINPUT83), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n277), .B1(G1), .B2(new_n261), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  XNOR2_X1  g0281(.A(new_n361), .B(KEYINPUT84), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G45), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(G1), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT81), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n279), .A2(G45), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT81), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n487), .A2(new_n490), .A3(G250), .A4(new_n286), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(new_n287), .B2(new_n488), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(G238), .A2(G1698), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n212), .B2(G1698), .ZN(new_n495));
  OR2_X1    g0295(.A1(KEYINPUT82), .A2(G116), .ZN(new_n496));
  NAND2_X1  g0296(.A1(KEYINPUT82), .A2(G116), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n416), .A2(new_n495), .B1(G33), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n493), .B1(new_n499), .B2(new_n299), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n378), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n495), .A2(new_n410), .A3(new_n330), .ZN(new_n502));
  INV_X1    g0302(.A(new_n498), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n502), .B1(new_n261), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n492), .B1(new_n504), .B2(new_n300), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n309), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n484), .A2(new_n501), .A3(new_n506), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n472), .A2(new_n478), .B1(G87), .B2(new_n481), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n500), .A2(G200), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n505), .A2(G190), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n274), .A2(new_n498), .ZN(new_n513));
  OR2_X1    g0313(.A1(new_n513), .A2(KEYINPUT85), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(KEYINPUT85), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n261), .A2(G97), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G283), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n357), .A2(new_n517), .A3(new_n358), .A4(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n496), .A2(G20), .A3(new_n497), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n262), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT20), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n262), .A2(KEYINPUT20), .A3(new_n519), .A4(new_n520), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n277), .B(G116), .C1(G1), .C2(new_n261), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n516), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(G257), .A2(G1698), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n214), .B2(G1698), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(new_n410), .A3(new_n330), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n370), .A2(G303), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n300), .ZN(new_n533));
  XNOR2_X1  g0333(.A(KEYINPUT5), .B(G41), .ZN(new_n534));
  INV_X1    g0334(.A(new_n231), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n534), .A2(new_n486), .B1(new_n535), .B2(new_n285), .ZN(new_n536));
  OR2_X1    g0336(.A1(KEYINPUT5), .A2(G41), .ZN(new_n537));
  NAND2_X1  g0337(.A1(KEYINPUT5), .A2(G41), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n488), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n536), .A2(G270), .B1(new_n342), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n378), .B1(new_n533), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n527), .A2(new_n541), .A3(KEYINPUT21), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n342), .A2(new_n539), .ZN(new_n543));
  INV_X1    g0343(.A(G270), .ZN(new_n544));
  INV_X1    g0344(.A(new_n538), .ZN(new_n545));
  NOR2_X1   g0345(.A1(KEYINPUT5), .A2(G41), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n486), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n286), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n543), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n299), .B1(new_n530), .B2(new_n531), .ZN(new_n550));
  NOR3_X1   g0350(.A1(new_n549), .A2(new_n550), .A3(new_n309), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n527), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n542), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(KEYINPUT21), .B1(new_n527), .B2(new_n541), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(G250), .A2(G1698), .ZN(new_n556));
  INV_X1    g0356(.A(G257), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n556), .B1(new_n557), .B2(G1698), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n558), .A2(new_n410), .A3(new_n330), .ZN(new_n559));
  INV_X1    g0359(.A(G294), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n559), .B1(new_n261), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n561), .A2(new_n300), .B1(G264), .B2(new_n536), .ZN(new_n562));
  AOI21_X1  g0362(.A(G169), .B1(new_n562), .B2(new_n543), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n536), .A2(G264), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n416), .A2(new_n558), .B1(G33), .B2(G294), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n564), .B(new_n543), .C1(new_n565), .C2(new_n299), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n566), .A2(G179), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  AND2_X1   g0368(.A1(KEYINPUT82), .A2(G116), .ZN(new_n569));
  NOR2_X1   g0369(.A1(KEYINPUT82), .A2(G116), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n263), .B(G33), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(KEYINPUT23), .A2(G107), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n237), .B2(new_n238), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n213), .A2(G20), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT23), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n571), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT87), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n571), .A2(new_n573), .A3(KEYINPUT87), .A4(new_n575), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n239), .A2(new_n293), .A3(G87), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT22), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n582), .A2(new_n465), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n410), .A2(new_n239), .A3(new_n330), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(KEYINPUT24), .B1(new_n580), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n586), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT24), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n578), .A2(new_n579), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n409), .B1(new_n587), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT25), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n274), .B2(G107), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n275), .A2(KEYINPUT25), .A3(new_n213), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n481), .A2(G107), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n568), .B1(new_n592), .B2(new_n597), .ZN(new_n598));
  NOR3_X1   g0398(.A1(new_n580), .A2(KEYINPUT24), .A3(new_n586), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n589), .B1(new_n588), .B2(new_n590), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n262), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n566), .A2(new_n303), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(G190), .B2(new_n566), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n603), .A3(new_n596), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n516), .A2(new_n525), .ZN(new_n605));
  OAI21_X1  g0405(.A(G200), .B1(new_n549), .B2(new_n550), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT86), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n605), .A2(new_n606), .A3(new_n607), .A4(new_n526), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n303), .B1(new_n533), .B2(new_n540), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT86), .B1(new_n527), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n434), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n533), .A2(new_n611), .A3(new_n540), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n608), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n555), .A2(new_n598), .A3(new_n604), .A4(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT80), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n275), .A2(new_n335), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(new_n480), .B2(new_n335), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT6), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n335), .A2(new_n213), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n618), .B1(new_n619), .B2(new_n464), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n213), .A2(KEYINPUT6), .A3(G97), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n622), .A2(new_n359), .B1(G77), .B2(new_n268), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n390), .A2(new_n395), .B1(new_n399), .B2(new_n400), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n623), .B1(new_n624), .B2(new_n213), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n617), .B1(new_n625), .B2(new_n262), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT79), .B1(new_n536), .B2(G257), .ZN(new_n627));
  AND4_X1   g0427(.A1(KEYINPUT79), .A2(new_n547), .A3(G257), .A4(new_n286), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n543), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT4), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n212), .A2(G1698), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n630), .B1(new_n411), .B2(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(KEYINPUT4), .A2(G244), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n330), .A2(new_n332), .A3(new_n634), .A4(new_n294), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n330), .A2(new_n332), .A3(G250), .A4(G1698), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n635), .A2(new_n636), .A3(new_n518), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n299), .B1(new_n633), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n378), .B1(new_n629), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT79), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n548), .B2(new_n557), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n536), .A2(KEYINPUT79), .A3(G257), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n641), .A2(new_n642), .B1(new_n342), .B2(new_n539), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT4), .B1(new_n416), .B2(new_n631), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n635), .A2(new_n636), .A3(new_n518), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n300), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n643), .A2(new_n646), .A3(new_n309), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n639), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n626), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n213), .B1(new_n396), .B2(new_n401), .ZN(new_n650));
  INV_X1    g0450(.A(new_n623), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n262), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n617), .ZN(new_n653));
  OAI21_X1  g0453(.A(G200), .B1(new_n629), .B2(new_n638), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n643), .A2(new_n646), .A3(G190), .ZN(new_n655));
  AND4_X1   g0455(.A1(new_n652), .A2(new_n653), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n615), .B1(new_n649), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n652), .A2(new_n653), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n658), .A2(new_n639), .A3(new_n647), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n626), .A2(new_n654), .A3(new_n655), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(KEYINPUT80), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  NOR4_X1   g0462(.A1(new_n458), .A2(new_n512), .A3(new_n614), .A4(new_n662), .ZN(G372));
  INV_X1    g0463(.A(new_n458), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT88), .B1(new_n499), .B2(new_n299), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT88), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n504), .A2(new_n666), .A3(new_n300), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n493), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n378), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n484), .A2(new_n670), .A3(new_n506), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(G200), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n508), .A2(new_n672), .A3(new_n510), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n671), .A2(new_n673), .A3(new_n649), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT89), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT89), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n674), .A2(new_n678), .A3(new_n675), .ZN(new_n679));
  INV_X1    g0479(.A(new_n512), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n680), .A2(KEYINPUT26), .A3(new_n649), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n677), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n671), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n555), .A2(new_n598), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n649), .A2(new_n656), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n684), .A2(new_n604), .A3(new_n685), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n671), .A2(new_n673), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n683), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n682), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n664), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n311), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n445), .A2(KEYINPUT18), .A3(new_n449), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n452), .ZN(new_n693));
  INV_X1    g0493(.A(new_n352), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n355), .B2(new_n381), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n441), .A2(new_n444), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n693), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n305), .A2(new_n308), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n691), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n690), .A2(new_n699), .ZN(G369));
  NAND2_X1  g0500(.A1(new_n239), .A2(new_n273), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT27), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n239), .A2(new_n703), .A3(new_n273), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n702), .A2(G213), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G343), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT90), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n526), .B2(new_n605), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n554), .B2(new_n553), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n555), .A2(new_n613), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n709), .B1(new_n710), .B2(new_n708), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G330), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT91), .ZN(new_n713));
  INV_X1    g0513(.A(new_n707), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n714), .B(new_n568), .C1(new_n592), .C2(new_n597), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n598), .A2(new_n604), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n707), .B1(new_n601), .B2(new_n596), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n713), .B(new_n715), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(KEYINPUT91), .A3(new_n568), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n712), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n718), .A2(new_n719), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n555), .A2(new_n714), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n598), .A2(new_n714), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n722), .A2(new_n725), .A3(new_n726), .ZN(G399));
  INV_X1    g0527(.A(new_n222), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G41), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n230), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n466), .A2(G116), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n731), .B(G1), .C1(G41), .C2(new_n728), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT92), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT28), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n687), .A2(KEYINPUT95), .A3(KEYINPUT26), .A4(new_n649), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n688), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT26), .B1(new_n680), .B2(new_n649), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT95), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(new_n674), .B2(new_n675), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  OAI211_X1 g0541(.A(KEYINPUT29), .B(new_n707), .C1(new_n737), .C2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n714), .B1(new_n682), .B2(new_n688), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n742), .B1(KEYINPUT29), .B2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(G330), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n564), .B1(new_n565), .B2(new_n299), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n500), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n533), .A2(G179), .A3(new_n540), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(KEYINPUT93), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n629), .A2(new_n638), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT93), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n533), .A2(new_n751), .A3(G179), .A4(new_n540), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n747), .A2(new_n749), .A3(new_n750), .A4(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT30), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n566), .B1(new_n629), .B2(new_n638), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(KEYINPUT94), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT94), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n566), .B(new_n758), .C1(new_n629), .C2(new_n638), .ZN(new_n759));
  AOI21_X1  g0559(.A(G179), .B1(new_n533), .B2(new_n540), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n757), .A2(new_n669), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  AND4_X1   g0561(.A1(new_n505), .A2(new_n562), .A3(new_n643), .A4(new_n646), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n762), .A2(KEYINPUT30), .A3(new_n752), .A4(new_n749), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n755), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n714), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT31), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n764), .A2(KEYINPUT31), .A3(new_n714), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n662), .A2(new_n614), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(new_n680), .A3(new_n707), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n745), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n744), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n735), .B1(new_n774), .B2(G1), .ZN(G364));
  NOR2_X1   g0575(.A1(new_n359), .A2(new_n272), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n279), .B1(new_n776), .B2(G45), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n729), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(new_n711), .B2(G330), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(G330), .B2(new_n711), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n293), .A2(new_n222), .ZN(new_n782));
  INV_X1    g0582(.A(G355), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n782), .A2(new_n783), .B1(G116), .B2(new_n222), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT96), .Z(new_n785));
  NAND2_X1  g0585(.A1(new_n230), .A2(new_n485), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n416), .A2(new_n728), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n253), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n788), .B1(new_n789), .B2(G45), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n785), .B1(new_n786), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n236), .B1(G20), .B2(new_n378), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G13), .A2(G33), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(G20), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n779), .B1(new_n791), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n303), .A2(G179), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n799), .A2(G20), .A3(G190), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT98), .Z(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G303), .ZN(new_n803));
  INV_X1    g0603(.A(G283), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n359), .A2(new_n354), .A3(new_n799), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n802), .A2(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(G179), .A2(G200), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n359), .A2(new_n354), .A3(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n806), .B1(G329), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n239), .B1(G190), .B2(new_n807), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n293), .B1(new_n812), .B2(G294), .ZN(new_n813));
  INV_X1    g0613(.A(G311), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n359), .A2(G179), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT97), .ZN(new_n816));
  AND3_X1   g0616(.A1(new_n816), .A2(new_n354), .A3(new_n303), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n810), .B(new_n813), .C1(new_n814), .C2(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n816), .A2(new_n354), .A3(G200), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(KEYINPUT33), .B(G317), .ZN(new_n822));
  AND3_X1   g0622(.A1(new_n816), .A2(new_n303), .A3(new_n611), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n821), .A2(new_n822), .B1(new_n823), .B2(G322), .ZN(new_n824));
  INV_X1    g0624(.A(G326), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n816), .A2(G200), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(new_n434), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n824), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n821), .A2(G68), .B1(new_n823), .B2(G58), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n211), .B2(new_n818), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n293), .B1(new_n800), .B2(new_n465), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n805), .A2(new_n213), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n832), .B(new_n833), .C1(G97), .C2(new_n812), .ZN(new_n834));
  INV_X1    g0634(.A(G159), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n808), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT32), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n834), .B(new_n837), .C1(new_n828), .C2(new_n226), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n819), .A2(new_n829), .B1(new_n831), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n798), .B1(new_n839), .B2(new_n792), .ZN(new_n840));
  INV_X1    g0640(.A(new_n795), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n711), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n781), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(G396));
  AND2_X1   g0644(.A1(new_n367), .A2(new_n714), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n380), .B1(new_n845), .B2(new_n376), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n381), .A2(new_n707), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n743), .B(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n779), .B1(new_n849), .B2(new_n773), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n773), .B2(new_n849), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n817), .A2(G159), .B1(new_n823), .B2(G143), .ZN(new_n852));
  INV_X1    g0652(.A(G137), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n852), .B1(new_n853), .B2(new_n828), .C1(new_n267), .C2(new_n820), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT34), .Z(new_n855));
  INV_X1    g0655(.A(G132), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n416), .B1(new_n808), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n805), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n812), .A2(G58), .B1(new_n858), .B2(G68), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n802), .B2(new_n226), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n855), .A2(new_n857), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n808), .A2(new_n814), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n805), .A2(new_n465), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n862), .B(new_n863), .C1(new_n801), .C2(G107), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n293), .B1(new_n812), .B2(G97), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n864), .B(new_n865), .C1(new_n804), .C2(new_n820), .ZN(new_n866));
  INV_X1    g0666(.A(new_n823), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n560), .A2(new_n867), .B1(new_n818), .B2(new_n503), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n866), .B(new_n868), .C1(G303), .C2(new_n827), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n792), .B1(new_n861), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n779), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n792), .A2(new_n793), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT99), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n871), .B1(new_n874), .B2(new_n211), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n870), .B(new_n875), .C1(new_n794), .C2(new_n848), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n851), .A2(new_n876), .ZN(G384));
  OR2_X1    g0677(.A1(new_n622), .A2(KEYINPUT35), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n622), .A2(KEYINPUT35), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(G116), .A3(new_n240), .A4(new_n879), .ZN(new_n880));
  XOR2_X1   g0680(.A(KEYINPUT100), .B(KEYINPUT36), .Z(new_n881));
  XNOR2_X1  g0681(.A(new_n880), .B(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n230), .A2(G77), .A3(new_n403), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(G50), .B2(new_n202), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n279), .A2(G13), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n847), .B(KEYINPUT101), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n743), .B2(new_n848), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n714), .A2(new_n322), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT102), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n352), .A2(new_n890), .A3(new_n355), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n352), .A2(KEYINPUT102), .A3(new_n355), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n889), .A2(new_n351), .A3(new_n349), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n889), .A2(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n888), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n405), .A2(new_n406), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n239), .A2(new_n393), .ZN(new_n899));
  OAI21_X1  g0699(.A(G68), .B1(new_n416), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n393), .B1(new_n411), .B2(new_n263), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n898), .B(KEYINPUT16), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n262), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n418), .A2(KEYINPUT16), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n424), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n705), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n420), .A2(new_n424), .A3(new_n437), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT78), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n439), .A2(KEYINPUT78), .A3(new_n437), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n443), .B1(new_n911), .B2(KEYINPUT17), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT76), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n692), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(new_n450), .A3(new_n452), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n906), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT37), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n439), .B2(new_n448), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n438), .A2(new_n918), .A3(new_n440), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n898), .B1(new_n624), .B2(new_n202), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n903), .B1(new_n383), .B2(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(KEYINPUT103), .B(new_n705), .C1(new_n921), .C2(new_n423), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT103), .ZN(new_n923));
  INV_X1    g0723(.A(new_n705), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n923), .B1(new_n439), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n905), .B1(new_n449), .B2(new_n705), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n909), .A2(new_n910), .A3(new_n927), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n919), .A2(new_n926), .B1(KEYINPUT37), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n897), .B1(new_n916), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n906), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n456), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n918), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n926), .A2(new_n909), .A3(new_n910), .A4(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n928), .A2(KEYINPUT37), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n932), .A2(KEYINPUT38), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n930), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n693), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n896), .A2(new_n938), .B1(new_n939), .B2(new_n924), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n916), .A2(new_n929), .A3(new_n897), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT38), .B1(new_n932), .B2(new_n936), .ZN(new_n942));
  OAI21_X1  g0742(.A(KEYINPUT39), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT104), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n938), .A2(KEYINPUT104), .A3(KEYINPUT39), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n926), .B1(new_n912), .B2(new_n693), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n442), .A2(new_n454), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n926), .A2(new_n948), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n926), .A2(new_n919), .B1(new_n949), .B2(KEYINPUT37), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n897), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT39), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n951), .A2(new_n952), .A3(new_n937), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(KEYINPUT105), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT105), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n951), .A2(new_n937), .A3(new_n955), .A4(new_n952), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n945), .A2(new_n946), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n694), .A2(new_n707), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n940), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n699), .B1(new_n744), .B2(new_n458), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NOR4_X1   g0761(.A1(new_n662), .A2(new_n614), .A3(new_n512), .A4(new_n714), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n767), .A2(new_n768), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n848), .B(new_n894), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n930), .B2(new_n937), .ZN(new_n965));
  INV_X1    g0765(.A(new_n926), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n696), .B2(new_n939), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n454), .B(new_n442), .C1(new_n922), .C2(new_n925), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n934), .B1(new_n968), .B2(new_n917), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT38), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n941), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n769), .A2(new_n771), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n972), .A2(KEYINPUT40), .A3(new_n848), .A4(new_n894), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n965), .A2(KEYINPUT40), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n458), .B1(new_n771), .B2(new_n769), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n745), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n976), .B2(new_n975), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n961), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n279), .B2(new_n776), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n961), .A2(new_n978), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n886), .B1(new_n980), .B2(new_n981), .ZN(G367));
  NAND2_X1  g0782(.A1(new_n249), .A2(new_n787), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n796), .B(new_n983), .C1(new_n222), .C2(new_n361), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n871), .B1(new_n984), .B2(KEYINPUT107), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(KEYINPUT107), .B2(new_n984), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n828), .A2(new_n814), .B1(new_n867), .B2(new_n803), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G294), .B2(new_n821), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n817), .A2(G283), .ZN(new_n989));
  INV_X1    g0789(.A(new_n800), .ZN(new_n990));
  AOI21_X1  g0790(.A(KEYINPUT46), .B1(new_n990), .B2(new_n498), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n416), .B(new_n991), .C1(G317), .C2(new_n809), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n805), .A2(new_n335), .ZN(new_n993));
  AND3_X1   g0793(.A1(new_n801), .A2(KEYINPUT46), .A3(G116), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n993), .B(new_n994), .C1(G107), .C2(new_n812), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n988), .A2(new_n989), .A3(new_n992), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n827), .A2(G143), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n202), .B2(new_n811), .C1(new_n267), .C2(new_n867), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT108), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n818), .A2(new_n226), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n805), .A2(new_n211), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n293), .B1(new_n201), .B2(new_n800), .C1(new_n808), .C2(new_n853), .ZN(new_n1003));
  NOR3_X1   g0803(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1000), .B(new_n1004), .C1(new_n835), .C2(new_n820), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n998), .A2(new_n999), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n996), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT47), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n986), .B1(new_n1008), .B2(new_n792), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n508), .A2(new_n707), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT106), .Z(new_n1011));
  OR2_X1    g0811(.A1(new_n1011), .A2(new_n687), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n671), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1009), .B1(new_n1015), .B2(new_n841), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n725), .A2(new_n726), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n685), .B1(new_n626), .B2(new_n707), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n659), .B2(new_n707), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT45), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1019), .B1(new_n725), .B2(new_n726), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT44), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n721), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n712), .B(new_n720), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(new_n724), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1022), .A2(new_n722), .A3(new_n1024), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1026), .A2(new_n774), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n774), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n729), .B(KEYINPUT41), .Z(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n778), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n723), .A2(new_n724), .A3(new_n1019), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1035), .A2(KEYINPUT42), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1018), .A2(new_n598), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n714), .B1(new_n1037), .B2(new_n659), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n1035), .B2(KEYINPUT42), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1036), .A2(new_n1039), .B1(KEYINPUT43), .B2(new_n1015), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1015), .A2(KEYINPUT43), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1040), .B(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n722), .A2(new_n1020), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1042), .B(new_n1043), .Z(new_n1044));
  OAI21_X1  g0844(.A(new_n1016), .B1(new_n1034), .B2(new_n1044), .ZN(G387));
  NOR2_X1   g0845(.A1(new_n774), .A2(new_n1028), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n774), .A2(new_n1028), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n729), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1046), .B1(new_n1048), .B2(KEYINPUT112), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(KEYINPUT112), .B2(new_n1048), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n782), .A2(new_n731), .B1(G107), .B2(new_n222), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n788), .B1(new_n246), .B2(G45), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n731), .B(new_n485), .C1(new_n202), .C2(new_n211), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT109), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  OAI21_X1  g0856(.A(KEYINPUT50), .B1(new_n266), .B2(G50), .ZN(new_n1057));
  OR3_X1    g0857(.A1(new_n266), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1051), .B1(new_n1052), .B2(new_n1059), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n779), .B1(new_n797), .B2(new_n1060), .C1(new_n723), .C2(new_n841), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n827), .A2(G159), .B1(new_n823), .B2(G50), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n416), .B1(new_n211), .B2(new_n800), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1063), .A2(new_n993), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n812), .A2(new_n482), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(new_n267), .C2(new_n808), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n817), .B2(G68), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1062), .B(new_n1067), .C1(new_n266), .C2(new_n820), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n811), .A2(new_n804), .B1(new_n560), .B2(new_n800), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n817), .A2(G303), .B1(new_n823), .B2(G317), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(KEYINPUT110), .B(G322), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1070), .B1(new_n814), .B2(new_n820), .C1(new_n828), .C2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT48), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1069), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n1073), .B2(new_n1072), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT49), .Z(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(KEYINPUT111), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n416), .B1(new_n809), .B2(G326), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(new_n503), .C2(new_n805), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1076), .A2(KEYINPUT111), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1068), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1061), .B1(new_n1081), .B2(new_n792), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n778), .B2(new_n1028), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1050), .A2(new_n1083), .ZN(G393));
  INV_X1    g0884(.A(new_n1029), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n722), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1085), .A2(new_n777), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1020), .A2(new_n795), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n796), .B1(new_n335), .B2(new_n222), .C1(new_n256), .C2(new_n788), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n779), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n827), .A2(G317), .B1(new_n823), .B2(G311), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT52), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n811), .A2(new_n503), .B1(new_n808), .B2(new_n1071), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n370), .B1(new_n800), .B2(new_n804), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n1093), .A2(new_n833), .A3(new_n1094), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1095), .B1(new_n803), .B2(new_n820), .C1(new_n818), .C2(new_n560), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n827), .A2(G150), .B1(new_n823), .B2(G159), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT51), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n811), .A2(new_n211), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n416), .B1(new_n202), .B2(new_n800), .C1(new_n805), .C2(new_n465), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1099), .B(new_n1100), .C1(G143), .C2(new_n809), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1101), .B1(new_n226), .B2(new_n820), .C1(new_n266), .C2(new_n818), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n1092), .A2(new_n1096), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1090), .B1(new_n1103), .B2(new_n792), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1087), .B1(new_n1088), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1047), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1106), .A2(new_n1030), .A3(new_n729), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1107), .ZN(G390));
  NAND2_X1  g0908(.A1(new_n772), .A2(new_n848), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n895), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n772), .A2(new_n848), .A3(new_n894), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n743), .A2(new_n848), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1112), .B1(new_n1113), .B2(new_n887), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n707), .B(new_n846), .C1(new_n737), .C2(new_n741), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1110), .A2(new_n847), .A3(new_n1111), .A4(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n664), .A2(new_n772), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n699), .B(new_n1118), .C1(new_n744), .C2(new_n458), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1111), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n895), .B1(new_n1115), .B2(new_n847), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n951), .A2(new_n937), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n958), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n958), .B1(new_n888), .B2(new_n895), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1122), .B(new_n1126), .C1(new_n957), .C2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n954), .A2(new_n956), .ZN(new_n1129));
  AOI21_X1  g0929(.A(KEYINPUT104), .B1(new_n938), .B2(KEYINPUT39), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n946), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1129), .B(new_n1127), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1126), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1111), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1121), .B1(new_n1128), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n1122), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1132), .A2(new_n1111), .A3(new_n1133), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1119), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1135), .A2(new_n1140), .A3(new_n729), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1128), .A2(new_n1134), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n957), .A2(new_n793), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n873), .A2(new_n421), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n827), .A2(G128), .B1(new_n823), .B2(G132), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT113), .Z(new_n1146));
  NAND2_X1  g0946(.A1(new_n821), .A2(G137), .ZN(new_n1147));
  XOR2_X1   g0947(.A(KEYINPUT54), .B(G143), .Z(new_n1148));
  NAND2_X1  g0948(.A1(new_n817), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT53), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n990), .B2(G150), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n800), .A2(KEYINPUT53), .A3(new_n267), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1151), .A2(new_n370), .A3(new_n1152), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n811), .A2(new_n835), .B1(new_n805), .B2(new_n226), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(G125), .B2(new_n809), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1147), .A2(new_n1149), .A3(new_n1153), .A4(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n827), .A2(G283), .B1(new_n817), .B2(G97), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n213), .B2(new_n820), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n823), .A2(G116), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n293), .B1(new_n858), .B2(G68), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n808), .A2(new_n560), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1161), .B(new_n1099), .C1(new_n801), .C2(G87), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1159), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n1146), .A2(new_n1156), .B1(new_n1158), .B2(new_n1163), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n871), .B(new_n1144), .C1(new_n1164), .C2(new_n792), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1142), .A2(new_n778), .B1(new_n1143), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1141), .A2(new_n1166), .ZN(G378));
  AOI22_X1  g0967(.A1(G97), .A2(new_n821), .B1(new_n817), .B2(new_n482), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT114), .Z(new_n1169));
  AOI22_X1  g0969(.A1(new_n812), .A2(G68), .B1(new_n990), .B2(G77), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n805), .A2(new_n201), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n416), .A2(G41), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(G283), .C2(new_n809), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1170), .B(new_n1173), .C1(new_n867), .C2(new_n213), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G116), .B2(new_n827), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1169), .A2(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT115), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1177), .A2(KEYINPUT58), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(KEYINPUT58), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1172), .B(new_n226), .C1(G33), .C2(G41), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n827), .A2(G125), .B1(G150), .B2(new_n812), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT116), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n821), .A2(G132), .B1(new_n823), .B2(G128), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n817), .A2(G137), .B1(new_n990), .B2(new_n1148), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1182), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n858), .A2(G159), .ZN(new_n1190));
  AOI211_X1 g0990(.A(G33), .B(G41), .C1(new_n809), .C2(G124), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .A4(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n792), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n871), .B1(new_n226), .B2(new_n872), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n282), .A2(new_n705), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n312), .B(new_n1197), .Z(new_n1198));
  XNOR2_X1  g0998(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1198), .B(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1196), .B1(new_n793), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1202), .B1(new_n974), .B2(new_n745), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n964), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n938), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT40), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1124), .A2(KEYINPUT40), .A3(new_n1205), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1208), .A2(new_n1201), .A3(G330), .A4(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1204), .A2(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n940), .B(KEYINPUT118), .C1(new_n957), .C2(new_n958), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(KEYINPUT117), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1204), .A2(KEYINPUT117), .A3(new_n1210), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(KEYINPUT118), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1211), .A2(new_n1213), .B1(new_n1215), .B2(new_n959), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1203), .B1(new_n1216), .B2(new_n778), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1119), .B1(new_n1142), .B2(new_n1117), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n959), .A2(new_n1211), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n959), .A2(new_n1211), .ZN(new_n1220));
  OAI21_X1  g1020(.A(KEYINPUT57), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n729), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1140), .A2(new_n1120), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT57), .B1(new_n1223), .B2(new_n1216), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1217), .B1(new_n1222), .B2(new_n1224), .ZN(G375));
  INV_X1    g1025(.A(new_n1117), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n1119), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1227), .A2(new_n1033), .A3(new_n1121), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1065), .B1(new_n803), .B2(new_n808), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(G97), .B2(new_n801), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1002), .A2(new_n293), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(new_n828), .C2(new_n560), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n498), .A2(new_n821), .B1(new_n817), .B2(G107), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT119), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1232), .B(new_n1234), .C1(G283), .C2(new_n823), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1235), .A2(KEYINPUT120), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n828), .A2(new_n856), .B1(new_n867), .B2(new_n853), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n821), .B2(new_n1148), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n817), .A2(G150), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1171), .A2(new_n411), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n802), .A2(new_n835), .B1(new_n226), .B2(new_n811), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(G128), .B2(new_n809), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .A4(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1235), .B2(KEYINPUT120), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n792), .B1(new_n1236), .B2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n871), .B1(new_n874), .B2(new_n202), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1245), .B(new_n1246), .C1(new_n794), .C2(new_n894), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n1226), .B2(new_n777), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1228), .A2(new_n1249), .ZN(G381));
  XOR2_X1   g1050(.A(G375), .B(KEYINPUT121), .Z(new_n1251));
  AND2_X1   g1051(.A1(new_n1141), .A2(new_n1166), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1253));
  INV_X1    g1053(.A(G384), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1253), .A2(new_n1254), .A3(new_n1249), .A4(new_n1228), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1050), .A2(new_n1083), .A3(new_n843), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1255), .A2(G387), .A3(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1251), .A2(new_n1252), .A3(new_n1257), .ZN(G407));
  INV_X1    g1058(.A(G213), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1259), .A2(G343), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(G378), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1251), .A2(new_n1262), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1263), .B(KEYINPUT122), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1065(.A(KEYINPUT127), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(G387), .A2(new_n1253), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1256), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n843), .B1(new_n1050), .B2(new_n1083), .ZN(new_n1269));
  OAI21_X1  g1069(.A(KEYINPUT124), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(G393), .A2(G396), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT124), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(new_n1272), .A3(new_n1256), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G390), .B(new_n1016), .C1(new_n1034), .C2(new_n1044), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1267), .A2(new_n1270), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n1267), .A2(new_n1274), .B1(new_n1270), .B2(new_n1273), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1266), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1267), .A2(new_n1274), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(KEYINPUT127), .A3(new_n1275), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1283));
  XOR2_X1   g1083(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1284));
  OAI211_X1 g1084(.A(G378), .B(new_n1217), .C1(new_n1222), .C2(new_n1224), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1223), .A2(new_n1216), .A3(new_n1033), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n959), .B(new_n1211), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1203), .B1(new_n1287), .B2(new_n778), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1252), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1260), .B1(new_n1285), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT60), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1227), .B1(new_n1292), .B2(new_n1139), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1226), .A2(KEYINPUT60), .A3(new_n1119), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(new_n729), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1249), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1254), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1295), .A2(G384), .A3(new_n1249), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1284), .B1(new_n1291), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT125), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1285), .A2(new_n1290), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1302), .B1(new_n1303), .B2(new_n1261), .ZN(new_n1304));
  AOI211_X1 g1104(.A(KEYINPUT125), .B(new_n1260), .C1(new_n1285), .C2(new_n1290), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1300), .A2(KEYINPUT62), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1301), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1260), .A2(G2897), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(new_n1299), .B(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1310), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT61), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1283), .B1(new_n1308), .B2(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1312), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1291), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1315), .B1(new_n1316), .B2(new_n1310), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT63), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1299), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1306), .A2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT63), .B1(new_n1291), .B2(new_n1300), .ZN(new_n1321));
  OR2_X1    g1121(.A1(new_n1321), .A2(KEYINPUT123), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(KEYINPUT123), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1317), .A2(new_n1320), .A3(new_n1322), .A4(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1314), .A2(new_n1324), .ZN(G405));
  NAND2_X1  g1125(.A1(G375), .A2(new_n1252), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1285), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(new_n1327), .B(new_n1300), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(new_n1283), .B(new_n1328), .ZN(G402));
endmodule


