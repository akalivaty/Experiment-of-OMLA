//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n816, new_n817, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT1), .ZN(new_n205));
  XNOR2_X1  g004(.A(G127gat), .B(G134gat), .ZN(new_n206));
  INV_X1    g005(.A(G120gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n207), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n208));
  NAND4_X1  g007(.A1(new_n204), .A2(new_n205), .A3(new_n206), .A4(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n206), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(KEYINPUT1), .B2(new_n202), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT73), .ZN(new_n214));
  XNOR2_X1  g013(.A(G141gat), .B(G148gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n216), .B1(G155gat), .B2(G162gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n214), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(G155gat), .B(G162gat), .Z(new_n219));
  AND2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n218), .A2(new_n219), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(KEYINPUT74), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n213), .B1(new_n223), .B2(KEYINPUT3), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n220), .A2(new_n221), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT75), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT75), .B1(new_n222), .B2(KEYINPUT3), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n225), .A2(new_n213), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT4), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n222), .A2(new_n212), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n235), .A2(KEYINPUT4), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G225gat), .A2(G233gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n231), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT5), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n225), .B(KEYINPUT74), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n232), .B1(new_n241), .B2(new_n213), .ZN(new_n242));
  INV_X1    g041(.A(new_n238), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n239), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G1gat), .B(G29gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT0), .ZN(new_n247));
  XNOR2_X1  g046(.A(G57gat), .B(G85gat), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n247), .B(new_n248), .Z(new_n249));
  INV_X1    g048(.A(KEYINPUT76), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n250), .B1(new_n234), .B2(new_n236), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n232), .A2(new_n233), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n235), .A2(KEYINPUT4), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(KEYINPUT76), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n255), .A2(new_n231), .A3(new_n240), .A4(new_n238), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n245), .A2(new_n249), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT77), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n245), .A2(new_n256), .ZN(new_n259));
  INV_X1    g058(.A(new_n249), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT6), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT77), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n245), .A2(new_n263), .A3(new_n249), .A4(new_n256), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n258), .A2(new_n261), .A3(new_n262), .A4(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT78), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n264), .A2(new_n262), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n268), .A2(KEYINPUT78), .A3(new_n261), .A4(new_n258), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n249), .B1(new_n245), .B2(new_n256), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT6), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n267), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(G183gat), .A2(G190gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT24), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n274), .A2(KEYINPUT64), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT64), .B1(new_n274), .B2(new_n275), .ZN(new_n277));
  OAI221_X1 g076(.A(new_n273), .B1(G183gat), .B2(G190gat), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT65), .B(G176gat), .ZN(new_n279));
  INV_X1    g078(.A(G169gat), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n280), .A2(KEYINPUT23), .ZN(new_n281));
  INV_X1    g080(.A(G176gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT23), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n279), .A2(new_n281), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n278), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n273), .B1(G183gat), .B2(G190gat), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n288), .B1(new_n275), .B2(new_n274), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n281), .A2(new_n282), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n285), .A2(new_n283), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT25), .ZN(new_n292));
  OAI22_X1  g091(.A1(new_n287), .A2(KEYINPUT25), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT26), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n283), .A2(new_n294), .A3(new_n284), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n295), .B(new_n274), .C1(new_n294), .C2(new_n283), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT68), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n297), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT28), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT66), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n301), .B(KEYINPUT67), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT27), .B(G183gat), .ZN(new_n303));
  INV_X1    g102(.A(G190gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  OR2_X1    g105(.A1(new_n302), .A2(new_n305), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n298), .A2(new_n299), .A3(new_n306), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G226gat), .A2(G233gat), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n311), .B(KEYINPUT72), .Z(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n309), .B1(KEYINPUT29), .B2(new_n312), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G211gat), .B(G218gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n320));
  OR2_X1    g119(.A1(G197gat), .A2(G204gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(G197gat), .A2(G204gat), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n319), .B(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n316), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n314), .A2(new_n324), .A3(new_n315), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G8gat), .B(G36gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(G64gat), .B(G92gat), .ZN(new_n330));
  XOR2_X1   g129(.A(new_n329), .B(new_n330), .Z(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n326), .A2(new_n327), .A3(new_n331), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(KEYINPUT30), .A3(new_n334), .ZN(new_n335));
  OR3_X1    g134(.A1(new_n328), .A2(KEYINPUT30), .A3(new_n332), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n272), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT80), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT79), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT3), .B1(new_n324), .B2(new_n341), .ZN(new_n342));
  OAI211_X1 g141(.A(G228gat), .B(G233gat), .C1(new_n241), .C2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT29), .B1(new_n228), .B2(new_n229), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n344), .A2(new_n324), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n340), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G228gat), .A2(G233gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n324), .A2(new_n341), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(new_n227), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n347), .B1(new_n349), .B2(new_n223), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n350), .B(KEYINPUT79), .C1(new_n324), .C2(new_n344), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G22gat), .ZN(new_n353));
  OAI22_X1  g152(.A1(new_n344), .A2(new_n324), .B1(new_n225), .B2(new_n342), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n347), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n353), .B1(new_n352), .B2(new_n355), .ZN(new_n358));
  OAI21_X1  g157(.A(G78gat), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n358), .ZN(new_n360));
  INV_X1    g159(.A(G78gat), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(new_n361), .A3(new_n356), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT31), .B(G50gat), .ZN(new_n363));
  INV_X1    g162(.A(G106gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n359), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n365), .B1(new_n359), .B2(new_n362), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n339), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n365), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n361), .B1(new_n360), .B2(new_n356), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n357), .A2(new_n358), .A3(G78gat), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n359), .A2(new_n362), .A3(new_n365), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(KEYINPUT80), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n338), .A2(new_n368), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT86), .ZN(new_n376));
  INV_X1    g175(.A(new_n337), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n238), .B1(new_n255), .B2(new_n231), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT39), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n235), .B1(new_n223), .B2(new_n212), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT82), .B1(new_n381), .B2(new_n238), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT82), .ZN(new_n383));
  NOR3_X1   g182(.A1(new_n242), .A2(new_n383), .A3(new_n243), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n380), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT81), .B(KEYINPUT39), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n378), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n385), .A2(KEYINPUT40), .A3(new_n249), .A4(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT40), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n384), .A2(new_n382), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n390), .A2(new_n378), .A3(new_n379), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n387), .A2(new_n249), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n389), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n259), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n245), .A2(KEYINPUT83), .A3(new_n256), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(new_n260), .A3(new_n396), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n377), .A2(new_n388), .A3(new_n393), .A4(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n372), .A2(new_n398), .A3(new_n373), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n270), .A2(KEYINPUT85), .A3(KEYINPUT6), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT85), .B1(new_n270), .B2(KEYINPUT6), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n397), .A2(new_n268), .A3(new_n258), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n328), .A2(KEYINPUT37), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT37), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n326), .A2(new_n327), .A3(new_n405), .ZN(new_n406));
  XOR2_X1   g205(.A(KEYINPUT84), .B(KEYINPUT38), .Z(new_n407));
  NAND4_X1  g206(.A1(new_n404), .A2(new_n406), .A3(new_n332), .A4(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n334), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n331), .B1(new_n328), .B2(KEYINPUT37), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n407), .B1(new_n410), .B2(new_n406), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n402), .A2(new_n403), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n376), .B1(new_n399), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n366), .A2(new_n367), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n402), .A2(new_n403), .A3(new_n412), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n415), .A2(KEYINPUT86), .A3(new_n416), .A4(new_n398), .ZN(new_n417));
  INV_X1    g216(.A(G227gat), .ZN(new_n418));
  INV_X1    g217(.A(G233gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n310), .A2(new_n213), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n309), .A2(new_n212), .ZN(new_n421));
  AOI211_X1 g220(.A(new_n418), .B(new_n419), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT32), .ZN(new_n424));
  XOR2_X1   g223(.A(G71gat), .B(G99gat), .Z(new_n425));
  XNOR2_X1  g224(.A(G15gat), .B(G43gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n424), .B(new_n427), .C1(KEYINPUT33), .C2(new_n422), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n420), .B(new_n421), .C1(new_n418), .C2(new_n419), .ZN(new_n429));
  XOR2_X1   g228(.A(new_n429), .B(KEYINPUT34), .Z(new_n430));
  INV_X1    g229(.A(KEYINPUT70), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n427), .A2(new_n431), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT33), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n423), .B(KEYINPUT32), .C1(new_n432), .C2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n428), .A2(new_n430), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n430), .B1(new_n428), .B2(new_n435), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT36), .ZN(new_n440));
  INV_X1    g239(.A(new_n438), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n436), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT36), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n375), .A2(new_n414), .A3(new_n417), .A4(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n439), .A2(new_n372), .A3(new_n373), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT35), .B1(new_n447), .B2(new_n338), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT35), .B1(new_n402), .B2(new_n403), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n415), .A2(new_n337), .A3(new_n439), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(G229gat), .A2(G233gat), .ZN(new_n453));
  XOR2_X1   g252(.A(new_n453), .B(KEYINPUT13), .Z(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G15gat), .B(G22gat), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT16), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n457), .A2(G1gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n459), .B1(G1gat), .B2(new_n456), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT90), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n461), .B1(new_n456), .B2(G1gat), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(G8gat), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(G8gat), .ZN(new_n464));
  OAI221_X1 g263(.A(new_n459), .B1(new_n461), .B2(new_n464), .C1(G1gat), .C2(new_n456), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT87), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g269(.A(KEYINPUT87), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT14), .ZN(new_n472));
  INV_X1    g271(.A(G29gat), .ZN(new_n473));
  INV_X1    g272(.A(G36gat), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n470), .A2(new_n471), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT88), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n470), .A2(KEYINPUT88), .A3(new_n471), .A4(new_n475), .ZN(new_n479));
  NAND2_X1  g278(.A1(G29gat), .A2(G36gat), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(G50gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(G43gat), .ZN(new_n483));
  INV_X1    g282(.A(G43gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(G50gat), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n485), .A3(KEYINPUT15), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n480), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT15), .B1(new_n483), .B2(new_n485), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n475), .A2(KEYINPUT89), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n475), .A2(KEYINPUT89), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n468), .A3(new_n492), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n481), .A2(new_n487), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n467), .A2(new_n494), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n476), .A2(new_n477), .B1(G29gat), .B2(G36gat), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n486), .B1(new_n496), .B2(new_n479), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n490), .A2(new_n493), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n466), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n455), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n467), .B1(new_n494), .B2(KEYINPUT17), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT17), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n497), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n453), .B(new_n499), .C1(new_n501), .C2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT18), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n500), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G113gat), .B(G141gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(G197gat), .ZN(new_n508));
  XOR2_X1   g307(.A(KEYINPUT11), .B(G169gat), .Z(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n510), .B(KEYINPUT12), .Z(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n494), .A2(KEYINPUT17), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n502), .B1(new_n497), .B2(new_n498), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n514), .A3(new_n467), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n515), .A2(KEYINPUT18), .A3(new_n453), .A4(new_n499), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n506), .A2(new_n512), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n512), .B1(new_n506), .B2(new_n516), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT91), .ZN(new_n521));
  XNOR2_X1  g320(.A(G57gat), .B(G64gat), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G71gat), .B(G78gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT21), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G231gat), .A2(G233gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(G127gat), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n467), .B1(new_n527), .B2(new_n526), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT92), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n531), .B(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(G155gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(G183gat), .B(G211gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n534), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G99gat), .B(G106gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(G85gat), .A2(G92gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT7), .ZN(new_n542));
  INV_X1    g341(.A(G92gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT93), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT93), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(G92gat), .ZN(new_n546));
  INV_X1    g345(.A(G85gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT94), .ZN(new_n549));
  INV_X1    g348(.A(G99gat), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT8), .B1(new_n550), .B2(new_n364), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n549), .B1(new_n548), .B2(new_n551), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n540), .B(new_n542), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n548), .A2(new_n551), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT94), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n540), .B1(new_n559), .B2(new_n542), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n513), .B(new_n514), .C1(new_n555), .C2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n542), .B1(new_n552), .B2(new_n553), .ZN(new_n562));
  INV_X1    g361(.A(new_n540), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n564), .B(new_n554), .C1(new_n497), .C2(new_n498), .ZN(new_n565));
  NAND3_X1  g364(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n565), .A2(KEYINPUT95), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT95), .B1(new_n565), .B2(new_n566), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n561), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G190gat), .B(G218gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n570), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n572), .B(new_n561), .C1(new_n567), .C2(new_n568), .ZN(new_n573));
  XNOR2_X1  g372(.A(G134gat), .B(G162gat), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n571), .A2(KEYINPUT96), .A3(new_n573), .A4(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT96), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n580), .A2(new_n576), .B1(new_n571), .B2(new_n573), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n539), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(G230gat), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(new_n419), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n526), .B1(new_n560), .B2(new_n555), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT10), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n524), .B(new_n525), .Z(new_n588));
  NAND3_X1  g387(.A1(new_n564), .A2(new_n588), .A3(new_n554), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT97), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT97), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n586), .A2(new_n592), .A3(new_n589), .A4(new_n587), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n564), .A2(new_n588), .A3(KEYINPUT10), .A4(new_n554), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n585), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n585), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n597), .B1(new_n586), .B2(new_n589), .ZN(new_n598));
  XOR2_X1   g397(.A(G120gat), .B(G148gat), .Z(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT98), .ZN(new_n600));
  XNOR2_X1  g399(.A(G176gat), .B(G204gat), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n600), .B(new_n601), .Z(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  OR3_X1    g402(.A1(new_n596), .A2(new_n598), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n603), .B1(new_n596), .B2(new_n598), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n583), .A2(new_n606), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n452), .A2(new_n520), .A3(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n272), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(G1gat), .ZN(G1324gat));
  INV_X1    g410(.A(new_n608), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n457), .A2(new_n464), .ZN(new_n613));
  NOR2_X1   g412(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n614));
  NOR4_X1   g413(.A1(new_n612), .A2(new_n337), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n464), .B1(new_n608), .B2(new_n377), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT42), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n617), .B1(KEYINPUT42), .B2(new_n615), .ZN(G1325gat));
  OAI21_X1  g417(.A(G15gat), .B1(new_n612), .B2(new_n445), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n442), .A2(G15gat), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n619), .B1(new_n612), .B2(new_n620), .ZN(G1326gat));
  NAND2_X1  g420(.A1(new_n368), .A2(new_n374), .ZN(new_n622));
  OR3_X1    g421(.A1(new_n612), .A2(KEYINPUT99), .A3(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(KEYINPUT99), .B1(new_n612), .B2(new_n622), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT43), .B(G22gat), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n625), .B1(new_n623), .B2(new_n624), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(G1327gat));
  INV_X1    g427(.A(new_n539), .ZN(new_n629));
  INV_X1    g428(.A(new_n606), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n517), .A2(new_n518), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n504), .A2(new_n505), .ZN(new_n634));
  INV_X1    g433(.A(new_n500), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(new_n516), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n511), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n506), .A2(new_n512), .A3(new_n516), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT100), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n631), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT44), .ZN(new_n643));
  INV_X1    g442(.A(new_n582), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n643), .B1(new_n452), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(new_n578), .B2(new_n581), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n580), .A2(new_n576), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n571), .A2(new_n573), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n650), .A2(KEYINPUT101), .A3(new_n577), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(KEYINPUT44), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n654), .B1(new_n446), .B2(new_n451), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n609), .B(new_n642), .C1(new_n645), .C2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(G29gat), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n631), .A2(new_n582), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n272), .A2(G29gat), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n452), .A2(new_n520), .A3(new_n658), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT45), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1328gat));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n452), .A2(new_n520), .A3(new_n658), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n337), .A2(G36gat), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(KEYINPUT103), .Z(new_n669));
  NAND3_X1  g468(.A1(new_n666), .A2(new_n665), .A3(new_n667), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n670), .B(KEYINPUT104), .Z(new_n671));
  NAND2_X1  g470(.A1(new_n452), .A2(new_n653), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n582), .B1(new_n446), .B2(new_n451), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n672), .B1(new_n673), .B2(new_n643), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(new_n377), .A3(new_n642), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(G36gat), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n669), .A2(new_n671), .A3(new_n676), .ZN(G1329gat));
  INV_X1    g476(.A(new_n445), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n678), .B(new_n642), .C1(new_n645), .C2(new_n655), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(G43gat), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n666), .A2(new_n484), .A3(new_n439), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT47), .B1(new_n682), .B2(KEYINPUT105), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT105), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT47), .ZN(new_n685));
  AOI211_X1 g484(.A(new_n684), .B(new_n685), .C1(new_n680), .C2(new_n681), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n683), .A2(new_n686), .ZN(G1330gat));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n622), .A2(G50gat), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n452), .A2(new_n520), .A3(new_n658), .A4(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT48), .ZN(new_n691));
  INV_X1    g490(.A(new_n415), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n674), .A2(new_n692), .A3(new_n642), .ZN(new_n693));
  AOI211_X1 g492(.A(new_n688), .B(new_n691), .C1(new_n693), .C2(G50gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n690), .B(KEYINPUT106), .ZN(new_n695));
  INV_X1    g494(.A(new_n622), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n696), .B(new_n642), .C1(new_n645), .C2(new_n655), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n695), .B1(new_n698), .B2(new_n482), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT48), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n691), .B1(new_n693), .B2(G50gat), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(KEYINPUT107), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n694), .B1(new_n701), .B2(new_n703), .ZN(G1331gat));
  NOR3_X1   g503(.A1(new_n583), .A2(new_n630), .A3(new_n640), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n452), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n272), .B(KEYINPUT108), .Z(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g509(.A(new_n337), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT109), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n706), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT110), .ZN(new_n714));
  NOR2_X1   g513(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1333gat));
  INV_X1    g515(.A(G71gat), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n706), .A2(new_n717), .A3(new_n439), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n706), .A2(new_n678), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(new_n717), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n696), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g522(.A1(new_n539), .A2(new_n640), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n673), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT51), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n725), .A2(KEYINPUT51), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n730), .A2(new_n547), .A3(new_n609), .A4(new_n606), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n539), .A2(new_n630), .A3(new_n640), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n674), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733), .B2(new_n272), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(new_n734), .ZN(G1336gat));
  NAND3_X1  g534(.A1(new_n674), .A2(new_n377), .A3(new_n732), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n544), .A2(new_n546), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n630), .A2(new_n337), .A3(G92gat), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT111), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n728), .A2(new_n729), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n738), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n727), .A2(KEYINPUT112), .ZN(new_n744));
  XOR2_X1   g543(.A(new_n725), .B(new_n744), .Z(new_n745));
  AOI22_X1  g544(.A1(new_n745), .A2(new_n740), .B1(new_n736), .B2(new_n737), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n743), .B1(new_n746), .B2(new_n742), .ZN(G1337gat));
  NAND4_X1  g546(.A1(new_n730), .A2(new_n550), .A3(new_n439), .A4(new_n606), .ZN(new_n748));
  OAI21_X1  g547(.A(G99gat), .B1(new_n733), .B2(new_n445), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(G1338gat));
  OAI21_X1  g549(.A(G106gat), .B1(new_n733), .B2(new_n415), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT53), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n415), .A2(G106gat), .A3(new_n630), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n728), .A2(new_n729), .A3(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n751), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n753), .B(KEYINPUT113), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n674), .A2(new_n696), .A3(new_n732), .ZN(new_n757));
  AOI22_X1  g556(.A1(new_n745), .A2(new_n756), .B1(new_n757), .B2(G106gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n755), .B1(new_n758), .B2(new_n752), .ZN(G1339gat));
  AOI21_X1  g558(.A(new_n453), .B1(new_n515), .B2(new_n499), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n495), .A2(new_n499), .A3(new_n455), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n510), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n638), .A2(new_n762), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n647), .A2(new_n651), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT54), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n602), .B1(new_n596), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n595), .A2(new_n585), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n594), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(KEYINPUT114), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n594), .A2(new_n771), .A3(new_n768), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n595), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n591), .B2(new_n593), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT54), .B1(new_n775), .B2(new_n585), .ZN(new_n776));
  OAI211_X1 g575(.A(KEYINPUT55), .B(new_n766), .C1(new_n773), .C2(new_n776), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n777), .A2(new_n604), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT115), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780));
  AOI211_X1 g579(.A(KEYINPUT114), .B(new_n767), .C1(new_n591), .C2(new_n593), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n771), .B1(new_n594), .B2(new_n768), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n776), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n594), .A2(new_n595), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n784), .A2(new_n765), .A3(new_n597), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n603), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n780), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n764), .A2(new_n778), .A3(new_n779), .A4(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(new_n604), .A3(new_n777), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n647), .A2(new_n651), .A3(new_n763), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT115), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n787), .A2(new_n640), .A3(new_n604), .A4(new_n777), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n606), .A2(new_n763), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n652), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n794), .B1(new_n793), .B2(new_n795), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n792), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n629), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n607), .A2(new_n641), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n707), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n447), .A2(new_n377), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(G113gat), .B1(new_n805), .B2(new_n640), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n696), .B1(new_n800), .B2(new_n801), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n272), .A2(new_n377), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n439), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(G113gat), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n809), .A2(new_n810), .A3(new_n519), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n806), .A2(new_n811), .ZN(G1340gat));
  AOI21_X1  g611(.A(G120gat), .B1(new_n805), .B2(new_n606), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n809), .A2(new_n207), .A3(new_n630), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(G1341gat));
  OR3_X1    g614(.A1(new_n804), .A2(G127gat), .A3(new_n629), .ZN(new_n816));
  OAI21_X1  g615(.A(G127gat), .B1(new_n809), .B2(new_n629), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1342gat));
  NOR3_X1   g617(.A1(new_n804), .A2(G134gat), .A3(new_n582), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n820), .A2(KEYINPUT56), .ZN(new_n821));
  OAI21_X1  g620(.A(G134gat), .B1(new_n809), .B2(new_n582), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(KEYINPUT56), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(G1343gat));
  NAND2_X1  g623(.A1(new_n445), .A2(new_n808), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n696), .A2(KEYINPUT57), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n783), .B2(new_n786), .ZN(new_n829));
  OAI211_X1 g628(.A(KEYINPUT117), .B(new_n766), .C1(new_n773), .C2(new_n776), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n780), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n778), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT118), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n831), .A2(new_n778), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(new_n520), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n644), .B1(new_n836), .B2(new_n795), .ZN(new_n837));
  INV_X1    g636(.A(new_n792), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n629), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n827), .B1(new_n839), .B2(new_n801), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n800), .A2(new_n801), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT57), .B1(new_n841), .B2(new_n692), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n826), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G141gat), .B1(new_n843), .B2(new_n519), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n678), .A2(new_n377), .A3(new_n415), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n802), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n519), .A2(G141gat), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT121), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n850), .A2(KEYINPUT121), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n844), .A2(new_n849), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n640), .B(new_n826), .C1(new_n840), .C2(new_n842), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n854), .A2(KEYINPUT119), .A3(G141gat), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT119), .B1(new_n854), .B2(G141gat), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n847), .A2(KEYINPUT120), .A3(new_n848), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n858));
  INV_X1    g657(.A(new_n848), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n846), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n855), .A2(new_n856), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n853), .B1(new_n862), .B2(new_n850), .ZN(G1344gat));
  INV_X1    g662(.A(G148gat), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n847), .A2(new_n864), .A3(new_n606), .ZN(new_n865));
  INV_X1    g664(.A(new_n843), .ZN(new_n866));
  AOI211_X1 g665(.A(KEYINPUT59), .B(new_n864), .C1(new_n866), .C2(new_n606), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n696), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n644), .A2(new_n763), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n789), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n629), .B1(new_n837), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n607), .A2(new_n519), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n870), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n869), .B1(new_n841), .B2(new_n692), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n630), .B1(new_n825), .B2(KEYINPUT122), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n877), .B(new_n878), .C1(KEYINPUT122), .C2(new_n825), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n868), .B1(new_n879), .B2(G148gat), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n865), .B1(new_n867), .B2(new_n880), .ZN(G1345gat));
  OAI21_X1  g680(.A(G155gat), .B1(new_n843), .B2(new_n629), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n629), .A2(G155gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n846), .B2(new_n883), .ZN(G1346gat));
  AOI21_X1  g683(.A(G162gat), .B1(new_n847), .B2(new_n644), .ZN(new_n885));
  INV_X1    g684(.A(new_n652), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n886), .A2(G162gat), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n885), .B1(new_n866), .B2(new_n887), .ZN(G1347gat));
  NOR2_X1   g687(.A1(new_n708), .A2(new_n337), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n807), .A3(new_n439), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n890), .A2(new_n280), .A3(new_n519), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n609), .B1(new_n800), .B2(new_n801), .ZN(new_n892));
  AND4_X1   g691(.A1(new_n377), .A2(new_n892), .A3(new_n415), .A4(new_n439), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n640), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n891), .B1(new_n280), .B2(new_n894), .ZN(G1348gat));
  NOR3_X1   g694(.A1(new_n890), .A2(new_n279), .A3(new_n630), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n893), .A2(new_n606), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n282), .B2(new_n897), .ZN(G1349gat));
  NAND3_X1  g697(.A1(new_n893), .A2(new_n303), .A3(new_n539), .ZN(new_n899));
  OAI21_X1  g698(.A(G183gat), .B1(new_n890), .B2(new_n629), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g700(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n902));
  XOR2_X1   g701(.A(new_n901), .B(new_n902), .Z(G1350gat));
  NAND3_X1  g702(.A1(new_n893), .A2(new_n304), .A3(new_n886), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n890), .A2(new_n582), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n905), .A2(new_n304), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n906), .A2(new_n907), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n904), .B1(new_n909), .B2(new_n910), .ZN(G1351gat));
  NAND3_X1  g710(.A1(new_n445), .A2(new_n377), .A3(new_n692), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT124), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n892), .ZN(new_n914));
  OR3_X1    g713(.A1(new_n914), .A2(G197gat), .A3(new_n641), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n889), .A2(new_n520), .A3(new_n445), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n841), .A2(new_n692), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(KEYINPUT57), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n873), .A2(new_n874), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n918), .B(new_n919), .C1(new_n920), .C2(new_n870), .ZN(new_n921));
  OAI21_X1  g720(.A(KEYINPUT125), .B1(new_n875), .B2(new_n876), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n916), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n923), .A2(KEYINPUT126), .ZN(new_n924));
  OAI21_X1  g723(.A(G197gat), .B1(new_n923), .B2(KEYINPUT126), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n915), .B1(new_n924), .B2(new_n925), .ZN(G1352gat));
  INV_X1    g725(.A(G204gat), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n606), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT62), .B1(new_n914), .B2(new_n928), .ZN(new_n929));
  OR3_X1    g728(.A1(new_n914), .A2(KEYINPUT62), .A3(new_n928), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n889), .A2(new_n445), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n931), .B1(new_n921), .B2(new_n922), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n932), .A2(new_n606), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n929), .B(new_n930), .C1(new_n933), .C2(new_n927), .ZN(G1353gat));
  OR3_X1    g733(.A1(new_n914), .A2(G211gat), .A3(new_n629), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n877), .A2(new_n445), .A3(new_n539), .A4(new_n889), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n936), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT63), .B1(new_n936), .B2(G211gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(G1354gat));
  INV_X1    g738(.A(new_n914), .ZN(new_n940));
  AOI21_X1  g739(.A(G218gat), .B1(new_n940), .B2(new_n886), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n644), .A2(G218gat), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n941), .B1(new_n932), .B2(new_n942), .ZN(G1355gat));
endmodule


