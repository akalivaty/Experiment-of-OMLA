//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G210), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT27), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G101), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT67), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT67), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G119), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n196), .A3(G116), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n193), .A2(G116), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G113), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT2), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G113), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n200), .A2(new_n202), .A3(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT67), .B(G119), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n198), .B1(new_n206), .B2(G116), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n202), .A2(new_n204), .ZN(new_n208));
  AOI21_X1  g022(.A(KEYINPUT68), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n197), .A2(new_n208), .A3(KEYINPUT68), .A4(new_n199), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n205), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G137), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G134), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT11), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(KEYINPUT64), .A3(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n214), .A2(G134), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n216), .B1(new_n215), .B2(KEYINPUT64), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n220), .A2(G131), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G131), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n215), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n214), .A2(KEYINPUT65), .A3(G134), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n223), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G146), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G143), .ZN(new_n229));
  INV_X1    g043(.A(G143), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G146), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(new_n233), .A3(G128), .ZN(new_n234));
  INV_X1    g048(.A(G128), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n229), .B(new_n231), .C1(KEYINPUT1), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  OR3_X1    g051(.A1(new_n222), .A2(new_n227), .A3(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(G131), .B1(new_n220), .B2(new_n221), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n215), .A2(KEYINPUT64), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT11), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n241), .A2(new_n217), .A3(new_n223), .A4(new_n219), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT0), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n229), .B(new_n231), .C1(new_n245), .C2(new_n235), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n235), .ZN(new_n247));
  NOR2_X1   g061(.A1(KEYINPUT0), .A2(G128), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(G143), .B(G146), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n246), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n232), .B1(new_n248), .B2(new_n247), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(KEYINPUT69), .A3(new_n246), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n213), .B(new_n238), .C1(new_n244), .C2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT28), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n222), .A2(new_n237), .A3(new_n227), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n239), .A2(new_n242), .B1(new_n254), .B2(new_n246), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n212), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n259), .B1(new_n258), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n192), .B1(new_n260), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT30), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n266), .B1(new_n261), .B2(new_n262), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT66), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n238), .B(KEYINPUT30), .C1(new_n257), .C2(new_n244), .ZN(new_n270));
  OAI211_X1 g084(.A(KEYINPUT66), .B(new_n266), .C1(new_n261), .C2(new_n262), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n269), .A2(new_n212), .A3(new_n270), .A4(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT31), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n272), .A2(new_n273), .A3(new_n258), .A4(new_n191), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n265), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n272), .A2(new_n258), .A3(new_n191), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT31), .ZN(new_n277));
  AOI21_X1  g091(.A(G902), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n279));
  INV_X1    g093(.A(G472), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n278), .A2(new_n279), .A3(KEYINPUT32), .A4(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n277), .A2(new_n274), .A3(new_n265), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n282), .A2(KEYINPUT32), .A3(new_n280), .A4(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT70), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n282), .A2(new_n280), .A3(new_n283), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT32), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n238), .B1(new_n257), .B2(new_n244), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n212), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n258), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n260), .B1(KEYINPUT28), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n192), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(G902), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  OR2_X1    g109(.A1(new_n260), .A2(new_n264), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n293), .B1(new_n296), .B2(new_n192), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n272), .A2(new_n258), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n299), .A2(new_n191), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n295), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G472), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n281), .A2(new_n285), .A3(new_n288), .A4(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(G214), .B1(G237), .B2(G902), .ZN(new_n304));
  XOR2_X1   g118(.A(new_n304), .B(KEYINPUT78), .Z(new_n305));
  OAI21_X1  g119(.A(G210), .B1(G237), .B2(G902), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT4), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT75), .ZN(new_n309));
  INV_X1    g123(.A(G107), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n309), .B1(new_n310), .B2(G104), .ZN(new_n311));
  INV_X1    g125(.A(G104), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(KEYINPUT75), .A3(G107), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT3), .B1(new_n312), .B2(G107), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n310), .A3(G104), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(KEYINPUT76), .B1(new_n314), .B2(new_n318), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n311), .A2(new_n315), .A3(new_n317), .A4(new_n313), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n308), .B(G101), .C1(new_n319), .C2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G101), .ZN(new_n324));
  AND4_X1   g138(.A1(new_n311), .A2(new_n315), .A3(new_n317), .A4(new_n313), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT76), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n320), .A2(new_n321), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n314), .A2(new_n318), .A3(new_n324), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT4), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n212), .B(new_n323), .C1(new_n328), .C2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n197), .A2(new_n199), .A3(new_n208), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT68), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n210), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n312), .A2(G107), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n310), .A2(G104), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n324), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n338), .B1(new_n325), .B2(new_n324), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT5), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n206), .A2(new_n340), .A3(G116), .ZN(new_n341));
  OAI211_X1 g155(.A(G113), .B(new_n341), .C1(new_n200), .C2(new_n340), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n335), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n331), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(G110), .B(G122), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  XOR2_X1   g160(.A(KEYINPUT80), .B(KEYINPUT6), .Z(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT81), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n345), .B1(new_n331), .B2(new_n343), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(KEYINPUT81), .A3(new_n347), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n331), .A2(new_n343), .A3(new_n345), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT79), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n331), .A2(new_n356), .A3(new_n343), .A4(new_n345), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT6), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n351), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n246), .B(G125), .C1(new_n249), .C2(new_n250), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT82), .ZN(new_n363));
  INV_X1    g177(.A(G125), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n237), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT82), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n254), .A2(new_n366), .A3(G125), .A4(new_n246), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n363), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G224), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(G953), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n368), .B(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n353), .A2(new_n361), .A3(new_n371), .ZN(new_n372));
  XOR2_X1   g186(.A(new_n345), .B(KEYINPUT8), .Z(new_n373));
  OAI21_X1  g187(.A(new_n342), .B1(new_n209), .B2(new_n211), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n336), .A2(new_n337), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G101), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n376), .B1(new_n320), .B2(G101), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n373), .B1(new_n378), .B2(new_n343), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT7), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n370), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n362), .ZN(new_n383));
  AOI21_X1  g197(.A(G125), .B1(new_n234), .B2(new_n236), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(new_n368), .B2(new_n382), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n379), .A2(KEYINPUT83), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT83), .ZN(new_n388));
  INV_X1    g202(.A(new_n373), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n335), .A2(new_n339), .A3(new_n342), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n339), .B1(new_n335), .B2(new_n342), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n381), .B1(new_n365), .B2(new_n362), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n363), .A2(new_n365), .A3(new_n367), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n394), .B2(new_n381), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n388), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n387), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(G902), .B1(new_n397), .B2(new_n358), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n372), .B1(KEYINPUT84), .B2(new_n398), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n355), .A2(new_n357), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT83), .B1(new_n379), .B2(new_n386), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n392), .A2(new_n395), .A3(new_n388), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n283), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT84), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n307), .B1(new_n399), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n405), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n398), .A2(KEYINPUT84), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n408), .A2(new_n409), .A3(new_n306), .A4(new_n372), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n305), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G469), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(new_n283), .ZN(new_n413));
  XNOR2_X1  g227(.A(G110), .B(G140), .ZN(new_n414));
  INV_X1    g228(.A(G953), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n415), .A2(G227), .ZN(new_n416));
  XOR2_X1   g230(.A(new_n414), .B(new_n416), .Z(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n323), .B(new_n256), .C1(new_n328), .C2(new_n330), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n234), .A2(new_n236), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n339), .A2(KEYINPUT10), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT10), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n377), .B2(new_n237), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n419), .A2(new_n424), .A3(new_n244), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n244), .B1(new_n419), .B2(new_n424), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n418), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n329), .A2(new_n376), .B1(new_n236), .B2(new_n234), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n377), .A2(new_n237), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n243), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT12), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g246(.A(KEYINPUT12), .B(new_n243), .C1(new_n428), .C2(new_n429), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n419), .A2(new_n424), .A3(new_n244), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n435), .A3(new_n417), .ZN(new_n436));
  AOI21_X1  g250(.A(G902), .B1(new_n427), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n413), .B1(new_n437), .B2(new_n412), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n434), .A2(new_n435), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n418), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT77), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n435), .A2(new_n441), .A3(new_n417), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n419), .A2(new_n424), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n243), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n441), .B1(new_n435), .B2(new_n417), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n440), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n438), .B1(new_n447), .B2(new_n412), .ZN(new_n448));
  XOR2_X1   g262(.A(KEYINPUT9), .B(G234), .Z(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G221), .B1(new_n450), .B2(G902), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT74), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G475), .ZN(new_n455));
  XNOR2_X1  g269(.A(G125), .B(G140), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n228), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(KEYINPUT72), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(new_n228), .B2(new_n456), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n460));
  AOI21_X1  g274(.A(G143), .B1(new_n187), .B2(G214), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(new_n223), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT18), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT18), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n462), .B1(new_n465), .B2(new_n223), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n459), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n456), .A2(KEYINPUT16), .ZN(new_n468));
  OR3_X1    g282(.A1(new_n364), .A2(KEYINPUT16), .A3(G140), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(G146), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(G146), .B1(new_n468), .B2(new_n469), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n463), .A2(KEYINPUT17), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n462), .B(new_n223), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n473), .B(new_n474), .C1(new_n475), .C2(KEYINPUT17), .ZN(new_n476));
  XNOR2_X1  g290(.A(G113), .B(G122), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT85), .B(G104), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n477), .B(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n467), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  XOR2_X1   g295(.A(new_n456), .B(KEYINPUT19), .Z(new_n482));
  OAI211_X1 g296(.A(new_n475), .B(new_n470), .C1(G146), .C2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n479), .B1(new_n467), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n455), .B(new_n283), .C1(new_n481), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT20), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n467), .A2(new_n483), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n480), .B1(new_n487), .B2(new_n479), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT20), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n488), .A2(new_n489), .A3(new_n455), .A4(new_n283), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n479), .B1(new_n467), .B2(new_n476), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n283), .B1(new_n481), .B2(new_n491), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n486), .A2(new_n490), .B1(G475), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(G234), .A2(G237), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(G952), .A3(new_n415), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(G902), .A3(G953), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT21), .B(G898), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n496), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G122), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G116), .ZN(new_n503));
  INV_X1    g317(.A(G116), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G122), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(new_n505), .A3(new_n310), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT88), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n506), .B(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n235), .A2(G143), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n235), .A2(G143), .ZN(new_n511));
  OAI21_X1  g325(.A(G134), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n230), .A2(G128), .ZN(new_n513));
  INV_X1    g327(.A(G134), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n509), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT14), .B1(new_n502), .B2(G116), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n517), .B1(new_n504), .B2(G122), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n505), .A2(KEYINPUT14), .ZN(new_n519));
  OAI21_X1  g333(.A(G107), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n508), .A2(new_n516), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n511), .B1(KEYINPUT13), .B2(new_n509), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n522), .A2(KEYINPUT86), .B1(KEYINPUT13), .B2(new_n511), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT13), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n513), .B1(new_n510), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT86), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n514), .B1(new_n523), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n503), .A2(new_n505), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G107), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT87), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n530), .A2(new_n506), .B1(new_n515), .B2(new_n531), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n515), .A2(new_n531), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n521), .B1(new_n528), .B2(new_n534), .ZN(new_n535));
  XOR2_X1   g349(.A(KEYINPUT71), .B(G217), .Z(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n537), .A2(new_n450), .A3(G953), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n521), .B(new_n538), .C1(new_n528), .C2(new_n534), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n283), .ZN(new_n543));
  INV_X1    g357(.A(G478), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(KEYINPUT15), .ZN(new_n545));
  XOR2_X1   g359(.A(new_n543), .B(new_n545), .Z(new_n546));
  NAND3_X1  g360(.A1(new_n493), .A2(new_n501), .A3(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n454), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n537), .B1(G234), .B2(new_n283), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT23), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n194), .B(new_n196), .C1(new_n551), .C2(G128), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(G128), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n235), .A2(KEYINPUT23), .A3(G119), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G110), .ZN(new_n556));
  NOR2_X1   g370(.A1(G119), .A2(G128), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n194), .A2(new_n196), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n557), .B1(new_n558), .B2(G128), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT24), .B(G110), .ZN(new_n560));
  OAI221_X1 g374(.A(new_n556), .B1(new_n559), .B2(new_n560), .C1(new_n471), .C2(new_n472), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n560), .ZN(new_n562));
  INV_X1    g376(.A(G110), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n552), .A2(new_n563), .A3(new_n553), .A4(new_n554), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n458), .A2(new_n565), .A3(new_n470), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT22), .B(G137), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n415), .A2(G221), .A3(G234), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n561), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n569), .B1(new_n561), .B2(new_n566), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n283), .B(new_n550), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT73), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n283), .B1(new_n570), .B2(new_n571), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT25), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g391(.A(KEYINPUT25), .B(new_n283), .C1(new_n570), .C2(new_n571), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n550), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n303), .A2(new_n411), .A3(new_n548), .A4(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(G101), .ZN(G3));
  NAND2_X1  g396(.A1(new_n282), .A2(new_n283), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G472), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n286), .ZN(new_n585));
  INV_X1    g399(.A(new_n580), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n585), .A2(new_n454), .A3(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(new_n587), .B(KEYINPUT89), .Z(new_n588));
  NAND3_X1  g402(.A1(new_n542), .A2(new_n544), .A3(new_n283), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT91), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n542), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT33), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n542), .A2(new_n590), .A3(KEYINPUT33), .ZN(new_n594));
  AOI21_X1  g408(.A(G902), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n589), .B1(new_n595), .B2(new_n544), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT92), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT92), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n589), .B(new_n598), .C1(new_n595), .C2(new_n544), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n493), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n305), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n358), .A2(new_n360), .B1(new_n350), .B2(new_n352), .ZN(new_n604));
  AOI22_X1  g418(.A1(new_n405), .A2(new_n404), .B1(new_n604), .B2(new_n371), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n306), .B1(new_n605), .B2(new_n409), .ZN(new_n606));
  AND4_X1   g420(.A1(new_n306), .A2(new_n408), .A3(new_n409), .A4(new_n372), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n603), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT90), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT90), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n411), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NOR4_X1   g427(.A1(new_n588), .A2(new_n500), .A3(new_n602), .A4(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT34), .B(G104), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  INV_X1    g430(.A(new_n546), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n493), .A2(new_n617), .ZN(new_n618));
  NOR4_X1   g432(.A1(new_n588), .A2(new_n500), .A3(new_n613), .A4(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(KEYINPUT93), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT35), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(new_n310), .ZN(G9));
  INV_X1    g436(.A(new_n585), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n561), .A2(new_n566), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n569), .A2(KEYINPUT36), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n626), .A2(new_n283), .A3(new_n550), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n579), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n411), .A2(new_n548), .A3(new_n623), .A4(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT37), .B(G110), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G12));
  XOR2_X1   g446(.A(new_n495), .B(KEYINPUT94), .Z(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(G900), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n634), .B1(new_n635), .B2(new_n498), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n618), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n638), .A2(new_n454), .A3(new_n628), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n407), .A2(new_n410), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n610), .B1(new_n640), .B2(new_n603), .ZN(new_n641));
  AOI211_X1 g455(.A(KEYINPUT90), .B(new_n305), .C1(new_n407), .C2(new_n410), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n303), .B(new_n639), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT95), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n612), .A2(KEYINPUT95), .A3(new_n303), .A4(new_n639), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G128), .ZN(G30));
  INV_X1    g462(.A(new_n454), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n636), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n653));
  OR2_X1    g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n640), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n652), .A2(new_n653), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n493), .A2(new_n546), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n603), .A3(new_n628), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT99), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n654), .A2(new_n656), .A3(new_n657), .A4(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n280), .B1(new_n291), .B2(new_n192), .ZN(new_n662));
  AOI22_X1  g476(.A1(new_n662), .A2(new_n276), .B1(G472), .B2(G902), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n663), .B(KEYINPUT97), .Z(new_n664));
  NAND4_X1  g478(.A1(new_n664), .A2(new_n281), .A3(new_n285), .A4(new_n288), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT98), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n230), .ZN(G45));
  AOI211_X1 g482(.A(new_n493), .B(new_n636), .C1(new_n597), .C2(new_n599), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n669), .B1(new_n641), .B2(new_n642), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT102), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n303), .A2(new_n629), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n673), .B(new_n669), .C1(new_n641), .C2(new_n642), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n671), .A2(new_n649), .A3(new_n672), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G146), .ZN(G48));
  AOI21_X1  g490(.A(new_n417), .B1(new_n444), .B2(new_n435), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n434), .A2(new_n435), .A3(new_n417), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n412), .B(new_n283), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT103), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n437), .A2(new_n412), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n437), .A2(KEYINPUT103), .A3(new_n412), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n453), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n283), .B1(new_n677), .B2(new_n678), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(G469), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(KEYINPUT103), .A3(new_n679), .ZN(new_n689));
  OR3_X1    g503(.A1(new_n437), .A2(KEYINPUT103), .A3(new_n412), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(KEYINPUT104), .A3(new_n453), .ZN(new_n692));
  AND4_X1   g506(.A1(new_n303), .A2(new_n686), .A3(new_n580), .A4(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n602), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n612), .A2(new_n693), .A3(new_n501), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT41), .B(G113), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G15));
  INV_X1    g511(.A(new_n618), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n612), .A2(new_n693), .A3(new_n501), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  INV_X1    g514(.A(new_n547), .ZN(new_n701));
  AOI21_X1  g515(.A(KEYINPUT104), .B1(new_n691), .B2(new_n453), .ZN(new_n702));
  AOI211_X1 g516(.A(new_n685), .B(new_n452), .C1(new_n689), .C2(new_n690), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n612), .A2(new_n701), .A3(new_n672), .A4(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT105), .B(G119), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G21));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n708), .B1(new_n574), .B2(new_n579), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n577), .A2(new_n578), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n549), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n572), .B(KEYINPUT73), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n712), .A3(KEYINPUT106), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n274), .B1(new_n292), .B2(new_n191), .ZN(new_n715));
  INV_X1    g529(.A(new_n277), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n280), .B(new_n283), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n584), .A2(new_n714), .A3(new_n717), .ZN(new_n718));
  NOR4_X1   g532(.A1(new_n702), .A2(new_n703), .A3(new_n718), .A4(new_n500), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n612), .A2(new_n719), .A3(new_n658), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  INV_X1    g535(.A(new_n636), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n600), .A2(new_n601), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n584), .A2(new_n629), .A3(new_n717), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n704), .B(new_n725), .C1(new_n641), .C2(new_n642), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G125), .ZN(G27));
  NAND3_X1  g541(.A1(new_n288), .A2(new_n302), .A3(new_n284), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n669), .A2(new_n728), .A3(new_n714), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n407), .A2(new_n603), .A3(new_n410), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT107), .B1(new_n445), .B2(new_n446), .ZN(new_n731));
  INV_X1    g545(.A(new_n446), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n733), .A3(new_n444), .A4(new_n442), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n731), .A2(new_n734), .A3(G469), .A4(new_n440), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n438), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT108), .B1(new_n736), .B2(new_n453), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n738));
  AOI211_X1 g552(.A(new_n738), .B(new_n452), .C1(new_n735), .C2(new_n438), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n729), .A2(new_n730), .A3(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT42), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n736), .A2(new_n453), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n738), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n736), .A2(KEYINPUT108), .A3(new_n453), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n730), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n746), .A2(new_n747), .A3(new_n303), .A4(new_n580), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n669), .A2(new_n742), .ZN(new_n749));
  OAI22_X1  g563(.A1(new_n741), .A2(new_n742), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(new_n223), .ZN(G33));
  NOR2_X1   g565(.A1(new_n748), .A2(new_n638), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n514), .ZN(G36));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n600), .A2(new_n493), .ZN(new_n755));
  XOR2_X1   g569(.A(new_n755), .B(KEYINPUT43), .Z(new_n756));
  NOR2_X1   g570(.A1(new_n623), .A2(new_n628), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT109), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n757), .A2(KEYINPUT109), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n754), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n731), .A2(new_n734), .A3(KEYINPUT45), .A4(new_n440), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n412), .B1(new_n447), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n413), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n765), .A2(KEYINPUT46), .ZN(new_n766));
  AOI22_X1  g580(.A1(new_n765), .A2(KEYINPUT46), .B1(new_n412), .B2(new_n437), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n452), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n768), .A2(new_n651), .ZN(new_n769));
  INV_X1    g583(.A(new_n760), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n770), .A2(KEYINPUT44), .A3(new_n756), .A4(new_n758), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n761), .A2(new_n747), .A3(new_n769), .A4(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G137), .ZN(G39));
  XNOR2_X1  g587(.A(new_n768), .B(KEYINPUT47), .ZN(new_n774));
  NOR4_X1   g588(.A1(new_n303), .A2(new_n730), .A3(new_n723), .A4(new_n580), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n777), .A2(KEYINPUT110), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(KEYINPUT110), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G140), .ZN(G42));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n782));
  AND4_X1   g596(.A1(new_n695), .A2(new_n699), .A3(new_n705), .A4(new_n720), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n725), .A2(new_n747), .A3(new_n746), .ZN(new_n784));
  NOR4_X1   g598(.A1(new_n601), .A2(new_n628), .A3(new_n617), .A4(new_n636), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n747), .A2(new_n303), .A3(new_n649), .A4(new_n785), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n784), .B(new_n786), .C1(new_n748), .C2(new_n638), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n618), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n493), .A2(new_n617), .A3(KEYINPUT113), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n500), .B1(new_n791), .B2(new_n602), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n411), .A3(new_n587), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n581), .A3(new_n630), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n750), .A2(new_n787), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n783), .A2(new_n795), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n743), .A2(new_n629), .A3(new_n636), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n612), .A2(new_n665), .A3(new_n658), .A4(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n675), .A2(new_n647), .A3(new_n726), .A4(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n726), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(new_n645), .B2(new_n646), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(KEYINPUT52), .A3(new_n675), .A4(new_n798), .ZN(new_n804));
  AOI211_X1 g618(.A(new_n782), .B(new_n796), .C1(new_n801), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT114), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n801), .A2(new_n804), .ZN(new_n807));
  INV_X1    g621(.A(new_n796), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n782), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n807), .A2(KEYINPUT53), .A3(new_n808), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n806), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT54), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n810), .A2(new_n816), .A3(new_n811), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT53), .B1(new_n807), .B2(new_n808), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(new_n805), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT115), .B1(new_n821), .B2(new_n816), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n815), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n756), .A2(new_n634), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n718), .ZN(new_n825));
  INV_X1    g639(.A(new_n704), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n656), .A2(new_n826), .A3(new_n603), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT50), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT117), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n828), .A2(new_n831), .A3(KEYINPUT50), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n828), .A2(KEYINPUT50), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n826), .A2(new_n730), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n580), .A2(new_n836), .A3(new_n496), .A4(new_n666), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n600), .A2(new_n601), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n836), .A2(new_n634), .A3(new_n756), .ZN(new_n839));
  INV_X1    g653(.A(new_n724), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n837), .A2(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n825), .A2(new_n747), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT116), .ZN(new_n843));
  INV_X1    g657(.A(new_n691), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n453), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n774), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n835), .A2(KEYINPUT51), .A3(new_n841), .A4(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n728), .A2(new_n714), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n839), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT48), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n613), .A2(new_n826), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n825), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n851), .A2(G952), .A3(new_n415), .A4(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n694), .B2(new_n837), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n848), .A2(new_n855), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n833), .A2(new_n834), .B1(new_n846), .B2(new_n843), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT51), .B1(new_n857), .B2(new_n841), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  OAI22_X1  g673(.A1(new_n823), .A2(new_n859), .B1(G952), .B2(G953), .ZN(new_n860));
  INV_X1    g674(.A(new_n755), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(new_n603), .A3(new_n453), .A4(new_n714), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(KEYINPUT111), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n862), .A2(KEYINPUT111), .ZN(new_n864));
  AOI211_X1 g678(.A(new_n863), .B(new_n864), .C1(KEYINPUT49), .C2(new_n844), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT112), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT49), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n656), .B1(new_n869), .B2(new_n691), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n867), .A2(new_n666), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n860), .A2(new_n871), .ZN(G75));
  NOR2_X1   g686(.A1(new_n821), .A2(new_n283), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT56), .B1(new_n873), .B2(G210), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n604), .B(new_n371), .ZN(new_n875));
  XOR2_X1   g689(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n876));
  XNOR2_X1  g690(.A(new_n875), .B(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n415), .A2(G952), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n880), .B1(new_n874), .B2(new_n877), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n878), .A2(new_n881), .ZN(G51));
  NOR2_X1   g696(.A1(new_n677), .A2(new_n678), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n413), .B(KEYINPUT57), .Z(new_n884));
  OAI21_X1  g698(.A(KEYINPUT54), .B1(new_n820), .B2(new_n805), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n884), .B1(new_n817), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n883), .B1(new_n886), .B2(KEYINPUT119), .ZN(new_n887));
  INV_X1    g701(.A(new_n884), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n820), .A2(new_n805), .A3(KEYINPUT54), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n816), .B1(new_n810), .B2(new_n811), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n887), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n762), .A2(new_n764), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT120), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n873), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n879), .B1(new_n894), .B2(new_n897), .ZN(G54));
  INV_X1    g712(.A(new_n488), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n810), .A2(new_n811), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(G902), .ZN(new_n901));
  NAND2_X1  g715(.A1(KEYINPUT58), .A2(G475), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n902), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n900), .A2(G902), .A3(new_n488), .A4(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n903), .A2(new_n880), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n903), .A2(KEYINPUT121), .A3(new_n880), .A4(new_n905), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(G60));
  NOR2_X1   g724(.A1(new_n889), .A2(new_n890), .ZN(new_n911));
  NAND2_X1  g725(.A1(G478), .A2(G902), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT59), .Z(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n593), .ZN(new_n915));
  INV_X1    g729(.A(new_n594), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n880), .B1(new_n911), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n823), .A2(new_n914), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n915), .A2(new_n916), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(G63));
  NAND2_X1  g735(.A1(G217), .A2(G902), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT60), .Z(new_n923));
  NAND2_X1  g737(.A1(new_n900), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n570), .A2(new_n571), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n879), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n924), .A2(new_n925), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n900), .A2(new_n626), .A3(new_n923), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n929), .A2(new_n880), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n928), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n926), .B(new_n930), .C1(new_n927), .C2(KEYINPUT61), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(G66));
  INV_X1    g749(.A(new_n783), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(new_n794), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n938), .A2(KEYINPUT123), .A3(new_n415), .ZN(new_n939));
  OAI21_X1  g753(.A(G953), .B1(new_n499), .B2(new_n369), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT123), .B1(new_n938), .B2(new_n415), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(G898), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n604), .B1(new_n944), .B2(G953), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n943), .B(new_n945), .ZN(G69));
  NAND3_X1  g760(.A1(new_n269), .A2(new_n271), .A3(new_n270), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(new_n482), .Z(new_n948));
  AND2_X1   g762(.A1(new_n791), .A2(new_n602), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n949), .A2(new_n652), .A3(new_n730), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n950), .A2(new_n303), .A3(new_n580), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n780), .A2(new_n772), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n803), .A2(new_n675), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n953), .A2(new_n667), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n952), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n948), .B1(new_n958), .B2(G953), .ZN(new_n959));
  INV_X1    g773(.A(new_n769), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n612), .A2(new_n658), .A3(new_n849), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n772), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(new_n778), .B2(new_n779), .ZN(new_n963));
  INV_X1    g777(.A(new_n953), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n750), .A2(new_n752), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT125), .Z(new_n966));
  NAND4_X1  g780(.A1(new_n963), .A2(new_n415), .A3(new_n964), .A4(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n948), .B1(G900), .B2(G953), .ZN(new_n968));
  AOI21_X1  g782(.A(KEYINPUT124), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n959), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n415), .B1(G227), .B2(G900), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(G72));
  AND2_X1   g786(.A1(new_n958), .A2(new_n937), .ZN(new_n973));
  NAND2_X1  g787(.A1(G472), .A2(G902), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT63), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n298), .B(new_n191), .C1(new_n973), .C2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n975), .ZN(new_n977));
  INV_X1    g791(.A(new_n276), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n814), .B(new_n977), .C1(new_n978), .C2(new_n300), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n963), .A2(new_n964), .A3(new_n937), .A4(new_n966), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n980), .A2(KEYINPUT126), .A3(new_n977), .ZN(new_n981));
  AOI21_X1  g795(.A(KEYINPUT126), .B1(new_n980), .B2(new_n977), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n299), .B(new_n192), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  AND4_X1   g797(.A1(new_n880), .A2(new_n976), .A3(new_n979), .A4(new_n983), .ZN(G57));
endmodule


