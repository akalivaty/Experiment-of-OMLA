//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n851, new_n852, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961;
  INV_X1    g000(.A(KEYINPUT24), .ZN(new_n202));
  INV_X1    g001(.A(G183gat), .ZN(new_n203));
  INV_X1    g002(.A(G190gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT68), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT68), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(G183gat), .B2(G190gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n209));
  NAND4_X1  g008(.A1(new_n205), .A2(new_n206), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT69), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G169gat), .ZN(new_n213));
  INV_X1    g012(.A(G176gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT23), .ZN(new_n215));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT67), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n213), .A2(new_n214), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(KEYINPUT65), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n222));
  NOR2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(KEYINPUT23), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT67), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n215), .A2(new_n226), .A3(new_n216), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n218), .A2(new_n225), .A3(KEYINPUT25), .A4(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT70), .B1(new_n212), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT25), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n205), .A2(KEYINPUT64), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n232), .B(new_n202), .C1(new_n203), .C2(new_n204), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n203), .A2(new_n204), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n231), .A2(new_n233), .A3(new_n234), .A4(new_n209), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n217), .B1(new_n224), .B2(new_n221), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AOI211_X1 g037(.A(KEYINPUT66), .B(new_n217), .C1(new_n224), .C2(new_n221), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n230), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n228), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT70), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n206), .A2(new_n208), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n243), .A2(new_n211), .A3(new_n205), .A4(new_n209), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n210), .A2(KEYINPUT69), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n241), .A2(new_n242), .A3(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n229), .A2(new_n240), .A3(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(KEYINPUT27), .B(G183gat), .Z(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT72), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT28), .B1(new_n250), .B2(G190gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT71), .ZN(new_n252));
  OR3_X1    g051(.A1(new_n252), .A2(new_n203), .A3(KEYINPUT27), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT27), .B1(new_n252), .B2(new_n203), .ZN(new_n254));
  NOR2_X1   g053(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT26), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n219), .A2(new_n257), .A3(new_n216), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n223), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n251), .A2(new_n256), .A3(new_n258), .A4(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n248), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT29), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G226gat), .A2(G233gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G197gat), .B(G204gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(G211gat), .A2(G218gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT22), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n267), .A2(KEYINPUT75), .A3(new_n268), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n267), .ZN(new_n271));
  NOR2_X1   g070(.A1(G211gat), .A2(G218gat), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT76), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n272), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT76), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(new_n275), .A3(new_n267), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT75), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n277), .B1(new_n271), .B2(KEYINPUT22), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n270), .A2(new_n273), .A3(new_n276), .A4(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n269), .A3(new_n266), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(new_n273), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT77), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n279), .A2(new_n282), .A3(KEYINPUT77), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n264), .B(KEYINPUT78), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n261), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n265), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n279), .A2(KEYINPUT77), .A3(new_n282), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT77), .B1(new_n279), .B2(new_n282), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n288), .B1(new_n261), .B2(new_n262), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n264), .B1(new_n248), .B2(new_n260), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G8gat), .B(G36gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(KEYINPUT79), .ZN(new_n298));
  XNOR2_X1  g097(.A(G64gat), .B(G92gat), .ZN(new_n299));
  XOR2_X1   g098(.A(new_n298), .B(new_n299), .Z(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n290), .A2(new_n296), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT80), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT30), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT80), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n290), .A2(new_n296), .A3(new_n305), .A4(new_n301), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n303), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n301), .B1(new_n290), .B2(new_n296), .ZN(new_n308));
  AND3_X1   g107(.A1(new_n290), .A2(new_n296), .A3(new_n301), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n308), .B1(new_n309), .B2(KEYINPUT30), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT5), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT84), .ZN(new_n313));
  XNOR2_X1  g112(.A(G141gat), .B(G148gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT83), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT2), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n316), .A2(new_n317), .B1(G155gat), .B2(G162gat), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n314), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT82), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n323));
  AND3_X1   g122(.A1(KEYINPUT81), .A2(G155gat), .A3(G162gat), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT81), .B1(G155gat), .B2(G162gat), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n322), .B(new_n323), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n313), .B1(new_n319), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n314), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n316), .A2(new_n317), .ZN(new_n329));
  NAND2_X1  g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(new_n315), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  OR2_X1    g131(.A1(new_n324), .A2(new_n325), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n322), .A2(new_n323), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .A4(KEYINPUT84), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n327), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n317), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n314), .B1(new_n330), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G127gat), .B(G134gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G113gat), .B(G120gat), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n342), .B1(KEYINPUT1), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n343), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT1), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(new_n341), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT85), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n344), .A2(new_n347), .A3(KEYINPUT85), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n340), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n338), .B1(new_n327), .B2(new_n335), .ZN(new_n354));
  INV_X1    g153(.A(new_n348), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G225gat), .A2(G233gat), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n312), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT4), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n352), .B1(new_n354), .B2(new_n363), .ZN(new_n364));
  AOI211_X1 g163(.A(KEYINPUT3), .B(new_n338), .C1(new_n327), .C2(new_n335), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n362), .B(new_n358), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT86), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n354), .A2(new_n367), .ZN(new_n368));
  AOI211_X1 g167(.A(KEYINPUT86), .B(new_n338), .C1(new_n327), .C2(new_n335), .ZN(new_n369));
  NOR4_X1   g168(.A1(new_n368), .A2(new_n369), .A3(new_n361), .A4(new_n348), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n360), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n312), .B(new_n358), .C1(new_n364), .C2(new_n365), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n340), .A2(KEYINPUT86), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n354), .A2(new_n367), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n374), .A2(new_n361), .A3(new_n355), .A4(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n356), .A2(KEYINPUT4), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n371), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G1gat), .B(G29gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT0), .ZN(new_n382));
  XNOR2_X1  g181(.A(G57gat), .B(G85gat), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n382), .B(new_n383), .Z(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n379), .A3(new_n384), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AOI211_X1 g188(.A(new_n387), .B(new_n384), .C1(new_n371), .C2(new_n379), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n311), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G78gat), .B(G106gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT31), .B(G50gat), .ZN(new_n395));
  XOR2_X1   g194(.A(new_n394), .B(new_n395), .Z(new_n396));
  XOR2_X1   g195(.A(KEYINPUT88), .B(G22gat), .Z(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT29), .B1(new_n354), .B2(new_n363), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n399), .A2(new_n287), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT29), .B1(new_n279), .B2(new_n282), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n401), .A2(KEYINPUT3), .ZN(new_n402));
  OAI211_X1 g201(.A(G228gat), .B(G233gat), .C1(new_n402), .C2(new_n354), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT87), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n405), .B1(new_n399), .B2(new_n287), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n293), .B(KEYINPUT87), .C1(new_n365), .C2(KEYINPUT29), .ZN(new_n407));
  OAI22_X1  g206(.A1(new_n368), .A2(new_n369), .B1(KEYINPUT3), .B2(new_n401), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(G228gat), .A2(G233gat), .ZN(new_n410));
  AOI211_X1 g209(.A(new_n398), .B(new_n404), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n410), .ZN(new_n412));
  INV_X1    g211(.A(new_n404), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n397), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n396), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT89), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT89), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n417), .B(new_n396), .C1(new_n411), .C2(new_n414), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n404), .B1(new_n409), .B2(new_n410), .ZN(new_n420));
  INV_X1    g219(.A(G22gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n422), .A2(new_n411), .A3(new_n396), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n355), .B1(new_n248), .B2(new_n260), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n248), .A2(new_n355), .A3(new_n260), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G227gat), .A2(G233gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT34), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT34), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n427), .A2(new_n433), .A3(new_n430), .A4(new_n428), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT73), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n248), .A2(new_n355), .A3(new_n260), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n431), .B1(new_n437), .B2(new_n426), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT32), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  XOR2_X1   g240(.A(G15gat), .B(G43gat), .Z(new_n442));
  XNOR2_X1  g241(.A(G71gat), .B(G99gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n439), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n444), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n438), .B(KEYINPUT32), .C1(new_n440), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n436), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n436), .A2(new_n448), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n393), .A2(new_n425), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT35), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT90), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n311), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n307), .A2(new_n310), .A3(KEYINPUT90), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n423), .B1(new_n416), .B2(new_n418), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n389), .A2(new_n391), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT35), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n448), .A2(KEYINPUT74), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT74), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n445), .A2(new_n464), .A3(new_n447), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n435), .A3(new_n465), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n448), .A2(KEYINPUT74), .A3(new_n432), .A4(new_n434), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n457), .A2(new_n462), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n378), .B1(new_n365), .B2(new_n364), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n359), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT39), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n357), .A2(new_n359), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT91), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n472), .B(new_n476), .C1(new_n475), .C2(new_n474), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n471), .A2(new_n473), .A3(new_n359), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n384), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT40), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n479), .A2(new_n480), .B1(new_n385), .B2(new_n380), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n455), .A2(new_n456), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n263), .A2(new_n264), .B1(new_n288), .B2(new_n261), .ZN(new_n484));
  OR3_X1    g283(.A1(new_n484), .A2(KEYINPUT92), .A3(new_n287), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT92), .B1(new_n484), .B2(new_n287), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n294), .A2(new_n295), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n485), .B(new_n486), .C1(new_n487), .C2(new_n293), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT37), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT37), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n290), .A2(new_n296), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n300), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n492), .A2(KEYINPUT38), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n389), .A2(new_n391), .A3(new_n303), .A4(new_n306), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n490), .B1(new_n290), .B2(new_n296), .ZN(new_n497));
  OAI211_X1 g296(.A(KEYINPUT93), .B(KEYINPUT38), .C1(new_n492), .C2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n290), .A2(new_n296), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT37), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n501), .A2(new_n300), .A3(new_n491), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT93), .B1(new_n502), .B2(KEYINPUT38), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n494), .B(new_n496), .C1(new_n499), .C2(new_n503), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n483), .A2(new_n504), .A3(new_n425), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n465), .A2(new_n435), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n464), .B1(new_n445), .B2(new_n447), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n467), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n419), .B(new_n424), .C1(new_n311), .C2(new_n392), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n449), .A2(KEYINPUT36), .A3(new_n450), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n470), .B1(new_n505), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT15), .ZN(new_n516));
  INV_X1    g315(.A(G43gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n517), .A2(G50gat), .ZN(new_n518));
  INV_X1    g317(.A(G50gat), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(G43gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n516), .B1(new_n521), .B2(KEYINPUT95), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT95), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n523), .B1(new_n518), .B2(new_n520), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT96), .B(G29gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(G36gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(G29gat), .A2(G36gat), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n528), .A2(KEYINPUT14), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(KEYINPUT14), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT97), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n519), .A2(G43gat), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n520), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n518), .A2(KEYINPUT97), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT15), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n525), .B1(new_n531), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n531), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n538), .A2(new_n524), .A3(new_n522), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT17), .ZN(new_n541));
  XNOR2_X1  g340(.A(G15gat), .B(G22gat), .ZN(new_n542));
  INV_X1    g341(.A(G1gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT16), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(G1gat), .B2(new_n542), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n546), .B(G8gat), .Z(new_n547));
  INV_X1    g346(.A(KEYINPUT17), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n537), .A2(new_n539), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n541), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G229gat), .A2(G233gat), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n547), .A2(new_n540), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT18), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n550), .A2(KEYINPUT18), .A3(new_n552), .A4(new_n551), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n551), .B(KEYINPUT13), .Z(new_n557));
  AND2_X1   g356(.A1(new_n547), .A2(new_n540), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n547), .A2(new_n540), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n555), .A2(new_n556), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G113gat), .B(G141gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT94), .B(G197gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT11), .B(G169gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT12), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n561), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n555), .A2(new_n556), .A3(new_n560), .A4(new_n567), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G71gat), .B(G78gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT98), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n575), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G57gat), .B(G64gat), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n573), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(G57gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(G64gat), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n572), .B1(KEYINPUT99), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n583), .B1(KEYINPUT99), .B2(new_n579), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT100), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n576), .A2(new_n585), .A3(new_n577), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n574), .A2(new_n575), .ZN(new_n587));
  NAND2_X1  g386(.A1(G71gat), .A2(G78gat), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT9), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n588), .A2(new_n575), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT100), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n584), .A2(new_n592), .A3(KEYINPUT101), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT101), .B1(new_n584), .B2(new_n592), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n580), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT21), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(KEYINPUT103), .B(KEYINPUT19), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G183gat), .B(G211gat), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n599), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n547), .B1(new_n595), .B2(new_n596), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n605), .A2(KEYINPUT104), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(KEYINPUT104), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G127gat), .B(G155gat), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT20), .ZN(new_n610));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n611), .B(KEYINPUT102), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n610), .B(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n608), .A2(new_n613), .ZN(new_n615));
  OR3_X1    g414(.A1(new_n604), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n604), .B1(new_n614), .B2(new_n615), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(KEYINPUT106), .B(G85gat), .Z(new_n619));
  INV_X1    g418(.A(G92gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(G99gat), .A2(G106gat), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n619), .A2(new_n620), .B1(KEYINPUT8), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G99gat), .B(G106gat), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT105), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(G85gat), .A3(G92gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT7), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n622), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n623), .B1(new_n622), .B2(new_n626), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n630), .A2(new_n540), .ZN(new_n631));
  AND2_X1   g430(.A1(G232gat), .A2(G233gat), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n631), .B1(KEYINPUT41), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n541), .A2(new_n549), .A3(new_n630), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G190gat), .B(G218gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT107), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n635), .B(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n632), .A2(KEYINPUT41), .ZN(new_n640));
  XNOR2_X1  g439(.A(G134gat), .B(G162gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n639), .A2(new_n642), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n595), .A2(new_n630), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT10), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n629), .B(new_n580), .C1(new_n593), .C2(new_n594), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n650), .A2(new_n649), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n647), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n646), .B1(new_n648), .B2(new_n650), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(G120gat), .B(G148gat), .Z(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT108), .ZN(new_n657));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n657), .B(new_n658), .Z(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n653), .A2(new_n654), .A3(new_n659), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n618), .A2(new_n645), .A3(new_n664), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n515), .A2(new_n571), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n392), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G1gat), .ZN(G1324gat));
  INV_X1    g467(.A(new_n666), .ZN(new_n669));
  OAI21_X1  g468(.A(G8gat), .B1(new_n669), .B2(new_n457), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT42), .ZN(new_n671));
  INV_X1    g470(.A(new_n457), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT16), .B(G8gat), .Z(new_n673));
  NAND3_X1  g472(.A1(new_n666), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  AND3_X1   g473(.A1(new_n674), .A2(KEYINPUT109), .A3(new_n671), .ZN(new_n675));
  AOI21_X1  g474(.A(KEYINPUT109), .B1(new_n674), .B2(new_n671), .ZN(new_n676));
  OAI221_X1 g475(.A(new_n670), .B1(new_n671), .B2(new_n674), .C1(new_n675), .C2(new_n676), .ZN(G1325gat));
  NAND2_X1  g476(.A1(new_n511), .A2(new_n513), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(G15gat), .B1(new_n669), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n468), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n681), .A2(G15gat), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n680), .B1(new_n669), .B2(new_n682), .ZN(G1326gat));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n458), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT43), .B(G22gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  NAND2_X1  g485(.A1(new_n502), .A2(KEYINPUT38), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT93), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n498), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n495), .B1(new_n489), .B2(new_n493), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n458), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n483), .ZN(new_n693));
  INV_X1    g492(.A(new_n514), .ZN(new_n694));
  AOI22_X1  g493(.A1(new_n693), .A2(new_n694), .B1(new_n453), .B2(new_n469), .ZN(new_n695));
  INV_X1    g494(.A(new_n571), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n618), .ZN(new_n698));
  INV_X1    g497(.A(new_n645), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n698), .A2(new_n699), .A3(new_n664), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n459), .A2(new_n526), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n697), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT45), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(new_n695), .B2(new_n699), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n515), .A2(KEYINPUT44), .A3(new_n645), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n569), .A2(KEYINPUT110), .A3(new_n570), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT110), .B1(new_n569), .B2(new_n570), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n698), .A2(new_n664), .A3(new_n710), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n705), .A2(new_n706), .A3(new_n392), .A4(new_n711), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n712), .A2(KEYINPUT111), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n526), .B1(new_n712), .B2(KEYINPUT111), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n703), .B1(new_n713), .B2(new_n714), .ZN(G1328gat));
  INV_X1    g514(.A(G36gat), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n697), .A2(new_n716), .A3(new_n672), .A4(new_n700), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT46), .Z(new_n718));
  AND4_X1   g517(.A1(new_n672), .A2(new_n705), .A3(new_n706), .A4(new_n711), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n716), .B2(new_n719), .ZN(G1329gat));
  NOR2_X1   g519(.A1(new_n679), .A2(new_n517), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n705), .A2(new_n706), .A3(new_n711), .A4(new_n721), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n697), .A2(new_n468), .A3(new_n700), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n723), .B2(G43gat), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g524(.A(KEYINPUT48), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(KEYINPUT112), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n697), .A2(new_n458), .A3(new_n700), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n727), .B1(new_n728), .B2(new_n519), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(KEYINPUT112), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n425), .A2(new_n519), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n705), .A2(new_n706), .A3(new_n711), .A4(new_n731), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n730), .B1(new_n729), .B2(new_n732), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(G1331gat));
  NOR4_X1   g534(.A1(new_n618), .A2(new_n645), .A3(new_n663), .A4(new_n709), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n515), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(new_n459), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(new_n581), .ZN(G1332gat));
  INV_X1    g538(.A(KEYINPUT113), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n515), .A2(KEYINPUT113), .A3(new_n736), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n457), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT114), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT114), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n741), .A2(new_n746), .A3(new_n742), .A4(new_n743), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT49), .ZN(new_n749));
  INV_X1    g548(.A(G64gat), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n745), .A2(new_n749), .A3(new_n750), .A4(new_n747), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(G1333gat));
  NAND4_X1  g553(.A1(new_n741), .A2(G71gat), .A3(new_n678), .A4(new_n742), .ZN(new_n755));
  INV_X1    g554(.A(G71gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n737), .B2(new_n681), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT50), .ZN(G1334gat));
  NAND3_X1  g558(.A1(new_n741), .A2(new_n458), .A3(new_n742), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G78gat), .ZN(G1335gat));
  OAI21_X1  g560(.A(KEYINPUT115), .B1(new_n698), .B2(new_n709), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT115), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n618), .A2(new_n763), .A3(new_n710), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n514), .B1(new_n483), .B2(new_n692), .ZN(new_n766));
  INV_X1    g565(.A(new_n461), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n468), .A2(new_n425), .A3(new_n767), .ZN(new_n768));
  AOI22_X1  g567(.A1(new_n768), .A2(new_n457), .B1(new_n452), .B2(KEYINPUT35), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n645), .B(new_n765), .C1(new_n766), .C2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n515), .A2(KEYINPUT51), .A3(new_n645), .A4(new_n765), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n392), .A2(new_n619), .A3(new_n664), .ZN(new_n777));
  INV_X1    g576(.A(new_n765), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(new_n663), .ZN(new_n779));
  AND4_X1   g578(.A1(new_n392), .A2(new_n705), .A3(new_n706), .A4(new_n779), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n776), .A2(new_n777), .B1(new_n780), .B2(new_n619), .ZN(G1336gat));
  NAND3_X1  g580(.A1(new_n772), .A2(KEYINPUT116), .A3(new_n774), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n770), .A2(new_n783), .A3(new_n771), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n457), .A2(G92gat), .A3(new_n663), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n782), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n705), .A2(new_n706), .A3(new_n672), .A4(new_n779), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G92gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT52), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n785), .B1(new_n773), .B2(new_n775), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n791), .A2(new_n788), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n790), .A2(new_n793), .ZN(G1337gat));
  NAND4_X1  g593(.A1(new_n705), .A2(new_n706), .A3(new_n678), .A4(new_n779), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT117), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(G99gat), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n795), .A2(new_n796), .ZN(new_n799));
  OR3_X1    g598(.A1(new_n681), .A2(G99gat), .A3(new_n663), .ZN(new_n800));
  OAI22_X1  g599(.A1(new_n798), .A2(new_n799), .B1(new_n776), .B2(new_n800), .ZN(G1338gat));
  NOR3_X1   g600(.A1(new_n425), .A2(G106gat), .A3(new_n663), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n782), .A2(new_n784), .A3(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n705), .A2(new_n706), .A3(new_n458), .A4(new_n779), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(G106gat), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT53), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n802), .B1(new_n773), .B2(new_n775), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n805), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n807), .A2(new_n810), .ZN(G1339gat));
  NAND2_X1  g610(.A1(new_n457), .A2(new_n392), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n653), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n651), .A2(new_n652), .A3(new_n815), .A4(new_n647), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n651), .A2(new_n652), .A3(new_n647), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT118), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n814), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n660), .B1(new_n653), .B2(new_n813), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n662), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI211_X1 g622(.A(new_n822), .B(new_n660), .C1(new_n653), .C2(new_n813), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT119), .B1(new_n819), .B2(new_n824), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n819), .A2(new_n824), .A3(KEYINPUT119), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n709), .B(new_n823), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n551), .B1(new_n550), .B2(new_n552), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n558), .A2(new_n559), .A3(new_n557), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n566), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n570), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n664), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n645), .B1(new_n827), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n645), .A2(new_n832), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n618), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n698), .A2(new_n699), .A3(new_n663), .A4(new_n710), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n812), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n458), .B1(new_n449), .B2(new_n450), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(G113gat), .B1(new_n842), .B2(new_n709), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n458), .B1(new_n838), .B2(new_n839), .ZN(new_n844));
  AND4_X1   g643(.A1(new_n392), .A2(new_n844), .A3(new_n457), .A4(new_n468), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n571), .A2(G113gat), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n843), .B1(new_n845), .B2(new_n846), .ZN(G1340gat));
  AOI21_X1  g646(.A(G120gat), .B1(new_n842), .B2(new_n664), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n664), .A2(G120gat), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n845), .B2(new_n849), .ZN(G1341gat));
  AND3_X1   g649(.A1(new_n845), .A2(G127gat), .A3(new_n698), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n842), .A2(new_n698), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(KEYINPUT120), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n853), .A2(G127gat), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(KEYINPUT120), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n851), .B1(new_n854), .B2(new_n855), .ZN(G1342gat));
  INV_X1    g655(.A(KEYINPUT56), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n699), .A2(G134gat), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n842), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n859), .B(KEYINPUT121), .Z(new_n860));
  AOI21_X1  g659(.A(new_n857), .B1(new_n842), .B2(new_n858), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n645), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n862), .B2(G134gat), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n860), .A2(new_n863), .ZN(G1343gat));
  NOR2_X1   g663(.A1(new_n812), .A2(new_n678), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n838), .A2(new_n839), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT57), .B1(new_n866), .B2(new_n458), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n458), .A2(KEYINPUT57), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n823), .B(new_n571), .C1(new_n825), .C2(new_n826), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n645), .B1(new_n869), .B2(new_n833), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n618), .B1(new_n870), .B2(new_n837), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n868), .B1(new_n871), .B2(new_n839), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n865), .B1(new_n867), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G141gat), .B1(new_n873), .B2(new_n696), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n678), .A2(new_n425), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n840), .A2(new_n875), .ZN(new_n876));
  OR3_X1    g675(.A1(new_n876), .A2(G141gat), .A3(new_n696), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n874), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G141gat), .B1(new_n873), .B2(new_n710), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n880), .A2(new_n877), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n879), .B1(new_n881), .B2(new_n878), .ZN(G1344gat));
  NAND2_X1  g681(.A1(new_n665), .A2(new_n696), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n871), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n458), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n886));
  INV_X1    g685(.A(new_n868), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n885), .A2(new_n886), .B1(new_n866), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n865), .A2(new_n664), .ZN(new_n889));
  OAI21_X1  g688(.A(G148gat), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(KEYINPUT59), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n664), .B(new_n865), .C1(new_n867), .C2(new_n872), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893));
  INV_X1    g692(.A(G148gat), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(KEYINPUT59), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n893), .B1(new_n892), .B2(new_n895), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n891), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n840), .A2(new_n894), .A3(new_n664), .A4(new_n875), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1345gat));
  OAI21_X1  g699(.A(G155gat), .B1(new_n873), .B2(new_n618), .ZN(new_n901));
  OR3_X1    g700(.A1(new_n876), .A2(G155gat), .A3(new_n618), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT123), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1346gat));
  NAND2_X1  g706(.A1(new_n645), .A2(G162gat), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n876), .A2(new_n699), .ZN(new_n909));
  OAI22_X1  g708(.A1(new_n873), .A2(new_n908), .B1(new_n909), .B2(G162gat), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT124), .ZN(G1347gat));
  NAND2_X1  g710(.A1(new_n672), .A2(new_n459), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n912), .B1(new_n838), .B2(new_n839), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n913), .A2(new_n841), .ZN(new_n914));
  AOI21_X1  g713(.A(G169gat), .B1(new_n914), .B2(new_n709), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n912), .A2(new_n681), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n844), .A2(new_n916), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n917), .A2(new_n213), .A3(new_n696), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n915), .A2(new_n918), .ZN(G1348gat));
  NAND3_X1  g718(.A1(new_n914), .A2(new_n214), .A3(new_n664), .ZN(new_n920));
  OAI21_X1  g719(.A(G176gat), .B1(new_n917), .B2(new_n663), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1349gat));
  INV_X1    g721(.A(new_n250), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n914), .A2(new_n923), .A3(new_n698), .ZN(new_n924));
  OAI21_X1  g723(.A(G183gat), .B1(new_n917), .B2(new_n618), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g725(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n927));
  XOR2_X1   g726(.A(new_n926), .B(new_n927), .Z(G1350gat));
  NAND3_X1  g727(.A1(new_n914), .A2(new_n204), .A3(new_n645), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n930));
  INV_X1    g729(.A(new_n917), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n645), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n930), .B1(new_n932), .B2(G190gat), .ZN(new_n933));
  AOI211_X1 g732(.A(KEYINPUT61), .B(new_n204), .C1(new_n931), .C2(new_n645), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(G1351gat));
  NAND2_X1  g734(.A1(new_n913), .A2(new_n875), .ZN(new_n936));
  OR3_X1    g735(.A1(new_n936), .A2(G197gat), .A3(new_n710), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT126), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n866), .A2(new_n887), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n425), .B1(new_n871), .B2(new_n883), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(KEYINPUT57), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n912), .A2(new_n678), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n938), .B1(new_n943), .B2(new_n696), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(G197gat), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n943), .A2(new_n938), .A3(new_n696), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n937), .B1(new_n945), .B2(new_n946), .ZN(G1352gat));
  NOR3_X1   g746(.A1(new_n936), .A2(G204gat), .A3(new_n663), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT62), .ZN(new_n949));
  OAI21_X1  g748(.A(G204gat), .B1(new_n943), .B2(new_n663), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1353gat));
  OR3_X1    g750(.A1(new_n936), .A2(G211gat), .A3(new_n618), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n941), .A2(new_n698), .A3(new_n942), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n953), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n954));
  AOI21_X1  g753(.A(KEYINPUT63), .B1(new_n953), .B2(G211gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(G1354gat));
  INV_X1    g755(.A(new_n936), .ZN(new_n957));
  AOI21_X1  g756(.A(G218gat), .B1(new_n957), .B2(new_n645), .ZN(new_n958));
  INV_X1    g757(.A(new_n943), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n645), .A2(G218gat), .ZN(new_n960));
  XOR2_X1   g759(.A(new_n960), .B(KEYINPUT127), .Z(new_n961));
  AOI21_X1  g760(.A(new_n958), .B1(new_n959), .B2(new_n961), .ZN(G1355gat));
endmodule


