//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XOR2_X1   g002(.A(G197gat), .B(G204gat), .Z(new_n204));
  OR2_X1    g003(.A1(KEYINPUT72), .A2(G218gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(KEYINPUT72), .A2(G218gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G211gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT22), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(KEYINPUT73), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT73), .ZN(new_n211));
  INV_X1    g010(.A(G211gat), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n212), .B1(new_n205), .B2(new_n206), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n211), .B1(new_n213), .B2(KEYINPUT22), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n204), .B1(new_n210), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n203), .B1(new_n215), .B2(KEYINPUT74), .ZN(new_n216));
  INV_X1    g015(.A(new_n204), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT73), .B1(new_n208), .B2(new_n209), .ZN(new_n218));
  NOR3_X1   g017(.A1(new_n213), .A2(new_n211), .A3(KEYINPUT22), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT74), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(new_n221), .A3(new_n202), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n216), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G226gat), .A2(G233gat), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT27), .B(G183gat), .ZN(new_n227));
  INV_X1    g026(.A(G190gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n229), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT26), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(KEYINPUT26), .ZN(new_n233));
  NOR2_X1   g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236));
  INV_X1    g035(.A(G169gat), .ZN(new_n237));
  INV_X1    g036(.A(G176gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(new_n231), .A3(KEYINPUT26), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n235), .A2(new_n236), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G183gat), .ZN(new_n242));
  OR3_X1    g041(.A1(new_n242), .A2(KEYINPUT66), .A3(KEYINPUT27), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT27), .B1(new_n242), .B2(KEYINPUT66), .ZN(new_n244));
  NOR2_X1   g043(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n241), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT23), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n248), .A2(G169gat), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT64), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n238), .ZN(new_n251));
  NAND2_X1  g050(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n236), .A2(KEYINPUT23), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(new_n239), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT65), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT24), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n257), .A2(G183gat), .A3(G190gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(G183gat), .B(G190gat), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n258), .B1(new_n259), .B2(new_n257), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n253), .A2(new_n255), .A3(KEYINPUT65), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT25), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n255), .B(KEYINPUT25), .C1(new_n248), .C2(new_n239), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(new_n260), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n247), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT29), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n226), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n265), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n253), .A2(KEYINPUT65), .A3(new_n255), .ZN(new_n270));
  NOR3_X1   g069(.A1(new_n270), .A2(new_n256), .A3(new_n260), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n269), .B1(new_n271), .B2(KEYINPUT25), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n225), .B1(new_n272), .B2(new_n247), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n224), .B1(new_n268), .B2(new_n273), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n230), .A2(new_n241), .A3(new_n246), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT65), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n237), .A2(KEYINPUT23), .ZN(new_n277));
  AND2_X1   g076(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n234), .B1(KEYINPUT23), .B2(new_n236), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n276), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n260), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(new_n283), .A3(new_n262), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT25), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n275), .B1(new_n286), .B2(new_n269), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n225), .B1(new_n287), .B2(KEYINPUT29), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n266), .A2(new_n226), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(new_n223), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n292));
  XNOR2_X1  g091(.A(G8gat), .B(G36gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(G64gat), .B(G92gat), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n293), .B(new_n294), .Z(new_n295));
  NAND4_X1  g094(.A1(new_n291), .A2(new_n292), .A3(KEYINPUT30), .A4(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT30), .ZN(new_n297));
  INV_X1    g096(.A(new_n295), .ZN(new_n298));
  AOI211_X1 g097(.A(new_n297), .B(new_n298), .C1(new_n274), .C2(new_n290), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n274), .A2(new_n298), .A3(new_n290), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT75), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n296), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NOR3_X1   g101(.A1(new_n268), .A2(new_n224), .A3(new_n273), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n223), .B1(new_n288), .B2(new_n289), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n295), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT76), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n307), .A3(new_n295), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n297), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n302), .A2(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT2), .ZN(new_n312));
  NOR2_X1   g111(.A1(G155gat), .A2(G162gat), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G141gat), .ZN(new_n315));
  INV_X1    g114(.A(G148gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G141gat), .A2(G148gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT78), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(G141gat), .A2(G148gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT78), .ZN(new_n324));
  NOR3_X1   g123(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n323), .B(new_n324), .C1(new_n311), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT77), .B1(new_n321), .B2(new_n322), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT77), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n317), .A2(new_n329), .A3(new_n318), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n330), .A3(new_n312), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n311), .A2(new_n313), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT3), .ZN(new_n335));
  INV_X1    g134(.A(G134gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G127gat), .ZN(new_n337));
  INV_X1    g136(.A(G127gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G134gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G120gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G113gat), .ZN(new_n343));
  INV_X1    g142(.A(G113gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G120gat), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT1), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT68), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n347), .B1(G127gat), .B2(new_n336), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n341), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n337), .A2(KEYINPUT68), .ZN(new_n350));
  XNOR2_X1  g149(.A(G113gat), .B(G120gat), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n340), .B(new_n350), .C1(new_n351), .C2(KEYINPUT1), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n349), .A2(KEYINPUT79), .A3(new_n352), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n320), .A2(new_n326), .B1(new_n331), .B2(new_n332), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT3), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n349), .A2(new_n352), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n335), .A2(new_n353), .A3(new_n356), .A4(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT69), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n349), .A2(KEYINPUT69), .A3(new_n352), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(new_n354), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n354), .A2(KEYINPUT4), .A3(new_n349), .A4(new_n352), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n360), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n359), .A2(new_n334), .A3(new_n353), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT80), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n354), .A2(new_n349), .A3(new_n352), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n359), .A2(new_n334), .A3(KEYINPUT80), .A4(new_n353), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n374), .A2(new_n369), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n371), .A2(KEYINPUT39), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT83), .B(KEYINPUT39), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n368), .A2(new_n370), .A3(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G1gat), .B(G29gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT0), .ZN(new_n383));
  XNOR2_X1  g182(.A(G57gat), .B(G85gat), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n383), .B(new_n384), .Z(new_n385));
  NAND2_X1  g184(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT84), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n381), .A2(KEYINPUT84), .A3(new_n385), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n379), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n366), .A2(new_n367), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT5), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n391), .A2(new_n392), .A3(new_n369), .A4(new_n360), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n394), .A2(new_n370), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n360), .A2(new_n369), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n375), .A2(new_n365), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(new_n365), .B2(new_n364), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT5), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n393), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n385), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n390), .A2(KEYINPUT40), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT85), .B1(new_n390), .B2(KEYINPUT40), .ZN(new_n403));
  INV_X1    g202(.A(new_n389), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT84), .B1(new_n381), .B2(new_n385), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n378), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT85), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT40), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n310), .A2(new_n402), .A3(new_n403), .A4(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G78gat), .B(G106gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT31), .B(G50gat), .ZN(new_n412));
  XOR2_X1   g211(.A(new_n411), .B(new_n412), .Z(new_n413));
  INV_X1    g212(.A(KEYINPUT82), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n267), .B1(new_n215), .B2(new_n203), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n220), .A2(new_n202), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n355), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n334), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n356), .A2(new_n267), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n223), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G228gat), .A2(G233gat), .ZN(new_n423));
  XOR2_X1   g222(.A(new_n423), .B(KEYINPUT81), .Z(new_n424));
  AOI21_X1  g223(.A(new_n415), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n421), .A2(G228gat), .A3(G233gat), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n216), .A2(new_n222), .A3(new_n267), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n354), .B1(new_n427), .B2(new_n355), .ZN(new_n428));
  OR2_X1    g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(G22gat), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n425), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n418), .A2(new_n334), .B1(new_n223), .B2(new_n420), .ZN(new_n434));
  INV_X1    g233(.A(new_n424), .ZN(new_n435));
  OAI22_X1  g234(.A1(new_n434), .A2(new_n435), .B1(new_n414), .B2(new_n413), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n426), .A2(new_n428), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n431), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n385), .A2(KEYINPUT6), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT6), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n401), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n400), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n394), .A2(new_n370), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n445), .B(KEYINPUT5), .C1(new_n396), .C2(new_n398), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n446), .A2(new_n442), .A3(new_n393), .A4(new_n401), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n306), .A2(new_n308), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n291), .A2(KEYINPUT37), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT37), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n274), .A2(new_n452), .A3(new_n290), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n298), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT38), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT38), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n454), .A2(new_n457), .A3(new_n298), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n450), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n410), .A2(new_n440), .A3(new_n459), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n349), .A2(KEYINPUT69), .A3(new_n352), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT69), .B1(new_n349), .B2(new_n352), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n272), .A2(new_n463), .A3(new_n247), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n362), .A2(new_n363), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n265), .B1(new_n284), .B2(new_n285), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n465), .B1(new_n466), .B2(new_n275), .ZN(new_n467));
  NAND2_X1  g266(.A1(G227gat), .A2(G233gat), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n464), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n469), .B(KEYINPUT34), .ZN(new_n470));
  XNOR2_X1  g269(.A(G15gat), .B(G43gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(KEYINPUT70), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(G71gat), .ZN(new_n473));
  OR2_X1    g272(.A1(new_n471), .A2(KEYINPUT70), .ZN(new_n474));
  INV_X1    g273(.A(G71gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n471), .A2(KEYINPUT70), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(G99gat), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n468), .B1(new_n464), .B2(new_n467), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(KEYINPUT33), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT32), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n464), .A2(new_n467), .ZN(new_n485));
  INV_X1    g284(.A(new_n468), .ZN(new_n486));
  AOI221_X4 g285(.A(new_n482), .B1(new_n479), .B2(KEYINPUT33), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n484), .A2(new_n487), .A3(KEYINPUT71), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT71), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n465), .A2(new_n466), .A3(new_n275), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n463), .B1(new_n272), .B2(new_n247), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n486), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT32), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT33), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n495), .A3(new_n479), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n483), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n489), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n470), .B1(new_n488), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT34), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n469), .B(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n496), .A2(new_n501), .A3(new_n497), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT36), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n484), .A2(new_n470), .A3(new_n487), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n501), .B1(new_n496), .B2(new_n497), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n302), .A2(new_n309), .A3(new_n448), .ZN(new_n510));
  AOI22_X1  g309(.A1(new_n505), .A2(new_n509), .B1(new_n439), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n439), .A2(new_n507), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n499), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT35), .B1(new_n513), .B2(new_n510), .ZN(new_n514));
  NOR4_X1   g313(.A1(new_n439), .A2(new_n507), .A3(new_n508), .A4(KEYINPUT35), .ZN(new_n515));
  INV_X1    g314(.A(new_n510), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n460), .A2(new_n511), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G43gat), .B(G50gat), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(KEYINPUT15), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(KEYINPUT15), .ZN(new_n521));
  INV_X1    g320(.A(G29gat), .ZN(new_n522));
  INV_X1    g321(.A(G36gat), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT86), .ZN(new_n526));
  NOR3_X1   g325(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  AOI211_X1 g327(.A(new_n520), .B(new_n524), .C1(new_n526), .C2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT87), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n527), .B(new_n530), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n531), .A2(new_n526), .B1(G29gat), .B2(G36gat), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n532), .A2(new_n521), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT17), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT92), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT92), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(new_n537), .A3(KEYINPUT17), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT17), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(new_n529), .B2(new_n533), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT88), .ZN(new_n542));
  INV_X1    g341(.A(G8gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(G15gat), .B(G22gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT16), .ZN(new_n545));
  AOI21_X1  g344(.A(G1gat), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(KEYINPUT89), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n544), .B(KEYINPUT89), .C1(new_n545), .C2(G1gat), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n543), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT90), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n548), .A2(new_n543), .A3(new_n549), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT91), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n542), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G229gat), .A2(G233gat), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n555), .B1(new_n533), .B2(new_n529), .ZN(new_n559));
  NOR2_X1   g358(.A1(KEYINPUT93), .A2(KEYINPUT18), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n557), .A2(new_n558), .A3(new_n559), .A4(new_n561), .ZN(new_n562));
  OR3_X1    g361(.A1(new_n556), .A2(KEYINPUT94), .A3(new_n534), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n558), .B(KEYINPUT13), .Z(new_n564));
  NAND3_X1  g363(.A1(new_n552), .A2(new_n534), .A3(new_n554), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n559), .A2(KEYINPUT94), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G113gat), .B(G141gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G197gat), .ZN(new_n571));
  XOR2_X1   g370(.A(KEYINPUT11), .B(G169gat), .Z(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n573), .B(KEYINPUT12), .Z(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n560), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n569), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n576), .A2(new_n560), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n574), .B1(new_n579), .B2(new_n568), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n518), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G57gat), .B(G64gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT9), .ZN(new_n585));
  NAND2_X1  g384(.A1(G71gat), .A2(G78gat), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n586), .ZN(new_n588));
  NOR2_X1   g387(.A1(G71gat), .A2(G78gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n586), .A2(KEYINPUT95), .ZN(new_n591));
  OR3_X1    g390(.A1(new_n587), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n590), .B1(new_n587), .B2(new_n591), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n555), .B1(KEYINPUT21), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT96), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n594), .A2(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(G127gat), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n596), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G183gat), .B(G211gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT97), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n606));
  INV_X1    g405(.A(G155gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n605), .B(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n603), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n601), .A2(new_n602), .A3(new_n609), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(G99gat), .B(G106gat), .Z(new_n614));
  INV_X1    g413(.A(KEYINPUT99), .ZN(new_n615));
  INV_X1    g414(.A(G85gat), .ZN(new_n616));
  INV_X1    g415(.A(G92gat), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT7), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT7), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n619), .A2(G85gat), .A3(G92gat), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n614), .A2(new_n615), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(G99gat), .ZN(new_n622));
  INV_X1    g421(.A(G106gat), .ZN(new_n623));
  OAI21_X1  g422(.A(KEYINPUT8), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT98), .B(G85gat), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n621), .B(new_n624), .C1(G92gat), .C2(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n614), .A2(new_n615), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n539), .A2(new_n542), .A3(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(G232gat), .A2(G233gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(KEYINPUT41), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n634), .B1(new_n631), .B2(new_n534), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(G190gat), .B(G218gat), .Z(new_n638));
  AND2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n633), .A2(KEYINPUT41), .ZN(new_n641));
  XNOR2_X1  g440(.A(G134gat), .B(G162gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  OR3_X1    g443(.A1(new_n639), .A2(new_n640), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n644), .B1(new_n639), .B2(new_n640), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n613), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G230gat), .A2(G233gat), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n630), .A2(new_n594), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT10), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n628), .A2(new_n593), .A3(new_n592), .A4(new_n629), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n630), .A2(KEYINPUT10), .A3(new_n594), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n651), .A2(new_n653), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n656), .B1(new_n657), .B2(new_n650), .ZN(new_n658));
  XNOR2_X1  g457(.A(G120gat), .B(G148gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(G176gat), .B(G204gat), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n659), .B(new_n660), .Z(new_n661));
  OR2_X1    g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n656), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n657), .A2(new_n650), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(new_n664), .A3(new_n661), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n648), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n583), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n448), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT100), .B(G1gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1324gat));
  AND2_X1   g471(.A1(new_n668), .A2(new_n310), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT16), .B(G8gat), .Z(new_n674));
  AND2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n673), .A2(new_n543), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT42), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(KEYINPUT42), .B2(new_n675), .ZN(G1325gat));
  INV_X1    g477(.A(G15gat), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n507), .A2(new_n508), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n668), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT71), .B1(new_n484), .B2(new_n487), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n496), .A2(new_n489), .A3(new_n497), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n501), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n509), .B1(new_n684), .B2(new_n503), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n668), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n681), .B1(new_n687), .B2(new_n679), .ZN(G1326gat));
  NAND2_X1  g487(.A1(new_n668), .A2(new_n439), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT43), .B(G22gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1327gat));
  XNOR2_X1  g490(.A(new_n613), .B(KEYINPUT102), .ZN(new_n692));
  INV_X1    g491(.A(new_n666), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n575), .B1(new_n569), .B2(new_n577), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n579), .A2(new_n568), .A3(new_n574), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n578), .A2(new_n580), .A3(KEYINPUT101), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n692), .A2(new_n693), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT103), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(new_n518), .B2(new_n647), .ZN(new_n704));
  INV_X1    g503(.A(new_n647), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n510), .A2(new_n439), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n685), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n457), .B1(new_n454), .B2(new_n298), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n708), .A2(new_n448), .A3(new_n449), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n439), .B1(new_n709), .B2(new_n458), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n707), .B1(new_n710), .B2(new_n410), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n516), .A2(new_n499), .A3(new_n512), .ZN(new_n712));
  AOI22_X1  g511(.A1(new_n712), .A2(KEYINPUT35), .B1(new_n516), .B2(new_n515), .ZN(new_n713));
  OAI211_X1 g512(.A(KEYINPUT44), .B(new_n705), .C1(new_n711), .C2(new_n713), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n704), .A2(new_n714), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n702), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G29gat), .B1(new_n717), .B2(new_n448), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n613), .A2(new_n647), .A3(new_n666), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n583), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n721), .A2(new_n522), .A3(new_n669), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT45), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n718), .A2(new_n723), .ZN(G1328gat));
  INV_X1    g523(.A(new_n310), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n720), .A2(G36gat), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT46), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n716), .A2(new_n310), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT104), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G36gat), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n728), .A2(new_n729), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n727), .B1(new_n731), .B2(new_n732), .ZN(G1329gat));
  OAI21_X1  g532(.A(G43gat), .B1(new_n717), .B2(new_n685), .ZN(new_n734));
  INV_X1    g533(.A(new_n680), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n720), .A2(G43gat), .A3(new_n735), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n736), .B(KEYINPUT105), .Z(new_n737));
  NAND2_X1  g536(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT47), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1330gat));
  OAI21_X1  g539(.A(G50gat), .B1(new_n717), .B2(new_n440), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n721), .A2(KEYINPUT106), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n721), .A2(KEYINPUT106), .ZN(new_n743));
  OR4_X1    g542(.A1(G50gat), .A2(new_n742), .A3(new_n743), .A4(new_n440), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT48), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1331gat));
  NOR3_X1   g546(.A1(new_n700), .A2(new_n648), .A3(new_n693), .ZN(new_n748));
  XOR2_X1   g547(.A(new_n748), .B(KEYINPUT107), .Z(new_n749));
  NOR2_X1   g548(.A1(new_n749), .A2(new_n518), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n669), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G57gat), .ZN(G1332gat));
  INV_X1    g551(.A(KEYINPUT49), .ZN(new_n753));
  INV_X1    g552(.A(G64gat), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n750), .B(new_n310), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(G1333gat));
  AOI21_X1  g556(.A(new_n475), .B1(new_n750), .B2(new_n686), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n735), .A2(G71gat), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n758), .B1(new_n750), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g560(.A1(new_n750), .A2(new_n439), .ZN(new_n762));
  XOR2_X1   g561(.A(KEYINPUT108), .B(G78gat), .Z(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(G1335gat));
  INV_X1    g563(.A(new_n613), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n699), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n460), .A2(new_n511), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n514), .A2(new_n517), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n647), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n766), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT110), .B1(new_n518), .B2(new_n647), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n771), .A2(KEYINPUT51), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT51), .B1(new_n771), .B2(new_n772), .ZN(new_n774));
  OR2_X1    g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n693), .A2(new_n448), .A3(new_n625), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI211_X1 g576(.A(new_n693), .B(new_n613), .C1(new_n697), .C2(new_n698), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n704), .A2(new_n714), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT109), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n704), .A2(new_n714), .A3(KEYINPUT109), .A4(new_n778), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n625), .B1(new_n783), .B2(new_n448), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n777), .A2(new_n784), .ZN(G1336gat));
  NAND3_X1  g584(.A1(new_n666), .A2(new_n617), .A3(new_n310), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT111), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n775), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789));
  OAI21_X1  g588(.A(G92gat), .B1(new_n779), .B2(new_n725), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(G92gat), .B1(new_n783), .B2(new_n725), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n793), .B2(new_n789), .ZN(G1337gat));
  NAND4_X1  g593(.A1(new_n775), .A2(new_n622), .A3(new_n680), .A4(new_n666), .ZN(new_n795));
  OAI21_X1  g594(.A(G99gat), .B1(new_n783), .B2(new_n685), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(G1338gat));
  NOR3_X1   g596(.A1(new_n693), .A2(G106gat), .A3(new_n440), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n798), .B1(new_n773), .B2(new_n774), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n800));
  OAI21_X1  g599(.A(G106gat), .B1(new_n779), .B2(new_n440), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n781), .A2(new_n439), .A3(new_n782), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(G106gat), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n799), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n803), .B1(new_n806), .B2(KEYINPUT53), .ZN(new_n807));
  AOI211_X1 g606(.A(KEYINPUT112), .B(new_n800), .C1(new_n805), .C2(new_n799), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n802), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT113), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n811), .B(new_n802), .C1(new_n807), .C2(new_n808), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(G1339gat));
  NAND3_X1  g612(.A1(new_n654), .A2(new_n655), .A3(new_n650), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n663), .A2(KEYINPUT54), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n661), .B1(new_n656), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(KEYINPUT55), .A3(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(new_n665), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n815), .A2(new_n817), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n697), .A2(new_n824), .A3(new_n698), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n557), .A2(new_n559), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n564), .B1(new_n563), .B2(new_n566), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n828));
  OAI22_X1  g627(.A1(new_n826), .A2(new_n558), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n573), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT115), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n833), .B(new_n573), .C1(new_n829), .C2(new_n830), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n832), .A2(new_n578), .A3(new_n666), .A4(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n705), .B1(new_n825), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n832), .A2(new_n578), .A3(new_n834), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n837), .A2(new_n647), .A3(new_n823), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n692), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n667), .A2(new_n699), .ZN(new_n840));
  AOI211_X1 g639(.A(new_n439), .B(new_n735), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n310), .A2(new_n448), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n843), .A2(new_n344), .A3(new_n582), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n448), .B1(new_n839), .B2(new_n840), .ZN(new_n845));
  INV_X1    g644(.A(new_n513), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n845), .A2(new_n725), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(G113gat), .B1(new_n847), .B2(new_n700), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n844), .A2(new_n848), .ZN(G1340gat));
  OAI21_X1  g648(.A(G120gat), .B1(new_n843), .B2(new_n693), .ZN(new_n850));
  XOR2_X1   g649(.A(new_n850), .B(KEYINPUT116), .Z(new_n851));
  NAND3_X1  g650(.A1(new_n847), .A2(new_n342), .A3(new_n666), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(G1341gat));
  OAI21_X1  g652(.A(G127gat), .B1(new_n843), .B2(new_n692), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n847), .A2(new_n338), .A3(new_n613), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT117), .ZN(G1342gat));
  NAND3_X1  g656(.A1(new_n847), .A2(new_n336), .A3(new_n705), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n858), .A2(KEYINPUT56), .ZN(new_n859));
  OAI21_X1  g658(.A(G134gat), .B1(new_n843), .B2(new_n647), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(KEYINPUT56), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(G1343gat));
  NOR2_X1   g661(.A1(new_n686), .A2(new_n440), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n845), .A2(new_n725), .A3(new_n863), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n864), .A2(new_n315), .A3(new_n581), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT120), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n439), .A2(KEYINPUT57), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT55), .B1(new_n820), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n870), .B1(new_n869), .B2(new_n820), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n581), .A2(new_n871), .A3(new_n819), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n835), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n647), .ZN(new_n874));
  OR3_X1    g673(.A1(new_n837), .A2(new_n647), .A3(new_n823), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n613), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n840), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n868), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n440), .B1(new_n839), .B2(new_n840), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(KEYINPUT57), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n685), .A2(new_n842), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n880), .A2(new_n581), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(G141gat), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT58), .B1(new_n866), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT58), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n315), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n880), .A2(KEYINPUT119), .A3(new_n881), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT119), .B1(new_n880), .B2(new_n881), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n886), .B1(new_n889), .B2(new_n699), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n865), .B1(KEYINPUT120), .B2(new_n885), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n884), .B1(new_n890), .B2(new_n891), .ZN(G1344gat));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893));
  AOI211_X1 g692(.A(new_n893), .B(G148gat), .C1(new_n864), .C2(new_n666), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n693), .A2(new_n893), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n705), .B1(new_n835), .B2(new_n872), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n765), .B1(new_n896), .B2(new_n838), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n667), .A2(new_n582), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT57), .B1(new_n899), .B2(new_n439), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n867), .B1(new_n839), .B2(new_n840), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n881), .B(new_n895), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n887), .A2(new_n888), .A3(new_n693), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(KEYINPUT59), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n894), .B1(new_n904), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g704(.A(G155gat), .B1(new_n889), .B2(new_n692), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n864), .A2(new_n607), .A3(new_n613), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1346gat));
  AOI21_X1  g707(.A(G162gat), .B1(new_n864), .B2(new_n705), .ZN(new_n909));
  INV_X1    g708(.A(new_n889), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n705), .A2(G162gat), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(G1347gat));
  AOI21_X1  g711(.A(new_n669), .B1(new_n839), .B2(new_n840), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n310), .A3(new_n846), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT121), .ZN(new_n915));
  AOI21_X1  g714(.A(G169gat), .B1(new_n915), .B2(new_n700), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n725), .A2(new_n669), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n841), .A2(KEYINPUT122), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT122), .B1(new_n841), .B2(new_n917), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n582), .A2(new_n237), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n916), .B1(new_n920), .B2(new_n921), .ZN(G1348gat));
  AOI21_X1  g721(.A(new_n693), .B1(new_n251), .B2(new_n252), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n920), .A2(KEYINPUT123), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT123), .B1(new_n920), .B2(new_n923), .ZN(new_n925));
  AOI21_X1  g724(.A(G176gat), .B1(new_n915), .B2(new_n666), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(G1349gat));
  INV_X1    g726(.A(KEYINPUT60), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n928), .A2(KEYINPUT124), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n918), .A2(new_n919), .A3(new_n692), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n930), .A2(new_n242), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n613), .A2(new_n227), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n914), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n929), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n929), .ZN(new_n935));
  OAI221_X1 g734(.A(new_n935), .B1(new_n914), .B2(new_n932), .C1(new_n930), .C2(new_n242), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1350gat));
  NAND3_X1  g736(.A1(new_n915), .A2(new_n228), .A3(new_n705), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n920), .A2(new_n705), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(G190gat), .ZN(new_n941));
  AOI211_X1 g740(.A(KEYINPUT61), .B(new_n228), .C1(new_n920), .C2(new_n705), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(G1351gat));
  AND3_X1   g742(.A1(new_n913), .A2(new_n310), .A3(new_n863), .ZN(new_n944));
  INV_X1    g743(.A(G197gat), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n944), .A2(new_n945), .A3(new_n700), .ZN(new_n946));
  XOR2_X1   g745(.A(new_n946), .B(KEYINPUT125), .Z(new_n947));
  NAND2_X1  g746(.A1(new_n917), .A2(new_n685), .ZN(new_n948));
  OR3_X1    g747(.A1(new_n900), .A2(KEYINPUT126), .A3(new_n901), .ZN(new_n949));
  OAI21_X1  g748(.A(KEYINPUT126), .B1(new_n900), .B2(new_n901), .ZN(new_n950));
  AOI211_X1 g749(.A(new_n582), .B(new_n948), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n947), .B1(new_n945), .B2(new_n951), .ZN(G1352gat));
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n953));
  AOI21_X1  g752(.A(G204gat), .B1(new_n953), .B2(KEYINPUT62), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n944), .A2(new_n666), .A3(new_n954), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n955), .B(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n958), .A2(new_n666), .ZN(new_n959));
  INV_X1    g758(.A(G204gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(G1353gat));
  NAND3_X1  g760(.A1(new_n944), .A2(new_n212), .A3(new_n613), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n765), .A2(new_n948), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n963), .B1(new_n900), .B2(new_n901), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n964), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n964), .B2(G211gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(G1354gat));
  AOI21_X1  g766(.A(G218gat), .B1(new_n944), .B2(new_n705), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n647), .B1(new_n205), .B2(new_n206), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n958), .B2(new_n969), .ZN(G1355gat));
endmodule


