//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n786, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  INV_X1    g000(.A(KEYINPUT78), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G125), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT77), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n189), .A2(KEYINPUT77), .A3(G140), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n188), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n187), .B1(new_n196), .B2(new_n200), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n189), .A2(KEYINPUT77), .A3(G140), .ZN(new_n202));
  XNOR2_X1  g016(.A(G125), .B(G140), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(new_n193), .ZN(new_n204));
  OAI211_X1 g018(.A(KEYINPUT78), .B(new_n199), .C1(new_n204), .C2(new_n188), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n201), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n198), .B1(new_n196), .B2(new_n197), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT79), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT79), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n209), .B(new_n198), .C1(new_n196), .C2(new_n197), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n206), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n212));
  INV_X1    g026(.A(G119), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(G128), .ZN(new_n214));
  INV_X1    g028(.A(G128), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT23), .A3(G119), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n214), .B(new_n216), .C1(G119), .C2(new_n215), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT76), .ZN(new_n218));
  OR2_X1    g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G110), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n220), .B1(new_n217), .B2(new_n218), .ZN(new_n221));
  XNOR2_X1  g035(.A(G119), .B(G128), .ZN(new_n222));
  XOR2_X1   g036(.A(KEYINPUT24), .B(G110), .Z(new_n223));
  AOI22_X1  g037(.A1(new_n219), .A2(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n211), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n199), .B1(new_n204), .B2(new_n188), .ZN(new_n226));
  OAI22_X1  g040(.A1(new_n217), .A2(G110), .B1(new_n222), .B2(new_n223), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n203), .A2(new_n198), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT72), .A2(G953), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(KEYINPUT72), .A2(G953), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(G221), .A2(G234), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT80), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OR4_X1    g051(.A1(KEYINPUT80), .A2(new_n232), .A3(new_n233), .A4(new_n236), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT22), .B(G137), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n239), .B1(new_n237), .B2(new_n238), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT81), .ZN(new_n242));
  NOR3_X1   g056(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n237), .A2(new_n238), .ZN(new_n244));
  INV_X1    g058(.A(new_n239), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n247));
  AOI21_X1  g061(.A(KEYINPUT81), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(G902), .B1(new_n230), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n229), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n251), .B1(new_n211), .B2(new_n224), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n240), .A2(new_n241), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n252), .A2(KEYINPUT82), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT82), .B1(new_n252), .B2(new_n253), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n250), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT25), .ZN(new_n257));
  INV_X1    g071(.A(G217), .ZN(new_n258));
  INV_X1    g072(.A(G902), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n258), .B1(G234), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT25), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n250), .B(new_n261), .C1(new_n254), .C2(new_n255), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n257), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n255), .ZN(new_n264));
  INV_X1    g078(.A(new_n254), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n264), .A2(new_n265), .B1(new_n230), .B2(new_n249), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n260), .A2(G902), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT74), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT67), .ZN(new_n271));
  INV_X1    g085(.A(G137), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(KEYINPUT67), .A2(G137), .ZN(new_n274));
  AND2_X1   g088(.A1(KEYINPUT11), .A2(G134), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n272), .A2(G134), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT11), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT68), .B(G131), .ZN(new_n280));
  INV_X1    g094(.A(G134), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G137), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n276), .A2(new_n279), .A3(new_n280), .A4(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT69), .ZN(new_n284));
  INV_X1    g098(.A(G131), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT68), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G131), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n282), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT69), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n289), .A2(new_n290), .A3(new_n279), .A4(new_n276), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n293), .B1(new_n281), .B2(G137), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n272), .A2(KEYINPUT70), .A3(G134), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AND2_X1   g110(.A1(KEYINPUT67), .A2(G137), .ZN(new_n297));
  NOR2_X1   g111(.A1(KEYINPUT67), .A2(G137), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n281), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n285), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G143), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT1), .B1(new_n301), .B2(G146), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(G146), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n198), .A2(G143), .ZN(new_n304));
  OAI211_X1 g118(.A(G128), .B(new_n302), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n198), .A2(G143), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n301), .A2(G146), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n306), .B(new_n307), .C1(KEYINPUT1), .C2(new_n215), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n300), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n292), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT71), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n276), .A2(new_n279), .A3(new_n282), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G131), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n297), .A2(new_n298), .ZN(new_n316));
  AOI22_X1  g130(.A1(new_n316), .A2(new_n275), .B1(new_n278), .B2(new_n277), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n290), .B1(new_n317), .B2(new_n289), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n276), .A2(new_n279), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n282), .A2(new_n286), .A3(new_n288), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n319), .A2(KEYINPUT69), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n315), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(KEYINPUT0), .A2(G128), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n303), .A2(new_n304), .A3(new_n323), .ZN(new_n324));
  OAI22_X1  g138(.A1(new_n303), .A2(new_n304), .B1(KEYINPUT0), .B2(G128), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(KEYINPUT65), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT65), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(KEYINPUT0), .A3(G128), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT66), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n326), .A2(new_n328), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT66), .ZN(new_n332));
  NOR2_X1   g146(.A1(KEYINPUT0), .A2(G128), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n333), .B1(new_n306), .B2(new_n307), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n324), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n322), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n292), .A2(new_n310), .A3(KEYINPUT71), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n313), .A2(new_n337), .A3(KEYINPUT30), .A4(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n213), .A2(G116), .ZN(new_n340));
  INV_X1    g154(.A(G116), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G119), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  XOR2_X1   g158(.A(KEYINPUT2), .B(G113), .Z(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT2), .B(G113), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n284), .A2(new_n291), .B1(G131), .B2(new_n314), .ZN(new_n351));
  INV_X1    g165(.A(new_n324), .ZN(new_n352));
  XNOR2_X1  g166(.A(G143), .B(G146), .ZN(new_n353));
  NOR4_X1   g167(.A1(new_n329), .A2(new_n353), .A3(KEYINPUT66), .A4(new_n333), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n332), .B1(new_n331), .B2(new_n334), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n352), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n292), .A2(new_n310), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n350), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n339), .A2(new_n349), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n349), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n313), .A2(new_n337), .A3(new_n361), .A4(new_n338), .ZN(new_n362));
  INV_X1    g176(.A(G237), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n234), .A2(G210), .A3(new_n363), .ZN(new_n364));
  XOR2_X1   g178(.A(KEYINPUT73), .B(KEYINPUT27), .Z(new_n365));
  XNOR2_X1  g179(.A(new_n364), .B(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT26), .B(G101), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n366), .B(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT31), .B1(new_n360), .B2(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n311), .B(new_n361), .C1(new_n356), .C2(new_n351), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT28), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n349), .B1(new_n357), .B2(new_n358), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n373), .B(new_n374), .C1(new_n362), .C2(new_n372), .ZN(new_n375));
  INV_X1    g189(.A(new_n368), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n339), .A2(new_n349), .A3(new_n359), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT31), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n378), .A2(new_n379), .A3(new_n362), .A4(new_n368), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n370), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(G472), .A2(G902), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT32), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n270), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI211_X1 g199(.A(KEYINPUT74), .B(KEYINPUT32), .C1(new_n381), .C2(new_n382), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n375), .A2(new_n368), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n378), .A2(new_n362), .A3(new_n376), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT29), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n292), .A2(new_n310), .A3(KEYINPUT71), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT71), .B1(new_n292), .B2(new_n310), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n361), .B1(new_n395), .B2(new_n337), .ZN(new_n396));
  AND4_X1   g210(.A1(new_n361), .A2(new_n313), .A3(new_n337), .A4(new_n338), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT28), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n376), .A2(new_n391), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n373), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT75), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n398), .A2(KEYINPUT75), .A3(new_n373), .A4(new_n399), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n392), .A2(new_n402), .A3(new_n259), .A4(new_n403), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n381), .A2(new_n382), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n404), .A2(G472), .B1(new_n405), .B2(KEYINPUT32), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n269), .B1(new_n387), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT97), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT20), .ZN(new_n409));
  OR2_X1    g223(.A1(KEYINPUT72), .A2(G953), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n410), .A2(G214), .A3(new_n363), .A4(new_n231), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n411), .A2(new_n301), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n411), .A2(new_n301), .ZN(new_n413));
  OAI211_X1 g227(.A(KEYINPUT18), .B(G131), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n204), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n228), .B1(new_n415), .B2(new_n198), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n234), .A2(G143), .A3(G214), .A4(new_n363), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n411), .A2(new_n301), .ZN(new_n418));
  NAND2_X1  g232(.A1(KEYINPUT18), .A2(G131), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n414), .A2(new_n416), .A3(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(G113), .B(G122), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT93), .B(G104), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n422), .B(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n280), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n425), .B1(new_n412), .B2(new_n413), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT17), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n417), .A2(new_n418), .A3(new_n280), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n280), .B1(new_n417), .B2(new_n418), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n421), .B(new_n424), .C1(new_n432), .C2(new_n211), .ZN(new_n433));
  INV_X1    g247(.A(new_n428), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(new_n430), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT19), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(new_n194), .B2(new_n195), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n203), .A2(KEYINPUT19), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n226), .B1(new_n439), .B2(G146), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n421), .B1(new_n435), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n424), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n433), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(G475), .A2(G902), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n409), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n445), .ZN(new_n447));
  AOI211_X1 g261(.A(KEYINPUT20), .B(new_n447), .C1(new_n433), .C2(new_n443), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n421), .B1(new_n432), .B2(new_n211), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n442), .ZN(new_n450));
  AOI21_X1  g264(.A(G902), .B1(new_n450), .B2(new_n433), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT94), .B(G475), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  OAI22_X1  g267(.A1(new_n446), .A2(new_n448), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G122), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT14), .B1(new_n455), .B2(G116), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(KEYINPUT96), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n341), .A2(G122), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT14), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n455), .A2(G116), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G107), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n301), .A2(G128), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n215), .A2(G143), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT95), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(G128), .B(G143), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(KEYINPUT95), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n281), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n466), .A2(new_n467), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n469), .A2(KEYINPUT95), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n473), .A3(G134), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n458), .A2(new_n460), .ZN(new_n476));
  INV_X1    g290(.A(G107), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n463), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n476), .B(new_n477), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n469), .A2(KEYINPUT13), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n481), .B(G134), .C1(KEYINPUT13), .C2(new_n464), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n471), .A3(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT9), .B(G234), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n484), .A2(new_n258), .A3(G953), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n479), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n485), .B1(new_n479), .B2(new_n483), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n259), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G478), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n489), .A2(KEYINPUT15), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  OAI221_X1 g305(.A(new_n259), .B1(KEYINPUT15), .B2(new_n489), .C1(new_n486), .C2(new_n487), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n259), .B1(G234), .B2(G237), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n235), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT21), .B(G898), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G952), .ZN(new_n497));
  AOI211_X1 g311(.A(G953), .B(new_n497), .C1(G234), .C2(G237), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n491), .A2(new_n492), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n408), .B1(new_n454), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n447), .B1(new_n433), .B2(new_n443), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(new_n409), .ZN(new_n504));
  OR2_X1    g318(.A1(new_n451), .A2(new_n453), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n491), .A2(new_n492), .A3(new_n500), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .A4(KEYINPUT97), .ZN(new_n507));
  OAI21_X1  g321(.A(G214), .B1(G237), .B2(G902), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(G210), .B1(G237), .B2(G902), .ZN(new_n510));
  OAI211_X1 g324(.A(G125), .B(new_n352), .C1(new_n354), .C2(new_n355), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n309), .A2(G125), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(G953), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G224), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(KEYINPUT90), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n517), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n511), .B2(new_n513), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G104), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT3), .B1(new_n522), .B2(G107), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT3), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(new_n477), .A3(G104), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(G107), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT4), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n528), .A3(G101), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n527), .A2(G101), .ZN(new_n530));
  AOI21_X1  g344(.A(G101), .B1(new_n522), .B2(G107), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n523), .A2(new_n531), .A3(new_n525), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT4), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n349), .B(new_n529), .C1(new_n530), .C2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n344), .A2(KEYINPUT5), .ZN(new_n535));
  OAI21_X1  g349(.A(G113), .B1(new_n340), .B2(KEYINPUT5), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n523), .A2(new_n525), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT85), .B1(new_n477), .B2(G104), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT85), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(new_n522), .A3(G107), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n477), .A2(G104), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n539), .A2(new_n531), .B1(new_n544), .B2(G101), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n538), .A2(new_n545), .A3(new_n346), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n534), .A2(new_n546), .ZN(new_n547));
  XOR2_X1   g361(.A(G110), .B(G122), .Z(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n548), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n534), .A2(new_n550), .A3(new_n546), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(KEYINPUT6), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n534), .B2(new_n546), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT89), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT6), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n554), .B1(new_n553), .B2(new_n555), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n521), .B(new_n552), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n534), .A2(new_n546), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n516), .A2(KEYINPUT7), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n559), .A2(new_n550), .B1(new_n514), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT91), .B(KEYINPUT8), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n548), .B(new_n563), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n538), .A2(new_n346), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n544), .A2(G101), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n532), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n564), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT92), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n536), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n535), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n536), .A2(new_n569), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n346), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n545), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n512), .B1(new_n336), .B2(G125), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n568), .A2(new_n574), .B1(new_n575), .B2(new_n560), .ZN(new_n576));
  AOI21_X1  g390(.A(G902), .B1(new_n562), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n510), .B1(new_n558), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n558), .A2(new_n577), .A3(new_n510), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n509), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n502), .A2(new_n507), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G469), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT86), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n351), .A2(new_n584), .ZN(new_n585));
  AOI221_X4 g399(.A(KEYINPUT86), .B1(G131), .B2(new_n314), .C1(new_n284), .C2(new_n291), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n566), .A2(new_n308), .A3(new_n305), .A4(new_n532), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT10), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n305), .A2(new_n308), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n545), .A2(new_n591), .A3(KEYINPUT10), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n529), .B1(new_n530), .B2(new_n533), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n590), .B(new_n592), .C1(new_n356), .C2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT12), .ZN(new_n596));
  INV_X1    g410(.A(new_n588), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n566), .A2(new_n532), .B1(new_n308), .B2(new_n305), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n596), .B1(new_n599), .B2(new_n351), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n567), .A2(new_n309), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n588), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n602), .A2(new_n322), .A3(KEYINPUT12), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n587), .A2(new_n595), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(G110), .B(G140), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(KEYINPUT83), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n234), .A2(G227), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(KEYINPUT84), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n322), .A2(KEYINPUT86), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n351), .A2(new_n584), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n608), .B1(new_n612), .B2(new_n594), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n527), .A2(new_n528), .A3(G101), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n527), .A2(G101), .ZN(new_n615));
  INV_X1    g429(.A(new_n533), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n617), .A2(new_n336), .B1(new_n589), .B2(new_n588), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n351), .B1(new_n618), .B2(new_n592), .ZN(new_n619));
  OAI22_X1  g433(.A1(new_n604), .A2(new_n609), .B1(new_n613), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n583), .B1(new_n620), .B2(new_n259), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n602), .A2(new_n322), .A3(KEYINPUT12), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT12), .B1(new_n602), .B2(new_n322), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n613), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n618), .A2(new_n610), .A3(new_n592), .A4(new_n611), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n594), .A2(new_n322), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n608), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n583), .B(new_n259), .C1(new_n625), .C2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT87), .ZN(new_n630));
  INV_X1    g444(.A(new_n608), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n594), .A2(new_n585), .A3(new_n586), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n631), .B1(new_n632), .B2(new_n619), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n600), .A2(new_n603), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n634), .A2(new_n626), .A3(new_n608), .ZN(new_n635));
  AOI21_X1  g449(.A(G902), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT87), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n636), .A2(new_n637), .A3(new_n583), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n621), .B1(new_n630), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(G221), .B1(new_n484), .B2(G902), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(KEYINPUT88), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n613), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n634), .A2(new_n626), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT84), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n608), .B(new_n645), .ZN(new_n646));
  AOI22_X1  g460(.A1(new_n643), .A2(new_n627), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(G469), .B1(new_n647), .B2(G902), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n633), .A2(new_n635), .ZN(new_n649));
  AND4_X1   g463(.A1(new_n637), .A2(new_n649), .A3(new_n583), .A4(new_n259), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n637), .B1(new_n636), .B2(new_n583), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT88), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n652), .A2(new_n653), .A3(new_n640), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n582), .A2(new_n642), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n407), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G101), .ZN(G3));
  NAND2_X1  g471(.A1(new_n381), .A2(new_n259), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(G472), .ZN(new_n659));
  INV_X1    g473(.A(new_n260), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n256), .B2(KEYINPUT25), .ZN(new_n661));
  AOI22_X1  g475(.A1(new_n661), .A2(new_n262), .B1(new_n266), .B2(new_n267), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n659), .A2(new_n383), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n581), .A2(new_n500), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n489), .A2(new_n259), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n666), .B1(new_n488), .B2(G478), .ZN(new_n667));
  OAI21_X1  g481(.A(KEYINPUT33), .B1(new_n486), .B2(new_n487), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n479), .A2(new_n483), .ZN(new_n669));
  INV_X1    g483(.A(new_n485), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT33), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n479), .A2(new_n483), .A3(new_n485), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n667), .B1(G478), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n454), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n664), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n663), .A2(new_n642), .A3(new_n678), .A4(new_n654), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT34), .B(G104), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G6));
  AND2_X1   g495(.A1(new_n642), .A2(new_n654), .ZN(new_n682));
  INV_X1    g496(.A(new_n454), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n491), .A2(new_n492), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n664), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n682), .A2(new_n663), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT35), .B(G107), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G9));
  INV_X1    g503(.A(KEYINPUT99), .ZN(new_n690));
  INV_X1    g504(.A(new_n267), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n230), .A2(KEYINPUT98), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT36), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n693), .B1(new_n243), .B2(new_n248), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT98), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n252), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n692), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n252), .A2(new_n696), .ZN(new_n699));
  AOI211_X1 g513(.A(KEYINPUT98), .B(new_n251), .C1(new_n211), .C2(new_n224), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n694), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n691), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  AOI211_X1 g516(.A(new_n690), .B(new_n702), .C1(new_n661), .C2(new_n262), .ZN(new_n703));
  INV_X1    g517(.A(new_n702), .ZN(new_n704));
  AOI21_X1  g518(.A(KEYINPUT99), .B1(new_n263), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  AOI22_X1  g520(.A1(new_n658), .A2(G472), .B1(new_n382), .B2(new_n381), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n582), .A2(new_n642), .A3(new_n654), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT100), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT37), .B(G110), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G12));
  NAND2_X1  g527(.A1(new_n383), .A2(new_n384), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT74), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n404), .A2(G472), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n381), .A2(KEYINPUT32), .A3(new_n382), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n383), .A2(new_n270), .A3(new_n384), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n715), .A2(new_n716), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(G900), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n494), .A2(new_n720), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n721), .A2(KEYINPUT101), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(KEYINPUT101), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n722), .A2(new_n499), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n685), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n719), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n706), .A2(new_n642), .A3(new_n654), .A4(new_n581), .ZN(new_n727));
  OR2_X1    g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G128), .ZN(G30));
  XOR2_X1   g543(.A(new_n724), .B(KEYINPUT39), .Z(new_n730));
  NAND2_X1  g544(.A1(new_n682), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(KEYINPUT40), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n579), .A2(new_n580), .ZN(new_n733));
  XOR2_X1   g547(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n454), .A2(new_n684), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n735), .A2(new_n509), .A3(new_n736), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n396), .A2(new_n397), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n259), .B1(new_n738), .B2(new_n368), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n376), .B1(new_n378), .B2(new_n362), .ZN(new_n740));
  OAI21_X1  g554(.A(G472), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n715), .A2(new_n717), .A3(new_n718), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n263), .A2(new_n704), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n737), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT103), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n732), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n301), .ZN(G45));
  INV_X1    g564(.A(new_n724), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n454), .A2(new_n676), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n719), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n754), .A2(new_n727), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n198), .ZN(G48));
  NOR2_X1   g570(.A1(new_n636), .A2(new_n583), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n757), .B1(new_n630), .B2(new_n638), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n640), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n759), .B1(new_n387), .B2(new_n406), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n664), .A2(new_n269), .A3(new_n677), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(KEYINPUT41), .B(G113), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(G15));
  NOR3_X1   g578(.A1(new_n664), .A2(new_n269), .A3(new_n685), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n760), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G116), .ZN(G18));
  NAND3_X1  g581(.A1(new_n502), .A2(new_n507), .A3(new_n581), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n768), .A2(new_n703), .A3(new_n705), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n760), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G119), .ZN(G21));
  AND3_X1   g585(.A1(new_n558), .A2(new_n577), .A3(new_n510), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n508), .B1(new_n772), .B2(new_n578), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n736), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(new_n640), .A3(new_n500), .A4(new_n758), .ZN(new_n775));
  XNOR2_X1  g589(.A(KEYINPUT104), .B(G472), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n658), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n370), .A2(new_n380), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n368), .B1(new_n398), .B2(new_n373), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n382), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n777), .A2(new_n662), .A3(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n775), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n455), .ZN(G24));
  NOR2_X1   g597(.A1(new_n759), .A2(new_n773), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n777), .A2(new_n780), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(new_n743), .A3(new_n785), .A4(new_n753), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G125), .ZN(G27));
  NAND3_X1  g601(.A1(new_n716), .A2(new_n717), .A3(new_n714), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n579), .A2(new_n508), .A3(new_n580), .ZN(new_n789));
  NOR4_X1   g603(.A1(new_n639), .A2(new_n752), .A3(new_n789), .A4(new_n641), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n788), .A2(new_n790), .A3(new_n662), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n639), .A2(new_n641), .A3(new_n789), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT42), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n792), .A2(new_n793), .A3(new_n753), .ZN(new_n794));
  AOI22_X1  g608(.A1(KEYINPUT42), .A2(new_n791), .B1(new_n407), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G131), .ZN(G33));
  NAND3_X1  g610(.A1(new_n407), .A2(new_n725), .A3(new_n792), .ZN(new_n797));
  XNOR2_X1  g611(.A(KEYINPUT105), .B(G134), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n797), .B(new_n798), .ZN(G36));
  NAND2_X1  g613(.A1(new_n683), .A2(new_n676), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT43), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n801), .A2(new_n707), .A3(new_n744), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n789), .B1(new_n802), .B2(KEYINPUT44), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT107), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n647), .A2(KEYINPUT45), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n647), .A2(KEYINPUT45), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(G469), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(G469), .A2(G902), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(KEYINPUT46), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n630), .A2(new_n638), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(KEYINPUT106), .A3(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n807), .A2(new_n808), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n811), .B1(KEYINPUT46), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT106), .B1(new_n809), .B2(new_n810), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n815), .A2(new_n640), .A3(new_n730), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n804), .B(new_n817), .C1(KEYINPUT44), .C2(new_n802), .ZN(new_n818));
  XOR2_X1   g632(.A(KEYINPUT108), .B(G137), .Z(new_n819));
  XNOR2_X1  g633(.A(new_n818), .B(new_n819), .ZN(G39));
  NOR4_X1   g634(.A1(new_n719), .A2(new_n662), .A3(new_n752), .A4(new_n789), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n815), .A2(KEYINPUT47), .A3(new_n640), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT47), .B1(new_n815), .B2(new_n640), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n821), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT109), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT109), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n827), .B(new_n821), .C1(new_n823), .C2(new_n824), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(G140), .ZN(G42));
  AND4_X1   g644(.A1(new_n662), .A2(new_n642), .A3(new_n654), .A4(new_n707), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n831), .A2(new_n678), .B1(new_n407), .B2(new_n655), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT110), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n684), .B(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n683), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n664), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n659), .A2(new_n383), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n837), .A2(new_n703), .A3(new_n705), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n831), .A2(new_n836), .B1(new_n655), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT111), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n832), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n719), .A2(new_n662), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n679), .B1(new_n842), .B2(new_n709), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n663), .A2(new_n836), .A3(new_n642), .A4(new_n654), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n844), .B1(new_n709), .B2(new_n708), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT111), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n782), .B1(new_n760), .B2(new_n761), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n791), .A2(KEYINPUT42), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n407), .A2(new_n794), .ZN(new_n850));
  INV_X1    g664(.A(new_n759), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n719), .B(new_n851), .C1(new_n769), .C2(new_n765), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n848), .A2(new_n849), .A3(new_n850), .A4(new_n852), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n834), .A2(new_n789), .A3(new_n454), .A4(new_n724), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n682), .A2(new_n719), .A3(new_n706), .A4(new_n854), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n785), .A2(new_n743), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n790), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n797), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n853), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n786), .B1(new_n726), .B2(new_n727), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n860), .A2(new_n755), .ZN(new_n861));
  AND4_X1   g675(.A1(new_n640), .A2(new_n774), .A3(new_n652), .A4(new_n751), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n862), .A2(new_n742), .A3(new_n744), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT113), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n862), .A2(new_n742), .A3(KEYINPUT113), .A4(new_n744), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n861), .A2(KEYINPUT52), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT52), .B1(new_n861), .B2(new_n867), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n847), .B(new_n859), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n847), .A2(new_n859), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT52), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n754), .A2(new_n727), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n728), .A2(new_n875), .A3(new_n786), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n865), .A2(new_n866), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n861), .A2(KEYINPUT52), .A3(new_n867), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n873), .A2(KEYINPUT112), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT112), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n847), .A2(new_n859), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT53), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT114), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n872), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI211_X1 g699(.A(KEYINPUT114), .B(KEYINPUT53), .C1(new_n880), .C2(new_n882), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT54), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT116), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n858), .A2(new_n871), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n853), .A2(KEYINPUT115), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT115), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n795), .A2(new_n891), .A3(new_n848), .A4(new_n852), .ZN(new_n892));
  AND4_X1   g706(.A1(new_n847), .A2(new_n889), .A3(new_n890), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n878), .A2(new_n879), .ZN(new_n894));
  AOI22_X1  g708(.A1(new_n871), .A2(new_n870), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n888), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n870), .A2(new_n871), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n893), .A2(new_n894), .ZN(new_n899));
  AND4_X1   g713(.A1(new_n888), .A2(new_n898), .A3(new_n899), .A4(new_n896), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n887), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n789), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n498), .ZN(new_n904));
  NOR4_X1   g718(.A1(new_n742), .A2(new_n269), .A3(new_n759), .A4(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n454), .A2(new_n676), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n801), .A2(new_n499), .A3(new_n781), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n908), .A2(new_n509), .A3(new_n735), .A4(new_n851), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT50), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n801), .A2(new_n759), .A3(new_n904), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT119), .ZN(new_n912));
  AOI211_X1 g726(.A(new_n907), .B(new_n910), .C1(new_n856), .C2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n758), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n914), .A2(KEYINPUT118), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(KEYINPUT118), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n915), .A2(new_n916), .A3(new_n640), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n823), .A2(new_n824), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n908), .A2(new_n903), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT117), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT51), .B1(new_n913), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n269), .B1(new_n406), .B2(new_n714), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n912), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT48), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n905), .A2(new_n454), .A3(new_n676), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n908), .A2(new_n784), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n926), .A2(new_n927), .A3(G952), .A4(new_n515), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT120), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n925), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n922), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n913), .A2(new_n921), .A3(KEYINPUT51), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI22_X1  g749(.A1(new_n902), .A2(new_n935), .B1(G952), .B2(G953), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n914), .A2(KEYINPUT49), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n937), .A2(new_n735), .ZN(new_n938));
  NOR4_X1   g752(.A1(new_n269), .A2(new_n800), .A3(new_n641), .A4(new_n509), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n938), .B(new_n939), .C1(KEYINPUT49), .C2(new_n914), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n936), .B1(new_n742), .B2(new_n940), .ZN(G75));
  NOR2_X1   g755(.A1(new_n895), .A2(new_n259), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(G210), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT56), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(KEYINPUT55), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n552), .B1(new_n556), .B2(new_n557), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(new_n521), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT55), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n943), .A2(new_n949), .A3(new_n944), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n946), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n948), .B1(new_n946), .B2(new_n950), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n235), .A2(new_n497), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT121), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n951), .A2(new_n952), .A3(new_n955), .ZN(G51));
  XNOR2_X1  g770(.A(new_n895), .B(new_n896), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n808), .B(KEYINPUT57), .Z(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n649), .ZN(new_n960));
  OR3_X1    g774(.A1(new_n895), .A2(new_n259), .A3(new_n807), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n955), .B1(new_n960), .B2(new_n961), .ZN(G54));
  AND2_X1   g776(.A1(KEYINPUT58), .A2(G475), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n942), .A2(new_n963), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n964), .A2(new_n444), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n964), .A2(new_n444), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n954), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT122), .ZN(G60));
  XNOR2_X1  g782(.A(new_n665), .B(KEYINPUT59), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n675), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n955), .B1(new_n957), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n969), .B1(new_n887), .B2(new_n901), .ZN(new_n972));
  INV_X1    g786(.A(new_n675), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(KEYINPUT123), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT123), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n976), .B(new_n971), .C1(new_n972), .C2(new_n973), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(G63));
  NAND2_X1  g792(.A1(G217), .A2(G902), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT60), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n895), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n954), .B1(new_n981), .B2(new_n266), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n698), .A2(new_n701), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n982), .B1(new_n983), .B2(new_n981), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT61), .ZN(G66));
  INV_X1    g799(.A(G224), .ZN(new_n986));
  OAI21_X1  g800(.A(G953), .B1(new_n495), .B2(new_n986), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n847), .A2(new_n848), .A3(new_n852), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n987), .B1(new_n988), .B2(new_n235), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n947), .B1(G898), .B2(new_n234), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT124), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n989), .B(new_n991), .ZN(G69));
  AND2_X1   g806(.A1(new_n829), .A2(new_n818), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n923), .A2(new_n774), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n795), .B(new_n797), .C1(new_n816), .C2(new_n994), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n995), .A2(new_n876), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n339), .A2(new_n359), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(new_n439), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n999), .A2(new_n234), .ZN(new_n1000));
  AOI22_X1  g814(.A1(new_n997), .A2(new_n1000), .B1(new_n720), .B2(new_n235), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n749), .A2(new_n876), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT62), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n789), .B1(new_n835), .B2(new_n677), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n407), .A2(new_n682), .A3(new_n730), .A4(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n993), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n1006), .A2(new_n234), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1001), .B1(new_n1007), .B2(new_n999), .ZN(new_n1008));
  INV_X1    g822(.A(G227), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n235), .B1(new_n1009), .B2(new_n720), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1010), .B(KEYINPUT125), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1008), .B(new_n1012), .ZN(G72));
  NAND4_X1  g827(.A1(new_n829), .A2(new_n818), .A3(new_n988), .A4(new_n996), .ZN(new_n1014));
  NAND2_X1  g828(.A1(G472), .A2(G902), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1015), .B(KEYINPUT63), .Z(new_n1016));
  NAND2_X1  g830(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n389), .B(KEYINPUT126), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n955), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(KEYINPUT127), .ZN(new_n1020));
  INV_X1    g834(.A(new_n740), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n993), .A2(new_n988), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1021), .B1(new_n1022), .B2(new_n1016), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n885), .A2(new_n886), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1021), .A2(new_n389), .A3(new_n1016), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NOR3_X1   g840(.A1(new_n1020), .A2(new_n1023), .A3(new_n1026), .ZN(G57));
endmodule


