//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1264, new_n1265, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n201), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT64), .B(G238), .ZN(new_n216));
  AND2_X1   g0016(.A1(new_n216), .A2(G68), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G107), .A2(G264), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n209), .B1(new_n213), .B2(new_n215), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT65), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n230), .B(new_n233), .Z(G358));
  XOR2_X1   g0034(.A(G58), .B(G77), .Z(new_n235));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G87), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G97), .B(G107), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G351));
  NAND2_X1  g0041(.A1(KEYINPUT67), .A2(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT8), .ZN(new_n243));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  NOR2_X1   g0044(.A1(new_n244), .A2(G20), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NOR2_X1   g0046(.A1(G20), .A2(G33), .ZN(new_n247));
  AOI22_X1  g0047(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n210), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G13), .A3(G20), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(G50), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n251), .B1(new_n253), .B2(G20), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n255), .B1(new_n256), .B2(G50), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(G1), .A2(G13), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  OAI21_X1  g0064(.A(KEYINPUT66), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n244), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT66), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G77), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n262), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G222), .A2(G1698), .ZN(new_n274));
  INV_X1    g0074(.A(G223), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n274), .B1(new_n275), .B2(G1698), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n273), .B1(new_n271), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G45), .ZN(new_n279));
  AOI21_X1  g0079(.A(G1), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n262), .A2(G274), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n262), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n282), .B1(G226), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n277), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(G169), .ZN(new_n289));
  INV_X1    g0089(.A(G179), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n290), .A2(KEYINPUT68), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(KEYINPUT68), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI211_X1 g0093(.A(new_n259), .B(new_n289), .C1(new_n293), .C2(new_n288), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n258), .B(KEYINPUT9), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n288), .A2(G190), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n287), .A2(G200), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT10), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n295), .A2(new_n300), .A3(new_n296), .A4(new_n297), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n294), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n281), .A2(KEYINPUT70), .ZN(new_n303));
  INV_X1    g0103(.A(G274), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(new_n260), .B2(new_n261), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT70), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n305), .A2(new_n306), .A3(new_n280), .ZN(new_n307));
  INV_X1    g0107(.A(G238), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n303), .B(new_n307), .C1(new_n308), .C2(new_n284), .ZN(new_n309));
  MUX2_X1   g0109(.A(G226), .B(G232), .S(G1698), .Z(new_n310));
  NAND3_X1  g0110(.A1(new_n310), .A2(new_n265), .A3(new_n270), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G97), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n262), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT13), .B1(new_n309), .B2(new_n313), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n281), .A2(KEYINPUT70), .B1(new_n284), .B2(new_n308), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n306), .B1(new_n305), .B2(new_n280), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n311), .A2(new_n312), .ZN(new_n318));
  INV_X1    g0118(.A(new_n262), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT13), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n317), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n314), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G169), .ZN(new_n324));
  OAI211_X1 g0124(.A(KEYINPUT71), .B(KEYINPUT14), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT71), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n324), .B1(new_n314), .B2(new_n322), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT14), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n323), .A2(G179), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT72), .B(KEYINPUT14), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n325), .A2(new_n329), .A3(new_n330), .A4(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n256), .ZN(new_n334));
  INV_X1    g0134(.A(G68), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT12), .ZN(new_n336));
  INV_X1    g0136(.A(new_n254), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(new_n335), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n254), .A2(KEYINPUT12), .A3(G68), .ZN(new_n339));
  OAI22_X1  g0139(.A1(new_n334), .A2(new_n335), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n247), .A2(G50), .B1(G20), .B2(new_n335), .ZN(new_n341));
  INV_X1    g0141(.A(new_n245), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n341), .B1(new_n342), .B2(new_n272), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n343), .A2(KEYINPUT11), .A3(new_n251), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT11), .B1(new_n343), .B2(new_n251), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n340), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n333), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n314), .A2(new_n322), .A3(G190), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n346), .ZN(new_n350));
  INV_X1    g0150(.A(G200), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n351), .B1(new_n314), .B2(new_n322), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n337), .A2(new_n272), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(new_n334), .B2(new_n272), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT8), .B(G58), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n358), .A2(new_n247), .B1(G20), .B2(G77), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT15), .B(G87), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n359), .B1(new_n342), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n356), .B1(new_n251), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n271), .ZN(new_n364));
  NOR2_X1   g0164(.A1(G232), .A2(G1698), .ZN(new_n365));
  INV_X1    g0165(.A(G1698), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n216), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n364), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n368), .B(new_n319), .C1(G107), .C2(new_n364), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n282), .B1(G244), .B2(new_n285), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G190), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n363), .B1(new_n373), .B2(KEYINPUT69), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n351), .B1(new_n369), .B2(new_n370), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT69), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n375), .A2(new_n376), .B1(new_n371), .B2(new_n372), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n369), .A2(new_n293), .A3(new_n370), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n362), .B1(new_n371), .B2(new_n324), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n374), .A2(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n302), .A2(new_n348), .A3(new_n354), .A4(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n243), .A2(new_n337), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n334), .B2(new_n243), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n275), .A2(new_n366), .ZN(new_n385));
  OAI221_X1 g0185(.A(new_n385), .B1(G226), .B2(new_n366), .C1(new_n263), .C2(new_n264), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G87), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n319), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n262), .A2(G232), .A3(new_n283), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n281), .A2(new_n390), .A3(KEYINPUT73), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT73), .B1(new_n281), .B2(new_n390), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n389), .B(new_n372), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n262), .B1(new_n386), .B2(new_n387), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n281), .A2(new_n390), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n351), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n263), .A2(new_n264), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n398), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n399));
  AOI21_X1  g0199(.A(G20), .B1(new_n265), .B2(new_n270), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n399), .B1(new_n400), .B2(KEYINPUT7), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G68), .ZN(new_n402));
  INV_X1    g0202(.A(G58), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(new_n335), .ZN(new_n404));
  OAI21_X1  g0204(.A(G20), .B1(new_n404), .B2(new_n201), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n247), .A2(G159), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT16), .B1(new_n402), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n267), .A2(new_n269), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT7), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n410), .A2(new_n411), .A3(G20), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT7), .B1(new_n398), .B2(new_n211), .ZN(new_n413));
  OAI21_X1  g0213(.A(G68), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n414), .A2(KEYINPUT16), .A3(new_n408), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n251), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n384), .B(new_n397), .C1(new_n409), .C2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n251), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n411), .B1(new_n410), .B2(G20), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n399), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n407), .B1(new_n422), .B2(G68), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n420), .B1(new_n423), .B2(KEYINPUT16), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n407), .B1(new_n401), .B2(G68), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n424), .B1(KEYINPUT16), .B2(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n426), .A2(KEYINPUT17), .A3(new_n384), .A4(new_n397), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n419), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT74), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT18), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n384), .B1(new_n409), .B2(new_n416), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n389), .B(new_n293), .C1(new_n391), .C2(new_n392), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n324), .B1(new_n394), .B2(new_n395), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n431), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n428), .A2(new_n437), .ZN(new_n438));
  AOI211_X1 g0238(.A(KEYINPUT18), .B(new_n435), .C1(new_n426), .C2(new_n384), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n430), .B1(new_n432), .B2(new_n436), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT74), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n381), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n247), .A2(G77), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT6), .ZN(new_n445));
  INV_X1    g0245(.A(G97), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n445), .A2(new_n446), .A3(G107), .ZN(new_n447));
  XNOR2_X1  g0247(.A(G97), .B(G107), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n447), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n444), .B1(new_n449), .B2(new_n211), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n450), .B1(new_n401), .B2(G107), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n253), .A2(G33), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n254), .A2(new_n452), .A3(new_n210), .A4(new_n250), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G97), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n254), .A2(new_n446), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT75), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n454), .A2(KEYINPUT75), .A3(new_n455), .ZN(new_n457));
  OAI22_X1  g0257(.A1(new_n451), .A2(new_n420), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n279), .A2(G1), .ZN(new_n459));
  XNOR2_X1  g0259(.A(KEYINPUT5), .B(G41), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n305), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  AND2_X1   g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  NOR2_X1   g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n262), .ZN(new_n465));
  INV_X1    g0265(.A(G257), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(G244), .B(new_n366), .C1(new_n263), .C2(new_n264), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT4), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT76), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G33), .A2(G283), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT76), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n468), .A2(new_n473), .A3(new_n469), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G250), .A2(G1698), .ZN(new_n475));
  NAND2_X1  g0275(.A1(KEYINPUT4), .A2(G244), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n475), .B1(new_n476), .B2(G1698), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n265), .A2(new_n270), .A3(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n471), .A2(new_n472), .A3(new_n474), .A4(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n467), .B1(new_n479), .B2(new_n319), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n293), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n458), .B(new_n481), .C1(G169), .C2(new_n480), .ZN(new_n482));
  INV_X1    g0282(.A(new_n467), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n478), .A2(new_n472), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n468), .A2(new_n473), .A3(new_n469), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n473), .B1(new_n468), .B2(new_n469), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n483), .B1(new_n487), .B2(new_n262), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G200), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n457), .A2(new_n456), .ZN(new_n490));
  INV_X1    g0290(.A(new_n450), .ZN(new_n491));
  NOR3_X1   g0291(.A1(new_n263), .A2(new_n264), .A3(KEYINPUT66), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n268), .B1(new_n267), .B2(new_n269), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n211), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n412), .B1(new_n494), .B2(new_n411), .ZN(new_n495));
  INV_X1    g0295(.A(G107), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n491), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n490), .B1(new_n497), .B2(new_n251), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n480), .A2(G190), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n489), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(G250), .B(new_n366), .C1(new_n263), .C2(new_n264), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT85), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n410), .A2(KEYINPUT85), .A3(G250), .A4(new_n366), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(G257), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G294), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n465), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n510), .A2(new_n319), .B1(G264), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(G190), .A3(new_n461), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(G264), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n508), .B1(new_n504), .B2(new_n503), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n461), .B(new_n514), .C1(new_n515), .C2(new_n262), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G200), .ZN(new_n517));
  INV_X1    g0317(.A(G87), .ZN(new_n518));
  NOR3_X1   g0318(.A1(new_n518), .A2(KEYINPUT22), .A3(G20), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n265), .A2(new_n270), .A3(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n211), .B(G87), .C1(new_n263), .C2(new_n264), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT22), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT24), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT23), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n211), .B2(G107), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n496), .A2(KEYINPUT23), .A3(G20), .ZN(new_n527));
  INV_X1    g0327(.A(G116), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n244), .A2(new_n528), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n526), .A2(new_n527), .B1(new_n529), .B2(new_n211), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n523), .A2(new_n524), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n524), .B1(new_n523), .B2(new_n530), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n251), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT25), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n254), .B2(G107), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NOR3_X1   g0337(.A1(new_n254), .A2(new_n535), .A3(G107), .ZN(new_n538));
  OAI22_X1  g0338(.A1(new_n537), .A2(new_n538), .B1(new_n496), .B2(new_n453), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n513), .A2(new_n517), .A3(new_n534), .A4(new_n540), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n482), .A2(new_n500), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n308), .A2(new_n366), .ZN(new_n543));
  INV_X1    g0343(.A(G244), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G1698), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n543), .B(new_n545), .C1(new_n263), .C2(new_n264), .ZN(new_n546));
  INV_X1    g0346(.A(new_n529), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n262), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n262), .A2(G274), .A3(new_n459), .ZN(new_n549));
  INV_X1    g0349(.A(G250), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(new_n253), .B2(G45), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n262), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(G169), .B1(new_n548), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT77), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n305), .A2(new_n459), .B1(new_n262), .B2(new_n551), .ZN(new_n556));
  INV_X1    g0356(.A(new_n293), .ZN(new_n557));
  NOR2_X1   g0357(.A1(G238), .A2(G1698), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n558), .B1(new_n544), .B2(G1698), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n529), .B1(new_n559), .B2(new_n410), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n556), .B(new_n557), .C1(new_n560), .C2(new_n262), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n554), .A2(new_n555), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n555), .B1(new_n554), .B2(new_n561), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n360), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n565), .A2(new_n254), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n211), .B(G68), .C1(new_n263), .C2(new_n264), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT79), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT79), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n410), .A2(new_n569), .A3(new_n211), .A4(G68), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(KEYINPUT19), .B1(new_n245), .B2(G97), .ZN(new_n572));
  OR2_X1    g0372(.A1(KEYINPUT78), .A2(G87), .ZN(new_n573));
  NAND2_X1  g0373(.A1(KEYINPUT78), .A2(G87), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n573), .A2(new_n446), .A3(new_n496), .A4(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT19), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n312), .B2(new_n211), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n572), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n571), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n566), .B1(new_n579), .B2(new_n251), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n453), .A2(new_n360), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT80), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n420), .B1(new_n571), .B2(new_n578), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT80), .ZN(new_n585));
  NOR4_X1   g0385(.A1(new_n584), .A2(new_n585), .A3(new_n566), .A4(new_n581), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n564), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  OR2_X1    g0387(.A1(new_n453), .A2(new_n518), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n580), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n556), .B1(new_n560), .B2(new_n262), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G200), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n372), .B2(new_n590), .ZN(new_n592));
  OR2_X1    g0392(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n510), .A2(new_n319), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n594), .A2(new_n290), .A3(new_n461), .A4(new_n514), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n516), .A2(new_n324), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n523), .A2(new_n530), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT24), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n420), .B1(new_n598), .B2(new_n531), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n595), .B(new_n596), .C1(new_n599), .C2(new_n539), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n587), .A2(new_n593), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n542), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n337), .A2(new_n528), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n453), .B2(new_n528), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n250), .A2(new_n210), .B1(G20), .B2(new_n528), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n472), .B(new_n211), .C1(G33), .C2(new_n446), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT20), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n606), .A2(KEYINPUT20), .A3(new_n607), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n605), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n464), .A2(G270), .A3(new_n262), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT81), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n611), .A2(new_n612), .A3(new_n461), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n612), .B1(new_n611), .B2(new_n461), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(G264), .A2(G1698), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n271), .A2(G303), .B1(new_n410), .B2(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(G257), .B(new_n366), .C1(new_n263), .C2(new_n264), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT82), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n410), .A2(KEYINPUT82), .A3(G257), .A4(new_n366), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n262), .B1(new_n617), .B2(new_n622), .ZN(new_n623));
  OAI211_X1 g0423(.A(G169), .B(new_n610), .C1(new_n615), .C2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT21), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n271), .A2(G303), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n410), .A2(new_n616), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n622), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n319), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n611), .A2(new_n461), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT81), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n611), .A2(new_n461), .A3(new_n612), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n610), .A2(G179), .ZN(new_n635));
  OAI22_X1  g0435(.A1(new_n624), .A2(new_n625), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n609), .A2(new_n608), .ZN(new_n637));
  OAI21_X1  g0437(.A(G169), .B1(new_n637), .B2(new_n604), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n629), .B2(new_n633), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT83), .B1(new_n639), .B2(KEYINPUT21), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT83), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n624), .A2(new_n641), .A3(new_n625), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n636), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT84), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n634), .A2(G200), .ZN(new_n645));
  INV_X1    g0445(.A(new_n610), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n645), .B(new_n646), .C1(new_n372), .C2(new_n634), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n643), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n635), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n615), .A2(new_n623), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n639), .A2(KEYINPUT21), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n639), .A2(KEYINPUT83), .A3(KEYINPUT21), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n641), .B1(new_n624), .B2(new_n625), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n647), .B(new_n651), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(KEYINPUT84), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n602), .B1(new_n648), .B2(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n443), .A2(new_n656), .ZN(G372));
  NAND2_X1  g0457(.A1(new_n299), .A2(new_n301), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n379), .A2(new_n378), .ZN(new_n659));
  AOI211_X1 g0459(.A(new_n428), .B(new_n353), .C1(new_n348), .C2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n408), .B1(new_n495), .B2(new_n335), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT16), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n383), .B1(new_n663), .B2(new_n424), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT18), .B1(new_n664), .B2(new_n435), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n432), .A2(new_n436), .A3(new_n430), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n658), .B1(new_n660), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n294), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT26), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n554), .A2(new_n561), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n583), .B2(new_n586), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT86), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n593), .B(new_n673), .C1(new_n482), .C2(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n482), .A2(new_n674), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n671), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n587), .A2(new_n593), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n482), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(KEYINPUT26), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n673), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n643), .A2(new_n600), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n482), .A2(new_n500), .A3(new_n541), .ZN(new_n684));
  INV_X1    g0484(.A(new_n593), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n682), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n443), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n670), .A2(new_n689), .ZN(G369));
  NAND3_X1  g0490(.A1(new_n253), .A2(new_n211), .A3(G13), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G213), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g0494(.A(KEYINPUT87), .B(G343), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n646), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n698), .B1(new_n655), .B2(new_n648), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n700), .A2(new_n698), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n600), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n697), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n696), .B1(new_n599), .B2(new_n539), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n541), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n704), .B1(new_n706), .B2(new_n703), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n702), .A2(G330), .A3(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n700), .A2(new_n706), .A3(new_n600), .A4(new_n697), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n704), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n709), .A2(new_n712), .ZN(G399));
  INV_X1    g0513(.A(new_n207), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G41), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G1), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n575), .A2(G116), .ZN(new_n718));
  OAI22_X1  g0518(.A1(new_n717), .A2(new_n718), .B1(new_n215), .B2(new_n716), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  AOI211_X1 g0520(.A(KEYINPUT29), .B(new_n696), .C1(new_n681), .C2(new_n687), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT29), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n683), .A2(new_n686), .ZN(new_n723));
  OAI21_X1  g0523(.A(KEYINPUT26), .B1(new_n675), .B2(new_n676), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n679), .A2(new_n671), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n723), .A2(new_n724), .A3(new_n673), .A4(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n722), .B1(new_n726), .B2(new_n697), .ZN(new_n727));
  INV_X1    g0527(.A(G330), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n684), .A2(new_n678), .A3(new_n703), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n654), .A2(KEYINPUT84), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n644), .B1(new_n643), .B2(new_n647), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n729), .B(new_n697), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n590), .A2(new_n290), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n512), .A2(new_n629), .A3(new_n633), .A4(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n733), .B1(new_n735), .B2(new_n488), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n590), .A2(new_n293), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n488), .A2(new_n634), .A3(new_n516), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT88), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AND3_X1   g0541(.A1(new_n629), .A2(new_n633), .A3(new_n734), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(KEYINPUT30), .A3(new_n480), .A4(new_n512), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n736), .A2(KEYINPUT88), .A3(new_n738), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n741), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT31), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n697), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n736), .A2(new_n743), .A3(new_n738), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n696), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n745), .A2(new_n747), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n728), .B1(new_n732), .B2(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n721), .A2(new_n727), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n720), .B1(new_n752), .B2(G1), .ZN(G364));
  NAND2_X1  g0553(.A1(new_n702), .A2(G330), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n211), .A2(G13), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n253), .B1(new_n755), .B2(G45), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n715), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n699), .A2(new_n701), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(new_n728), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n754), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT89), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n762), .B(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n210), .B1(G20), .B2(new_n324), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n211), .A2(G190), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n767), .A2(new_n290), .A3(G200), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT91), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G283), .ZN(new_n774));
  INV_X1    g0574(.A(G311), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n293), .A2(new_n211), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G190), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n773), .A2(new_n774), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  AND3_X1   g0579(.A1(new_n290), .A2(new_n351), .A3(KEYINPUT90), .ZN(new_n780));
  AOI21_X1  g0580(.A(KEYINPUT90), .B1(new_n290), .B2(new_n351), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n767), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n779), .B1(G329), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G303), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n290), .A2(G20), .A3(G190), .A4(G200), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n211), .A2(new_n372), .A3(G200), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n557), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G322), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n271), .B1(new_n785), .B2(new_n786), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n776), .A2(G190), .A3(G200), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n790), .B1(G326), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n780), .A2(new_n781), .ZN(new_n794));
  OAI21_X1  g0594(.A(G20), .B1(new_n794), .B2(new_n372), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G294), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n776), .A2(new_n372), .A3(G200), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT94), .B(KEYINPUT33), .ZN(new_n799));
  INV_X1    g0599(.A(G317), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n784), .A2(new_n793), .A3(new_n796), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n772), .A2(G107), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n786), .B1(new_n573), .B2(new_n574), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n271), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT92), .Z(new_n808));
  INV_X1    g0608(.A(G159), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n782), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT32), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n778), .A2(new_n272), .B1(new_n788), .B2(new_n403), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G50), .B2(new_n792), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n808), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n795), .A2(G97), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n797), .B2(new_n335), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT93), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n803), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n766), .B1(new_n818), .B2(KEYINPUT95), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(KEYINPUT95), .B2(new_n818), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n271), .A2(new_n714), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n821), .A2(G355), .B1(new_n528), .B2(new_n714), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n237), .A2(new_n279), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n714), .A2(new_n410), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(G45), .B2(new_n215), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n822), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(G13), .A2(G33), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(G20), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(new_n765), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n759), .B1(new_n826), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n829), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n820), .B(new_n831), .C1(new_n702), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n764), .A2(new_n833), .ZN(G396));
  NAND2_X1  g0634(.A1(new_n688), .A2(new_n697), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n363), .A2(new_n696), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT97), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n659), .B2(new_n697), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n379), .A2(KEYINPUT97), .A3(new_n378), .A4(new_n696), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n380), .A2(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n380), .A2(new_n836), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n838), .A2(new_n839), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n688), .A2(new_n697), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n751), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n758), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n847), .B2(new_n846), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n765), .A2(new_n827), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n759), .B1(new_n272), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n772), .A2(G87), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n852), .B1(new_n528), .B2(new_n778), .C1(new_n775), .C2(new_n782), .ZN(new_n853));
  INV_X1    g0653(.A(new_n786), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n364), .B1(G107), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(G294), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n855), .B(new_n815), .C1(new_n856), .C2(new_n788), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n774), .A2(new_n797), .B1(new_n791), .B2(new_n785), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n853), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n778), .ZN(new_n860));
  INV_X1    g0660(.A(new_n788), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n860), .A2(G159), .B1(new_n861), .B2(G143), .ZN(new_n862));
  INV_X1    g0662(.A(G137), .ZN(new_n863));
  INV_X1    g0663(.A(G150), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n862), .B1(new_n863), .B2(new_n791), .C1(new_n864), .C2(new_n797), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT34), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n410), .B1(new_n786), .B2(new_n202), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n772), .B2(G68), .ZN(new_n868));
  INV_X1    g0668(.A(new_n795), .ZN(new_n869));
  INV_X1    g0669(.A(G132), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n868), .B1(new_n403), .B2(new_n869), .C1(new_n870), .C2(new_n782), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT96), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n859), .B1(new_n866), .B2(new_n872), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n851), .B1(new_n766), .B2(new_n873), .C1(new_n844), .C2(new_n828), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n849), .A2(new_n874), .ZN(G384));
  NAND2_X1  g0675(.A1(new_n448), .A2(new_n445), .ZN(new_n876));
  INV_X1    g0676(.A(new_n447), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n528), .B(new_n213), .C1(new_n878), .C2(KEYINPUT35), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(KEYINPUT35), .B2(new_n878), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT36), .Z(new_n881));
  OR3_X1    g0681(.A1(new_n215), .A2(new_n272), .A3(new_n404), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n335), .A2(G50), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT98), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n253), .B(G13), .C1(new_n882), .C2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n423), .A2(KEYINPUT16), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n384), .B1(new_n416), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n694), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(new_n438), .B2(new_n441), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n888), .B1(new_n436), .B2(new_n889), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n417), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(KEYINPUT37), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n432), .A2(new_n436), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n432), .A2(new_n889), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT37), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n895), .A2(new_n896), .A3(new_n897), .A4(new_n417), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT38), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n891), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n665), .A2(new_n666), .A3(new_n419), .A4(new_n427), .ZN(new_n902));
  INV_X1    g0702(.A(new_n896), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT99), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n895), .A2(new_n896), .A3(new_n417), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT37), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n898), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n902), .A2(KEYINPUT99), .A3(new_n903), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n906), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n901), .B1(new_n900), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n749), .A2(new_n746), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n748), .A2(KEYINPUT31), .A3(new_n696), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n732), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n346), .A2(new_n697), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n348), .A2(new_n354), .A3(new_n918), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n347), .B(new_n696), .C1(new_n333), .C2(new_n353), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n840), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n916), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT40), .B1(new_n912), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n913), .A2(new_n914), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n656), .B2(new_n697), .ZN(new_n925));
  INV_X1    g0725(.A(new_n920), .ZN(new_n926));
  AOI211_X1 g0726(.A(new_n353), .B(new_n917), .C1(new_n333), .C2(new_n347), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n844), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT40), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n900), .B1(new_n891), .B2(new_n899), .ZN(new_n931));
  INV_X1    g0731(.A(new_n890), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n429), .B1(new_n665), .B2(new_n666), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n435), .B1(new_n426), .B2(new_n384), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n419), .B(new_n427), .C1(new_n934), .C2(new_n431), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n932), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n894), .A2(new_n898), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(KEYINPUT38), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n931), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n929), .A2(new_n930), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n923), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT100), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n925), .A2(new_n381), .A3(new_n442), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n944), .A2(new_n945), .A3(new_n728), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n659), .A2(new_n696), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n845), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n926), .A2(new_n927), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n949), .A2(new_n939), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n667), .A2(new_n694), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n910), .A2(new_n909), .ZN(new_n955));
  AOI21_X1  g0755(.A(KEYINPUT99), .B1(new_n902), .B2(new_n903), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n900), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(KEYINPUT39), .B1(new_n957), .B2(new_n938), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n931), .A2(KEYINPUT39), .A3(new_n938), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n348), .A2(new_n696), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n958), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n954), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n443), .B1(new_n721), .B2(new_n727), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n670), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n964), .B(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(KEYINPUT101), .B1(new_n946), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n946), .A2(new_n967), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n968), .B(new_n969), .C1(new_n253), .C2(new_n755), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n946), .A2(KEYINPUT101), .A3(new_n967), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n886), .B1(new_n970), .B2(new_n971), .ZN(G367));
  NAND2_X1  g0772(.A1(new_n233), .A2(new_n824), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n973), .B(new_n830), .C1(new_n207), .C2(new_n360), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n772), .A2(G97), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n975), .B(new_n398), .C1(new_n856), .C2(new_n797), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(G107), .B2(new_n795), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n791), .A2(new_n775), .B1(new_n785), .B2(new_n788), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT104), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n860), .A2(G283), .B1(G317), .B2(new_n783), .ZN(new_n980));
  OAI21_X1  g0780(.A(KEYINPUT105), .B1(new_n786), .B2(new_n528), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT46), .Z(new_n982));
  NAND4_X1  g0782(.A1(new_n977), .A2(new_n979), .A3(new_n980), .A4(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT106), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n792), .A2(G143), .B1(G150), .B2(new_n861), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n869), .A2(new_n335), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n988), .A2(KEYINPUT107), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n364), .B1(new_n778), .B2(new_n202), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n773), .A2(new_n272), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n990), .B(new_n991), .C1(G159), .C2(new_n798), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n988), .A2(KEYINPUT107), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n782), .A2(new_n863), .B1(new_n403), .B2(new_n786), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT108), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n992), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n984), .B1(new_n989), .B2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT47), .Z(new_n998));
  OAI211_X1 g0798(.A(new_n758), .B(new_n974), .C1(new_n998), .C2(new_n766), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT109), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n589), .A2(new_n696), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n673), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n673), .A2(new_n593), .A3(new_n1001), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1000), .B1(new_n832), .B2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n715), .B(KEYINPUT41), .Z(new_n1006));
  INV_X1    g0806(.A(new_n482), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT102), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1007), .A2(new_n1008), .A3(new_n696), .ZN(new_n1009));
  OAI21_X1  g0809(.A(KEYINPUT102), .B1(new_n482), .B2(new_n697), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n482), .A2(new_n500), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n458), .A2(new_n696), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n1009), .A2(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n711), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT45), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n711), .A2(new_n1013), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT44), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n709), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n700), .A2(new_n697), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n707), .A2(new_n1022), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1023), .A2(new_n710), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n754), .A2(new_n1024), .ZN(new_n1025));
  OR3_X1    g0825(.A1(new_n760), .A2(new_n1024), .A3(new_n728), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1015), .A2(new_n709), .A3(new_n1018), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1021), .A2(new_n752), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1006), .B1(new_n1029), .B2(new_n752), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1030), .A2(new_n757), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1013), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1007), .B1(new_n1032), .B2(new_n703), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1033), .A2(new_n696), .ZN(new_n1034));
  OR3_X1    g0834(.A1(new_n1013), .A2(KEYINPUT42), .A3(new_n710), .ZN(new_n1035));
  OAI21_X1  g0835(.A(KEYINPUT42), .B1(new_n1013), .B2(new_n710), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1004), .A2(KEYINPUT43), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1004), .A2(KEYINPUT43), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1038), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n709), .A2(new_n1013), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT43), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1004), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1034), .A2(new_n1037), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1042), .A2(new_n1043), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT103), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1043), .B1(new_n1042), .B2(new_n1046), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1042), .A2(KEYINPUT103), .A3(new_n1043), .A4(new_n1046), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1049), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1005), .B1(new_n1031), .B2(new_n1053), .ZN(G387));
  AOI21_X1  g0854(.A(new_n410), .B1(new_n783), .B2(G326), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n869), .A2(new_n774), .B1(new_n856), .B2(new_n786), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n860), .A2(G303), .B1(new_n861), .B2(G317), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n775), .B2(new_n797), .C1(new_n789), .C2(new_n791), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT48), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n1059), .B2(new_n1058), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT49), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1055), .B1(new_n528), .B2(new_n773), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n786), .A2(new_n272), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n398), .B(new_n1066), .C1(new_n861), .C2(G50), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n975), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n778), .A2(new_n335), .B1(new_n864), .B2(new_n782), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n869), .A2(new_n360), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n243), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n809), .A2(new_n791), .B1(new_n797), .B2(new_n1071), .ZN(new_n1072));
  NOR4_X1   g0872(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n765), .B1(new_n1065), .B2(new_n1073), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n230), .A2(new_n279), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1075), .A2(new_n824), .B1(new_n718), .B2(new_n821), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n357), .A2(G50), .ZN(new_n1077));
  XOR2_X1   g0877(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1078));
  XNOR2_X1  g0878(.A(new_n1077), .B(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n279), .B1(new_n335), .B2(new_n272), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n1079), .A2(new_n718), .A3(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n1076), .A2(new_n1081), .B1(G107), .B2(new_n207), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n759), .B1(new_n1082), .B2(new_n830), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1074), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n707), .B2(new_n829), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n1027), .B2(new_n757), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1027), .A2(new_n752), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1087), .A2(KEYINPUT111), .A3(new_n715), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n752), .B2(new_n1027), .ZN(new_n1089));
  AOI21_X1  g0889(.A(KEYINPUT111), .B1(new_n1087), .B2(new_n715), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1086), .B1(new_n1089), .B2(new_n1090), .ZN(G393));
  NAND2_X1  g0891(.A1(new_n1021), .A2(new_n1028), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n1087), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1093), .A2(new_n715), .A3(new_n1029), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n240), .A2(new_n824), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1095), .B(new_n830), .C1(new_n446), .C2(new_n207), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n869), .A2(new_n272), .B1(new_n797), .B2(new_n202), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n860), .A2(new_n358), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n398), .B1(new_n854), .B2(G68), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n783), .A2(G143), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n852), .A2(new_n1098), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n792), .A2(G150), .B1(G159), .B2(new_n861), .ZN(new_n1102));
  XOR2_X1   g0902(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n1103));
  AOI211_X1 g0903(.A(new_n1097), .B(new_n1101), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n791), .A2(new_n800), .B1(new_n775), .B2(new_n788), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT52), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n798), .A2(G303), .B1(G116), .B2(new_n795), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n364), .B1(G283), .B2(new_n854), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n860), .A2(G294), .B1(G322), .B2(new_n783), .ZN(new_n1110));
  AND4_X1   g0910(.A1(new_n804), .A2(new_n1108), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1104), .A2(new_n1105), .B1(new_n1107), .B2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n758), .B(new_n1096), .C1(new_n1112), .C2(new_n766), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n1013), .B2(new_n829), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1092), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1114), .B1(new_n1115), .B2(new_n757), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1094), .A2(new_n1116), .ZN(G390));
  AOI21_X1  g0917(.A(new_n950), .B1(new_n845), .B2(new_n948), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1118), .A2(new_n961), .B1(new_n958), .B2(new_n960), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n957), .A2(new_n938), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n724), .A2(new_n725), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n696), .B1(new_n1121), .B2(new_n687), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n947), .B1(new_n1122), .B2(new_n844), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n962), .B(new_n1120), .C1(new_n1123), .C2(new_n950), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n925), .A2(new_n928), .A3(new_n728), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(KEYINPUT113), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n751), .A2(new_n844), .A3(new_n951), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1119), .B(new_n1124), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1119), .A2(new_n1124), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT113), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1125), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1129), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n443), .A2(G330), .A3(new_n916), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n965), .A2(new_n670), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n951), .B1(new_n751), .B2(new_n844), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n949), .B1(new_n1136), .B2(new_n1125), .ZN(new_n1137));
  NOR3_X1   g0937(.A1(new_n925), .A2(new_n728), .A3(new_n840), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1128), .B(new_n1123), .C1(new_n1138), .C2(new_n951), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1135), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1133), .A2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1129), .B(new_n1140), .C1(new_n1130), .C2(new_n1132), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n715), .A3(new_n1143), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1133), .A2(new_n756), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n850), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n783), .A2(G125), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n364), .B(new_n1147), .C1(new_n773), .C2(new_n202), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT114), .Z(new_n1149));
  OAI22_X1  g0949(.A1(new_n869), .A2(new_n809), .B1(new_n797), .B2(new_n863), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n786), .A2(new_n864), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT53), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT54), .B(G143), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1152), .B1(new_n788), .B2(new_n870), .C1(new_n778), .C2(new_n1153), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1150), .B(new_n1154), .C1(G128), .C2(new_n792), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n773), .A2(new_n335), .B1(new_n856), .B2(new_n782), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(G97), .B2(new_n860), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n271), .B1(new_n518), .B2(new_n786), .C1(new_n788), .C2(new_n528), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n496), .A2(new_n797), .B1(new_n791), .B2(new_n774), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1158), .B(new_n1159), .C1(G77), .C2(new_n795), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1149), .A2(new_n1155), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n758), .B1(new_n243), .B2(new_n1146), .C1(new_n1161), .C2(new_n766), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n959), .B1(new_n912), .B2(KEYINPUT39), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1162), .B1(new_n1163), .B2(new_n827), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1144), .A2(new_n1145), .A3(new_n1165), .ZN(G378));
  OR2_X1    g0966(.A1(new_n954), .A2(new_n963), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n259), .A2(new_n694), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT55), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n302), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n302), .A2(new_n1170), .ZN(new_n1172));
  XOR2_X1   g0972(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  OR3_X1    g0974(.A1(new_n1171), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1174), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n941), .B2(G330), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n930), .B1(new_n929), .B2(new_n1120), .ZN(new_n1179));
  AOI21_X1  g0979(.A(KEYINPUT38), .B1(new_n936), .B2(new_n937), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n930), .B1(new_n901), .B2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1181), .A2(new_n922), .ZN(new_n1182));
  OAI211_X1 g0982(.A(G330), .B(new_n1177), .C1(new_n1179), .C2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1167), .B1(new_n1178), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(G330), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1177), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1188), .A2(new_n964), .A3(new_n1183), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1185), .A2(KEYINPUT119), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1135), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1143), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT119), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1193), .B(new_n1167), .C1(new_n1178), .C2(new_n1184), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1190), .A2(new_n1192), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT57), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1196), .B1(new_n1143), .B2(new_n1191), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1185), .A2(new_n1189), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n716), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1190), .A2(new_n757), .A3(new_n1194), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1187), .A2(new_n827), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n758), .B1(G50), .B2(new_n1146), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n398), .A2(new_n278), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1205), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n773), .A2(new_n403), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n565), .B2(new_n860), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n788), .A2(new_n496), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1208), .B1(KEYINPUT115), .B2(new_n1209), .C1(new_n774), .C2(new_n782), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1066), .B(new_n1205), .C1(new_n1209), .C2(KEYINPUT115), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G97), .A2(new_n798), .B1(new_n792), .B2(G116), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1211), .A2(new_n1212), .A3(new_n987), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1206), .B1(new_n1214), .B2(KEYINPUT58), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(KEYINPUT58), .B2(new_n1214), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n792), .A2(G125), .B1(new_n860), .B2(G137), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n870), .B2(new_n797), .C1(new_n864), .C2(new_n869), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1153), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n861), .A2(G128), .B1(new_n854), .B2(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT116), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1218), .A2(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT117), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n783), .A2(G124), .ZN(new_n1225));
  AOI211_X1 g1025(.A(G33), .B(G41), .C1(new_n772), .C2(G159), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1216), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1204), .B1(new_n1229), .B2(new_n765), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1203), .A2(new_n1230), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1202), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1201), .A2(new_n1232), .ZN(G375));
  AND2_X1   g1033(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1135), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1006), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n1141), .A3(new_n1236), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT120), .Z(new_n1238));
  INV_X1    g1038(.A(new_n1234), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n950), .A2(new_n827), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n758), .B1(G68), .B2(new_n1146), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n991), .B1(G107), .B2(new_n860), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n785), .B2(new_n782), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n271), .B1(new_n446), .B2(new_n786), .C1(new_n788), .C2(new_n774), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n528), .A2(new_n797), .B1(new_n791), .B2(new_n856), .ZN(new_n1245));
  NOR4_X1   g1045(.A1(new_n1243), .A2(new_n1070), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1246), .A2(KEYINPUT121), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(KEYINPUT121), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n410), .B1(new_n786), .B2(new_n809), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n1249), .B(new_n1207), .C1(G137), .C2(new_n861), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n860), .A2(G150), .B1(G128), .B2(new_n783), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n795), .A2(G50), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(G132), .A2(new_n792), .B1(new_n798), .B2(new_n1219), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .A4(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1247), .A2(new_n1248), .A3(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1241), .B1(new_n1255), .B2(new_n765), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1239), .A2(new_n757), .B1(new_n1240), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1238), .A2(new_n1257), .ZN(G381));
  INV_X1    g1058(.A(G396), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1259), .B(new_n1086), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1260));
  OR4_X1    g1060(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1260), .ZN(new_n1261));
  OR4_X1    g1061(.A1(G378), .A2(new_n1261), .A3(G375), .A4(G381), .ZN(G407));
  NAND2_X1  g1062(.A1(new_n695), .A2(G213), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1263), .B(KEYINPUT122), .ZN(new_n1264));
  OR3_X1    g1064(.A1(G375), .A2(G378), .A3(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(G407), .A2(G213), .A3(new_n1265), .ZN(G409));
  INV_X1    g1066(.A(KEYINPUT63), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1201), .A2(G378), .A3(new_n1232), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1199), .A2(new_n757), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1269), .A2(KEYINPUT123), .A3(new_n1231), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT123), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n756), .B1(new_n1185), .B2(new_n1189), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1231), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1271), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1190), .A2(new_n1192), .A3(new_n1236), .A4(new_n1194), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1270), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(G378), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1268), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT60), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1235), .B1(new_n1280), .B2(new_n1140), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1234), .A2(KEYINPUT60), .A3(new_n1135), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1281), .A2(new_n715), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1257), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1284), .A2(new_n849), .A3(new_n874), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1283), .A2(G384), .A3(new_n1257), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  AND4_X1   g1087(.A1(KEYINPUT124), .A2(new_n1279), .A3(new_n1263), .A4(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1263), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1289), .B1(new_n1268), .B2(new_n1278), .ZN(new_n1290));
  AOI21_X1  g1090(.A(KEYINPUT124), .B1(new_n1290), .B2(new_n1287), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1267), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1279), .A2(new_n1264), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(KEYINPUT63), .A3(new_n1287), .ZN(new_n1294));
  INV_X1    g1094(.A(G2897), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1264), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1263), .A2(new_n1295), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1297), .B1(new_n1287), .B2(new_n1298), .ZN(new_n1299));
  OR2_X1    g1099(.A1(new_n1290), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(G393), .A2(G396), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1260), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1050), .B1(new_n1048), .B2(new_n1047), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1303), .B(new_n1052), .C1(new_n1030), .C2(new_n757), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1304), .A2(new_n1005), .A3(G390), .ZN(new_n1305));
  INV_X1    g1105(.A(G390), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(G387), .A2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1302), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT125), .ZN(new_n1309));
  OR2_X1    g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1311));
  OR2_X1    g1111(.A1(new_n1305), .A2(KEYINPUT126), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1305), .A2(KEYINPUT126), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1312), .A2(new_n1302), .A3(new_n1307), .A4(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1310), .A2(new_n1311), .A3(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT61), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1292), .A2(new_n1294), .A3(new_n1300), .A4(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1316), .B1(new_n1293), .B2(new_n1299), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT62), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1320), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1293), .A2(KEYINPUT62), .A3(new_n1287), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1319), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  XNOR2_X1  g1123(.A(new_n1315), .B(KEYINPUT127), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1318), .B1(new_n1323), .B2(new_n1324), .ZN(G405));
  XNOR2_X1  g1125(.A(G375), .B(G378), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(new_n1326), .B(new_n1287), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(new_n1327), .B(new_n1324), .ZN(G402));
endmodule


