

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741;

  XNOR2_X1 U370 ( .A(G116), .B(G107), .ZN(n457) );
  XNOR2_X1 U371 ( .A(G122), .B(G104), .ZN(n444) );
  XNOR2_X1 U372 ( .A(n407), .B(n406), .ZN(n722) );
  OR2_X2 U373 ( .A1(n701), .A2(n686), .ZN(n499) );
  XNOR2_X2 U374 ( .A(n540), .B(n539), .ZN(n622) );
  XNOR2_X1 U375 ( .A(n545), .B(KEYINPUT41), .ZN(n674) );
  OR2_X2 U376 ( .A1(n535), .A2(n645), .ZN(n570) );
  XNOR2_X1 U377 ( .A(n382), .B(n381), .ZN(n473) );
  XNOR2_X2 U378 ( .A(n570), .B(KEYINPUT19), .ZN(n559) );
  XNOR2_X2 U379 ( .A(n357), .B(G110), .ZN(n402) );
  XNOR2_X1 U380 ( .A(n353), .B(G131), .ZN(n728) );
  INV_X1 U381 ( .A(n638), .ZN(n600) );
  NAND2_X1 U382 ( .A1(n597), .A2(n596), .ZN(n601) );
  OR2_X1 U383 ( .A1(n624), .A2(G902), .ZN(n382) );
  BUF_X1 U384 ( .A(n472), .Z(n652) );
  XNOR2_X1 U385 ( .A(n728), .B(n360), .ZN(n706) );
  XNOR2_X1 U386 ( .A(n359), .B(n351), .ZN(n360) );
  NOR2_X1 U387 ( .A1(n599), .A2(n598), .ZN(n638) );
  INV_X1 U388 ( .A(n532), .ZN(n489) );
  INV_X1 U389 ( .A(n563), .ZN(n463) );
  XNOR2_X1 U390 ( .A(n477), .B(KEYINPUT32), .ZN(n614) );
  XOR2_X1 U391 ( .A(n475), .B(KEYINPUT78), .Z(n347) );
  XOR2_X1 U392 ( .A(n603), .B(n602), .Z(n348) );
  XOR2_X1 U393 ( .A(n434), .B(KEYINPUT34), .Z(n349) );
  XOR2_X1 U394 ( .A(KEYINPUT84), .B(KEYINPUT48), .Z(n350) );
  XOR2_X1 U395 ( .A(n402), .B(n358), .Z(n351) );
  AND2_X1 U396 ( .A1(n542), .A2(n469), .ZN(n352) );
  INV_X1 U397 ( .A(KEYINPUT75), .ZN(n388) );
  INV_X1 U398 ( .A(KEYINPUT76), .ZN(n357) );
  XNOR2_X1 U399 ( .A(n389), .B(n388), .ZN(n390) );
  NOR2_X1 U400 ( .A1(G953), .A2(G237), .ZN(n436) );
  XNOR2_X1 U401 ( .A(n391), .B(n390), .ZN(n396) );
  XNOR2_X1 U402 ( .A(G143), .B(G128), .ZN(n454) );
  XNOR2_X1 U403 ( .A(n356), .B(n727), .ZN(n359) );
  AND2_X1 U404 ( .A1(n658), .A2(n657), .ZN(n651) );
  NAND2_X1 U405 ( .A1(n651), .A2(n488), .ZN(n532) );
  XNOR2_X1 U406 ( .A(G140), .B(G137), .ZN(n727) );
  AND2_X1 U407 ( .A1(n472), .A2(n651), .ZN(n485) );
  AND2_X2 U408 ( .A1(n601), .A2(n600), .ZN(n627) );
  BUF_X1 U409 ( .A(n634), .Z(n732) );
  BUF_X1 U410 ( .A(n627), .Z(n712) );
  XNOR2_X1 U411 ( .A(n488), .B(KEYINPUT1), .ZN(n472) );
  INV_X1 U412 ( .A(n716), .ZN(n606) );
  OR2_X1 U413 ( .A1(n592), .A2(n694), .ZN(n540) );
  NAND2_X1 U414 ( .A1(n505), .A2(n504), .ZN(n613) );
  XNOR2_X1 U415 ( .A(n454), .B(KEYINPUT4), .ZN(n413) );
  XNOR2_X1 U416 ( .A(n413), .B(G134), .ZN(n353) );
  XOR2_X1 U417 ( .A(G107), .B(G104), .Z(n355) );
  XNOR2_X1 U418 ( .A(G101), .B(G146), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n355), .B(n354), .ZN(n356) );
  INV_X2 U420 ( .A(G953), .ZN(n733) );
  NAND2_X1 U421 ( .A1(G227), .A2(n733), .ZN(n358) );
  NOR2_X1 U422 ( .A1(n706), .A2(G902), .ZN(n363) );
  INV_X1 U423 ( .A(KEYINPUT68), .ZN(n361) );
  XNOR2_X1 U424 ( .A(n361), .B(G469), .ZN(n362) );
  XNOR2_X2 U425 ( .A(n363), .B(n362), .ZN(n488) );
  XNOR2_X1 U426 ( .A(G110), .B(G128), .ZN(n365) );
  XNOR2_X1 U427 ( .A(G119), .B(KEYINPUT23), .ZN(n364) );
  XNOR2_X1 U428 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n366), .B(n727), .ZN(n370) );
  NAND2_X1 U430 ( .A1(n733), .A2(G234), .ZN(n368) );
  XNOR2_X1 U431 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n368), .B(n367), .ZN(n451) );
  NAND2_X1 U433 ( .A1(n451), .A2(G221), .ZN(n369) );
  XNOR2_X1 U434 ( .A(n370), .B(n369), .ZN(n375) );
  XNOR2_X1 U435 ( .A(G146), .B(G125), .ZN(n409) );
  XNOR2_X1 U436 ( .A(n409), .B(KEYINPUT10), .ZN(n729) );
  XNOR2_X1 U437 ( .A(KEYINPUT24), .B(KEYINPUT77), .ZN(n372) );
  XNOR2_X1 U438 ( .A(KEYINPUT79), .B(KEYINPUT92), .ZN(n371) );
  XNOR2_X1 U439 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U440 ( .A(n729), .B(n373), .ZN(n374) );
  XNOR2_X1 U441 ( .A(n375), .B(n374), .ZN(n624) );
  XNOR2_X1 U442 ( .A(G902), .B(KEYINPUT15), .ZN(n523) );
  NAND2_X1 U443 ( .A1(n523), .A2(G234), .ZN(n376) );
  XNOR2_X1 U444 ( .A(n376), .B(KEYINPUT20), .ZN(n383) );
  NAND2_X1 U445 ( .A1(n383), .A2(G217), .ZN(n380) );
  XNOR2_X1 U446 ( .A(KEYINPUT93), .B(KEYINPUT94), .ZN(n378) );
  INV_X1 U447 ( .A(KEYINPUT25), .ZN(n377) );
  XNOR2_X1 U448 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U449 ( .A(n380), .B(n379), .ZN(n381) );
  INV_X1 U450 ( .A(n473), .ZN(n658) );
  NAND2_X1 U451 ( .A1(n383), .A2(G221), .ZN(n385) );
  XNOR2_X1 U452 ( .A(KEYINPUT95), .B(KEYINPUT21), .ZN(n384) );
  XNOR2_X1 U453 ( .A(n385), .B(n384), .ZN(n657) );
  XOR2_X1 U454 ( .A(G146), .B(KEYINPUT5), .Z(n387) );
  NAND2_X1 U455 ( .A1(n436), .A2(G210), .ZN(n386) );
  XNOR2_X1 U456 ( .A(n387), .B(n386), .ZN(n391) );
  XNOR2_X1 U457 ( .A(G137), .B(G116), .ZN(n389) );
  XNOR2_X1 U458 ( .A(G119), .B(G113), .ZN(n392) );
  XNOR2_X1 U459 ( .A(n392), .B(KEYINPUT3), .ZN(n395) );
  INV_X1 U460 ( .A(KEYINPUT69), .ZN(n393) );
  XNOR2_X1 U461 ( .A(n393), .B(G101), .ZN(n394) );
  XNOR2_X1 U462 ( .A(n395), .B(n394), .ZN(n406) );
  XNOR2_X1 U463 ( .A(n396), .B(n406), .ZN(n397) );
  XNOR2_X1 U464 ( .A(n728), .B(n397), .ZN(n603) );
  INV_X1 U465 ( .A(G902), .ZN(n417) );
  NAND2_X1 U466 ( .A1(n603), .A2(n417), .ZN(n398) );
  XNOR2_X2 U467 ( .A(n398), .B(G472), .ZN(n525) );
  INV_X1 U468 ( .A(KEYINPUT6), .ZN(n399) );
  XNOR2_X1 U469 ( .A(n525), .B(n399), .ZN(n568) );
  NAND2_X1 U470 ( .A1(n485), .A2(n568), .ZN(n401) );
  INV_X1 U471 ( .A(KEYINPUT33), .ZN(n400) );
  XNOR2_X1 U472 ( .A(n401), .B(n400), .ZN(n673) );
  INV_X1 U473 ( .A(n673), .ZN(n433) );
  XNOR2_X1 U474 ( .A(n402), .B(n444), .ZN(n405) );
  XNOR2_X1 U475 ( .A(KEYINPUT73), .B(KEYINPUT16), .ZN(n403) );
  XNOR2_X1 U476 ( .A(n457), .B(n403), .ZN(n404) );
  XNOR2_X1 U477 ( .A(n405), .B(n404), .ZN(n407) );
  XNOR2_X1 U478 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n408) );
  XNOR2_X1 U479 ( .A(n409), .B(n408), .ZN(n412) );
  NAND2_X1 U480 ( .A1(n733), .A2(G224), .ZN(n410) );
  XNOR2_X1 U481 ( .A(n410), .B(KEYINPUT88), .ZN(n411) );
  XNOR2_X1 U482 ( .A(n412), .B(n411), .ZN(n414) );
  XNOR2_X1 U483 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U484 ( .A(n722), .B(n415), .ZN(n616) );
  INV_X1 U485 ( .A(n523), .ZN(n595) );
  OR2_X2 U486 ( .A1(n616), .A2(n595), .ZN(n419) );
  INV_X1 U487 ( .A(G237), .ZN(n416) );
  NAND2_X1 U488 ( .A1(n417), .A2(n416), .ZN(n420) );
  NAND2_X1 U489 ( .A1(n420), .A2(G210), .ZN(n418) );
  XNOR2_X2 U490 ( .A(n419), .B(n418), .ZN(n535) );
  NAND2_X1 U491 ( .A1(n420), .A2(G214), .ZN(n421) );
  XNOR2_X1 U492 ( .A(n421), .B(KEYINPUT89), .ZN(n645) );
  XOR2_X1 U493 ( .A(KEYINPUT90), .B(KEYINPUT14), .Z(n423) );
  NAND2_X1 U494 ( .A1(G234), .A2(G237), .ZN(n422) );
  XNOR2_X1 U495 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U496 ( .A(KEYINPUT74), .B(n424), .Z(n426) );
  AND2_X1 U497 ( .A1(G953), .A2(n426), .ZN(n425) );
  NAND2_X1 U498 ( .A1(G902), .A2(n425), .ZN(n527) );
  NOR2_X1 U499 ( .A1(G898), .A2(n527), .ZN(n427) );
  NAND2_X1 U500 ( .A1(G952), .A2(n426), .ZN(n671) );
  NOR2_X1 U501 ( .A1(G953), .A2(n671), .ZN(n528) );
  OR2_X1 U502 ( .A1(n427), .A2(n528), .ZN(n429) );
  INV_X1 U503 ( .A(KEYINPUT91), .ZN(n428) );
  XNOR2_X1 U504 ( .A(n429), .B(n428), .ZN(n430) );
  NAND2_X1 U505 ( .A1(n559), .A2(n430), .ZN(n432) );
  INV_X1 U506 ( .A(KEYINPUT0), .ZN(n431) );
  XNOR2_X2 U507 ( .A(n432), .B(n431), .ZN(n490) );
  NAND2_X1 U508 ( .A1(n433), .A2(n490), .ZN(n435) );
  INV_X1 U509 ( .A(KEYINPUT71), .ZN(n434) );
  XNOR2_X1 U510 ( .A(n435), .B(n349), .ZN(n464) );
  XNOR2_X1 U511 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n449) );
  XOR2_X1 U512 ( .A(G131), .B(KEYINPUT12), .Z(n438) );
  NAND2_X1 U513 ( .A1(G214), .A2(n436), .ZN(n437) );
  XNOR2_X1 U514 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U515 ( .A(KEYINPUT11), .B(KEYINPUT97), .Z(n440) );
  XNOR2_X1 U516 ( .A(G140), .B(KEYINPUT98), .ZN(n439) );
  XNOR2_X1 U517 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U518 ( .A(n442), .B(n441), .ZN(n447) );
  XNOR2_X1 U519 ( .A(G113), .B(G143), .ZN(n443) );
  XNOR2_X1 U520 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U521 ( .A(n729), .B(n445), .ZN(n446) );
  XNOR2_X1 U522 ( .A(n447), .B(n446), .ZN(n629) );
  NOR2_X1 U523 ( .A1(G902), .A2(n629), .ZN(n448) );
  XNOR2_X1 U524 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U525 ( .A(n450), .B(G475), .ZN(n542) );
  XNOR2_X1 U526 ( .A(KEYINPUT101), .B(G478), .ZN(n461) );
  XOR2_X1 U527 ( .A(G122), .B(KEYINPUT9), .Z(n453) );
  NAND2_X1 U528 ( .A1(G217), .A2(n451), .ZN(n452) );
  XNOR2_X1 U529 ( .A(n453), .B(n452), .ZN(n459) );
  XOR2_X1 U530 ( .A(KEYINPUT7), .B(G134), .Z(n455) );
  XNOR2_X1 U531 ( .A(n454), .B(n455), .ZN(n456) );
  XNOR2_X1 U532 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U533 ( .A(n459), .B(n458), .ZN(n713) );
  NOR2_X1 U534 ( .A1(G902), .A2(n713), .ZN(n460) );
  XNOR2_X1 U535 ( .A(n461), .B(n460), .ZN(n497) );
  INV_X1 U536 ( .A(n497), .ZN(n541) );
  OR2_X1 U537 ( .A1(n542), .A2(n541), .ZN(n462) );
  XNOR2_X1 U538 ( .A(n462), .B(KEYINPUT104), .ZN(n563) );
  NAND2_X1 U539 ( .A1(n464), .A2(n463), .ZN(n466) );
  INV_X1 U540 ( .A(KEYINPUT35), .ZN(n465) );
  XNOR2_X2 U541 ( .A(n466), .B(n465), .ZN(n623) );
  NOR2_X1 U542 ( .A1(KEYINPUT44), .A2(KEYINPUT87), .ZN(n467) );
  NAND2_X1 U543 ( .A1(n623), .A2(n467), .ZN(n468) );
  NAND2_X1 U544 ( .A1(n468), .A2(KEYINPUT66), .ZN(n481) );
  AND2_X1 U545 ( .A1(n657), .A2(n541), .ZN(n469) );
  NAND2_X1 U546 ( .A1(n490), .A2(n352), .ZN(n471) );
  XNOR2_X1 U547 ( .A(KEYINPUT72), .B(KEYINPUT22), .ZN(n470) );
  XNOR2_X1 U548 ( .A(n471), .B(n470), .ZN(n500) );
  INV_X1 U549 ( .A(n500), .ZN(n476) );
  NAND2_X1 U550 ( .A1(n652), .A2(n473), .ZN(n474) );
  OR2_X1 U551 ( .A1(n474), .A2(n568), .ZN(n475) );
  NAND2_X1 U552 ( .A1(n476), .A2(n347), .ZN(n477) );
  INV_X1 U553 ( .A(n525), .ZN(n493) );
  INV_X1 U554 ( .A(n493), .ZN(n656) );
  OR2_X1 U555 ( .A1(n656), .A2(n658), .ZN(n478) );
  OR2_X1 U556 ( .A1(n652), .A2(n478), .ZN(n479) );
  OR2_X1 U557 ( .A1(n500), .A2(n479), .ZN(n612) );
  NAND2_X1 U558 ( .A1(n614), .A2(n612), .ZN(n513) );
  INV_X1 U559 ( .A(n513), .ZN(n480) );
  NAND2_X1 U560 ( .A1(n481), .A2(n480), .ZN(n484) );
  INV_X1 U561 ( .A(n623), .ZN(n482) );
  NAND2_X1 U562 ( .A1(n482), .A2(KEYINPUT44), .ZN(n483) );
  NAND2_X1 U563 ( .A1(n484), .A2(n483), .ZN(n510) );
  NAND2_X1 U564 ( .A1(n485), .A2(n656), .ZN(n663) );
  INV_X1 U565 ( .A(n490), .ZN(n486) );
  OR2_X2 U566 ( .A1(n663), .A2(n486), .ZN(n487) );
  XNOR2_X2 U567 ( .A(n487), .B(KEYINPUT31), .ZN(n701) );
  NAND2_X1 U568 ( .A1(n490), .A2(n489), .ZN(n492) );
  INV_X1 U569 ( .A(KEYINPUT96), .ZN(n491) );
  XNOR2_X1 U570 ( .A(n492), .B(n491), .ZN(n494) );
  AND2_X1 U571 ( .A1(n494), .A2(n493), .ZN(n686) );
  XNOR2_X1 U572 ( .A(n542), .B(KEYINPUT100), .ZN(n498) );
  NAND2_X1 U573 ( .A1(n498), .A2(n497), .ZN(n496) );
  INV_X1 U574 ( .A(KEYINPUT102), .ZN(n495) );
  XNOR2_X1 U575 ( .A(n496), .B(n495), .ZN(n700) );
  OR2_X1 U576 ( .A1(n498), .A2(n497), .ZN(n694) );
  INV_X1 U577 ( .A(n694), .ZN(n697) );
  OR2_X1 U578 ( .A1(n700), .A2(n697), .ZN(n640) );
  NAND2_X1 U579 ( .A1(n499), .A2(n640), .ZN(n506) );
  INV_X1 U580 ( .A(n568), .ZN(n501) );
  NAND2_X1 U581 ( .A1(n476), .A2(n501), .ZN(n503) );
  INV_X1 U582 ( .A(KEYINPUT86), .ZN(n502) );
  XNOR2_X1 U583 ( .A(n503), .B(n502), .ZN(n505) );
  NOR2_X1 U584 ( .A1(n652), .A2(n473), .ZN(n504) );
  NAND2_X1 U585 ( .A1(n506), .A2(n613), .ZN(n508) );
  INV_X1 U586 ( .A(KEYINPUT103), .ZN(n507) );
  XNOR2_X1 U587 ( .A(n508), .B(n507), .ZN(n509) );
  NOR2_X1 U588 ( .A1(n510), .A2(n509), .ZN(n520) );
  NAND2_X1 U589 ( .A1(n623), .A2(KEYINPUT87), .ZN(n512) );
  INV_X1 U590 ( .A(KEYINPUT44), .ZN(n511) );
  NAND2_X1 U591 ( .A1(n512), .A2(n511), .ZN(n514) );
  NAND2_X1 U592 ( .A1(n514), .A2(n513), .ZN(n515) );
  NAND2_X1 U593 ( .A1(n515), .A2(KEYINPUT66), .ZN(n518) );
  INV_X1 U594 ( .A(KEYINPUT66), .ZN(n516) );
  NAND2_X1 U595 ( .A1(n516), .A2(KEYINPUT44), .ZN(n517) );
  NAND2_X1 U596 ( .A1(n518), .A2(n517), .ZN(n519) );
  NAND2_X1 U597 ( .A1(n520), .A2(n519), .ZN(n522) );
  XNOR2_X1 U598 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n521) );
  XNOR2_X2 U599 ( .A(n522), .B(n521), .ZN(n635) );
  NOR2_X2 U600 ( .A1(n635), .A2(n523), .ZN(n524) );
  XNOR2_X1 U601 ( .A(n524), .B(KEYINPUT80), .ZN(n594) );
  INV_X1 U602 ( .A(n645), .ZN(n544) );
  AND2_X1 U603 ( .A1(n525), .A2(n544), .ZN(n526) );
  XNOR2_X1 U604 ( .A(n526), .B(KEYINPUT30), .ZN(n530) );
  NOR2_X1 U605 ( .A1(G900), .A2(n527), .ZN(n529) );
  OR2_X1 U606 ( .A1(n529), .A2(n528), .ZN(n546) );
  AND2_X1 U607 ( .A1(n530), .A2(n546), .ZN(n534) );
  INV_X1 U608 ( .A(KEYINPUT108), .ZN(n531) );
  XNOR2_X1 U609 ( .A(n532), .B(n531), .ZN(n533) );
  NAND2_X1 U610 ( .A1(n534), .A2(n533), .ZN(n562) );
  BUF_X2 U611 ( .A(n535), .Z(n585) );
  INV_X1 U612 ( .A(n585), .ZN(n536) );
  XNOR2_X1 U613 ( .A(n536), .B(KEYINPUT38), .ZN(n641) );
  NOR2_X1 U614 ( .A1(n562), .A2(n641), .ZN(n538) );
  XNOR2_X1 U615 ( .A(KEYINPUT70), .B(KEYINPUT39), .ZN(n537) );
  XNOR2_X1 U616 ( .A(n538), .B(n537), .ZN(n592) );
  XNOR2_X1 U617 ( .A(KEYINPUT110), .B(KEYINPUT40), .ZN(n539) );
  AND2_X1 U618 ( .A1(n542), .A2(n541), .ZN(n643) );
  INV_X1 U619 ( .A(n641), .ZN(n543) );
  AND2_X1 U620 ( .A1(n643), .A2(n543), .ZN(n647) );
  NAND2_X1 U621 ( .A1(n647), .A2(n544), .ZN(n545) );
  AND2_X1 U622 ( .A1(n546), .A2(n657), .ZN(n547) );
  NAND2_X1 U623 ( .A1(n473), .A2(n547), .ZN(n567) );
  INV_X1 U624 ( .A(n567), .ZN(n548) );
  NAND2_X1 U625 ( .A1(n656), .A2(n548), .ZN(n550) );
  XNOR2_X1 U626 ( .A(KEYINPUT109), .B(KEYINPUT28), .ZN(n549) );
  XNOR2_X1 U627 ( .A(n550), .B(n549), .ZN(n551) );
  AND2_X1 U628 ( .A1(n488), .A2(n551), .ZN(n558) );
  NAND2_X1 U629 ( .A1(n674), .A2(n558), .ZN(n554) );
  INV_X1 U630 ( .A(KEYINPUT111), .ZN(n552) );
  XNOR2_X1 U631 ( .A(n552), .B(KEYINPUT42), .ZN(n553) );
  XNOR2_X1 U632 ( .A(n554), .B(n553), .ZN(n610) );
  NAND2_X1 U633 ( .A1(n622), .A2(n610), .ZN(n557) );
  XNOR2_X1 U634 ( .A(KEYINPUT85), .B(KEYINPUT46), .ZN(n555) );
  XNOR2_X1 U635 ( .A(n555), .B(KEYINPUT64), .ZN(n556) );
  XNOR2_X1 U636 ( .A(n557), .B(n556), .ZN(n578) );
  AND2_X1 U637 ( .A1(n559), .A2(n558), .ZN(n689) );
  NAND2_X1 U638 ( .A1(n640), .A2(n689), .ZN(n561) );
  INV_X1 U639 ( .A(KEYINPUT47), .ZN(n560) );
  XNOR2_X1 U640 ( .A(n561), .B(n560), .ZN(n566) );
  INV_X1 U641 ( .A(n562), .ZN(n565) );
  NOR2_X1 U642 ( .A1(n563), .A2(n585), .ZN(n564) );
  NAND2_X1 U643 ( .A1(n565), .A2(n564), .ZN(n609) );
  NAND2_X1 U644 ( .A1(n566), .A2(n609), .ZN(n576) );
  NOR2_X1 U645 ( .A1(n694), .A2(n567), .ZN(n569) );
  AND2_X1 U646 ( .A1(n569), .A2(n568), .ZN(n582) );
  INV_X1 U647 ( .A(n570), .ZN(n571) );
  NAND2_X1 U648 ( .A1(n582), .A2(n571), .ZN(n573) );
  INV_X1 U649 ( .A(KEYINPUT36), .ZN(n572) );
  XNOR2_X1 U650 ( .A(n573), .B(n572), .ZN(n574) );
  NAND2_X1 U651 ( .A1(n574), .A2(n652), .ZN(n705) );
  INV_X1 U652 ( .A(n705), .ZN(n575) );
  NOR2_X1 U653 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U654 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U655 ( .A(n579), .B(n350), .ZN(n589) );
  XNOR2_X1 U656 ( .A(KEYINPUT43), .B(KEYINPUT105), .ZN(n580) );
  XNOR2_X1 U657 ( .A(n580), .B(KEYINPUT106), .ZN(n584) );
  NOR2_X1 U658 ( .A1(n645), .A2(n652), .ZN(n581) );
  NAND2_X1 U659 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U660 ( .A(n584), .B(n583), .Z(n586) );
  NAND2_X1 U661 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U662 ( .A(n587), .B(KEYINPUT107), .ZN(n741) );
  INV_X1 U663 ( .A(n741), .ZN(n588) );
  NAND2_X1 U664 ( .A1(n589), .A2(n588), .ZN(n591) );
  INV_X1 U665 ( .A(KEYINPUT82), .ZN(n590) );
  XNOR2_X1 U666 ( .A(n591), .B(n590), .ZN(n593) );
  INV_X1 U667 ( .A(n700), .ZN(n690) );
  OR2_X1 U668 ( .A1(n592), .A2(n690), .ZN(n611) );
  NAND2_X2 U669 ( .A1(n593), .A2(n611), .ZN(n598) );
  XNOR2_X2 U670 ( .A(n598), .B(KEYINPUT81), .ZN(n634) );
  NAND2_X1 U671 ( .A1(n594), .A2(n634), .ZN(n597) );
  NAND2_X1 U672 ( .A1(n595), .A2(KEYINPUT2), .ZN(n596) );
  INV_X1 U673 ( .A(n635), .ZN(n717) );
  NAND2_X1 U674 ( .A1(n717), .A2(KEYINPUT2), .ZN(n599) );
  NAND2_X1 U675 ( .A1(n627), .A2(G472), .ZN(n604) );
  XOR2_X1 U676 ( .A(KEYINPUT112), .B(KEYINPUT62), .Z(n602) );
  XNOR2_X1 U677 ( .A(n604), .B(n348), .ZN(n607) );
  INV_X1 U678 ( .A(G952), .ZN(n605) );
  AND2_X1 U679 ( .A1(n605), .A2(G953), .ZN(n716) );
  NAND2_X1 U680 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U681 ( .A(n608), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U682 ( .A(n609), .B(G143), .ZN(G45) );
  XNOR2_X1 U683 ( .A(n610), .B(G137), .ZN(G39) );
  XNOR2_X1 U684 ( .A(n611), .B(G134), .ZN(G36) );
  XNOR2_X1 U685 ( .A(n612), .B(G110), .ZN(G12) );
  XNOR2_X1 U686 ( .A(n613), .B(G101), .ZN(G3) );
  XNOR2_X1 U687 ( .A(n614), .B(G119), .ZN(G21) );
  NAND2_X1 U688 ( .A1(n627), .A2(G210), .ZN(n618) );
  XOR2_X1 U689 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n615) );
  XNOR2_X1 U690 ( .A(n616), .B(n615), .ZN(n617) );
  XNOR2_X1 U691 ( .A(n618), .B(n617), .ZN(n619) );
  NOR2_X2 U692 ( .A1(n619), .A2(n716), .ZN(n621) );
  XOR2_X1 U693 ( .A(KEYINPUT83), .B(KEYINPUT56), .Z(n620) );
  XNOR2_X1 U694 ( .A(n621), .B(n620), .ZN(G51) );
  XNOR2_X1 U695 ( .A(n622), .B(G131), .ZN(G33) );
  XNOR2_X1 U696 ( .A(n623), .B(G122), .ZN(G24) );
  NAND2_X1 U697 ( .A1(n712), .A2(G217), .ZN(n625) );
  XNOR2_X1 U698 ( .A(n625), .B(n624), .ZN(n626) );
  NOR2_X1 U699 ( .A1(n626), .A2(n716), .ZN(G66) );
  NAND2_X1 U700 ( .A1(n627), .A2(G475), .ZN(n631) );
  XOR2_X1 U701 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n628) );
  XNOR2_X1 U702 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U703 ( .A(n631), .B(n630), .ZN(n632) );
  NOR2_X2 U704 ( .A1(n632), .A2(n716), .ZN(n633) );
  XNOR2_X1 U705 ( .A(n633), .B(KEYINPUT60), .ZN(G60) );
  INV_X1 U706 ( .A(n732), .ZN(n636) );
  NOR2_X1 U707 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U708 ( .A1(n637), .A2(KEYINPUT2), .ZN(n639) );
  OR2_X1 U709 ( .A1(n639), .A2(n638), .ZN(n679) );
  INV_X1 U710 ( .A(n640), .ZN(n642) );
  NOR2_X1 U711 ( .A1(n642), .A2(n641), .ZN(n644) );
  NOR2_X1 U712 ( .A1(n644), .A2(n643), .ZN(n646) );
  NOR2_X1 U713 ( .A1(n646), .A2(n645), .ZN(n648) );
  NOR2_X1 U714 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U715 ( .A(KEYINPUT121), .B(n649), .Z(n650) );
  NOR2_X1 U716 ( .A1(n650), .A2(n673), .ZN(n669) );
  NOR2_X1 U717 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U718 ( .A(KEYINPUT50), .B(n653), .Z(n654) );
  XNOR2_X1 U719 ( .A(KEYINPUT119), .B(n654), .ZN(n655) );
  NOR2_X1 U720 ( .A1(n656), .A2(n655), .ZN(n662) );
  XOR2_X1 U721 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n660) );
  NOR2_X1 U722 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U723 ( .A(n660), .B(n659), .Z(n661) );
  NAND2_X1 U724 ( .A1(n662), .A2(n661), .ZN(n664) );
  NAND2_X1 U725 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U726 ( .A(KEYINPUT51), .B(n665), .Z(n666) );
  NAND2_X1 U727 ( .A1(n666), .A2(n674), .ZN(n667) );
  XOR2_X1 U728 ( .A(KEYINPUT120), .B(n667), .Z(n668) );
  NOR2_X1 U729 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U730 ( .A(n670), .B(KEYINPUT52), .ZN(n672) );
  NOR2_X1 U731 ( .A1(n672), .A2(n671), .ZN(n677) );
  NAND2_X1 U732 ( .A1(n433), .A2(n674), .ZN(n675) );
  NAND2_X1 U733 ( .A1(n675), .A2(n733), .ZN(n676) );
  NOR2_X1 U734 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U735 ( .A1(n679), .A2(n678), .ZN(n681) );
  XOR2_X1 U736 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n680) );
  XNOR2_X1 U737 ( .A(n681), .B(n680), .ZN(G75) );
  NAND2_X1 U738 ( .A1(n686), .A2(n697), .ZN(n682) );
  XNOR2_X1 U739 ( .A(n682), .B(G104), .ZN(G6) );
  XOR2_X1 U740 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n684) );
  XNOR2_X1 U741 ( .A(G107), .B(KEYINPUT26), .ZN(n683) );
  XNOR2_X1 U742 ( .A(n684), .B(n683), .ZN(n685) );
  XOR2_X1 U743 ( .A(KEYINPUT113), .B(n685), .Z(n688) );
  NAND2_X1 U744 ( .A1(n686), .A2(n700), .ZN(n687) );
  XNOR2_X1 U745 ( .A(n688), .B(n687), .ZN(G9) );
  INV_X1 U746 ( .A(n689), .ZN(n695) );
  NOR2_X1 U747 ( .A1(n690), .A2(n695), .ZN(n692) );
  XNOR2_X1 U748 ( .A(KEYINPUT29), .B(KEYINPUT115), .ZN(n691) );
  XNOR2_X1 U749 ( .A(n692), .B(n691), .ZN(n693) );
  XOR2_X1 U750 ( .A(G128), .B(n693), .Z(G30) );
  NOR2_X1 U751 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U752 ( .A(G146), .B(n696), .Z(G48) );
  NAND2_X1 U753 ( .A1(n701), .A2(n697), .ZN(n698) );
  XNOR2_X1 U754 ( .A(n698), .B(KEYINPUT116), .ZN(n699) );
  XNOR2_X1 U755 ( .A(G113), .B(n699), .ZN(G15) );
  XOR2_X1 U756 ( .A(G116), .B(KEYINPUT117), .Z(n703) );
  NAND2_X1 U757 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U758 ( .A(n703), .B(n702), .ZN(G18) );
  XOR2_X1 U759 ( .A(G125), .B(KEYINPUT37), .Z(n704) );
  XNOR2_X1 U760 ( .A(n705), .B(n704), .ZN(G27) );
  NAND2_X1 U761 ( .A1(n712), .A2(G469), .ZN(n710) );
  XNOR2_X1 U762 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n708) );
  XNOR2_X1 U763 ( .A(n706), .B(KEYINPUT57), .ZN(n707) );
  XNOR2_X1 U764 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X1 U765 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U766 ( .A1(n716), .A2(n711), .ZN(G54) );
  NAND2_X1 U767 ( .A1(n712), .A2(G478), .ZN(n714) );
  XNOR2_X1 U768 ( .A(n714), .B(n713), .ZN(n715) );
  NOR2_X1 U769 ( .A1(n716), .A2(n715), .ZN(G63) );
  NAND2_X1 U770 ( .A1(n717), .A2(n733), .ZN(n721) );
  NAND2_X1 U771 ( .A1(G953), .A2(G224), .ZN(n718) );
  XNOR2_X1 U772 ( .A(KEYINPUT61), .B(n718), .ZN(n719) );
  NAND2_X1 U773 ( .A1(n719), .A2(G898), .ZN(n720) );
  NAND2_X1 U774 ( .A1(n721), .A2(n720), .ZN(n726) );
  XOR2_X1 U775 ( .A(KEYINPUT125), .B(n722), .Z(n724) );
  NOR2_X1 U776 ( .A1(G898), .A2(n733), .ZN(n723) );
  NOR2_X1 U777 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U778 ( .A(n726), .B(n725), .ZN(G69) );
  XNOR2_X1 U779 ( .A(n728), .B(n727), .ZN(n731) );
  XOR2_X1 U780 ( .A(KEYINPUT126), .B(n729), .Z(n730) );
  XNOR2_X1 U781 ( .A(n731), .B(n730), .ZN(n735) );
  XOR2_X1 U782 ( .A(n732), .B(n735), .Z(n734) );
  NAND2_X1 U783 ( .A1(n734), .A2(n733), .ZN(n740) );
  XNOR2_X1 U784 ( .A(G227), .B(n735), .ZN(n736) );
  NAND2_X1 U785 ( .A1(n736), .A2(G900), .ZN(n737) );
  XOR2_X1 U786 ( .A(KEYINPUT127), .B(n737), .Z(n738) );
  NAND2_X1 U787 ( .A1(G953), .A2(n738), .ZN(n739) );
  NAND2_X1 U788 ( .A1(n740), .A2(n739), .ZN(G72) );
  XOR2_X1 U789 ( .A(G140), .B(n741), .Z(G42) );
endmodule

