

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U550 ( .A1(G8), .A2(n669), .ZN(n678) );
  NOR2_X1 U551 ( .A1(G2104), .A2(G2105), .ZN(n545) );
  INV_X1 U552 ( .A(KEYINPUT17), .ZN(n544) );
  INV_X1 U553 ( .A(G2104), .ZN(n543) );
  NOR2_X1 U554 ( .A1(n535), .A2(n532), .ZN(n531) );
  AND2_X1 U555 ( .A1(n722), .A2(n518), .ZN(n535) );
  OR2_X1 U556 ( .A1(n671), .A2(n693), .ZN(n672) );
  NOR2_X1 U557 ( .A1(G164), .A2(G1384), .ZN(n622) );
  NOR2_X1 U558 ( .A1(n553), .A2(n552), .ZN(G160) );
  BUF_X2 U559 ( .A(n554), .Z(n517) );
  BUF_X2 U560 ( .A(n906), .Z(n516) );
  XNOR2_X1 U561 ( .A(n545), .B(n544), .ZN(n906) );
  OR2_X2 U562 ( .A1(n725), .A2(n723), .ZN(n669) );
  NOR2_X1 U563 ( .A1(n669), .A2(n961), .ZN(n624) );
  INV_X1 U564 ( .A(G2078), .ZN(n521) );
  NAND2_X1 U565 ( .A1(n721), .A2(n518), .ZN(n534) );
  INV_X1 U566 ( .A(KEYINPUT100), .ZN(n710) );
  INV_X1 U567 ( .A(KEYINPUT29), .ZN(n659) );
  NAND2_X1 U568 ( .A1(n705), .A2(n540), .ZN(n539) );
  XNOR2_X1 U569 ( .A(n622), .B(n621), .ZN(n723) );
  XNOR2_X1 U570 ( .A(G164), .B(n521), .ZN(n1002) );
  NAND2_X1 U571 ( .A1(n534), .A2(n533), .ZN(n532) );
  NAND2_X1 U572 ( .A1(n757), .A2(n537), .ZN(n533) );
  OR2_X1 U573 ( .A1(n721), .A2(KEYINPUT101), .ZN(n530) );
  INV_X1 U574 ( .A(n1013), .ZN(n522) );
  AND2_X1 U575 ( .A1(n538), .A2(KEYINPUT101), .ZN(n518) );
  NOR2_X1 U576 ( .A1(n725), .A2(n723), .ZN(n662) );
  XOR2_X1 U577 ( .A(KEYINPUT66), .B(n548), .Z(n519) );
  AND2_X1 U578 ( .A1(n626), .A2(n625), .ZN(n520) );
  AND2_X1 U579 ( .A1(n560), .A2(n561), .ZN(G164) );
  INV_X1 U580 ( .A(n757), .ZN(n538) );
  INV_X1 U581 ( .A(KEYINPUT101), .ZN(n537) );
  XNOR2_X1 U582 ( .A(n984), .B(G164), .ZN(n893) );
  NAND2_X1 U583 ( .A1(n520), .A2(n522), .ZN(n524) );
  AND2_X1 U584 ( .A1(n1019), .A2(n522), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n525), .A2(n523), .ZN(n652) );
  NAND2_X1 U586 ( .A1(n524), .A2(n528), .ZN(n523) );
  NAND2_X1 U587 ( .A1(n526), .A2(n647), .ZN(n525) );
  NAND2_X1 U588 ( .A1(n527), .A2(n520), .ZN(n526) );
  INV_X1 U589 ( .A(n1019), .ZN(n528) );
  NAND2_X1 U590 ( .A1(n531), .A2(n529), .ZN(n536) );
  OR2_X1 U591 ( .A1(n722), .A2(n530), .ZN(n529) );
  NAND2_X1 U592 ( .A1(n536), .A2(n771), .ZN(n772) );
  NAND2_X1 U593 ( .A1(n539), .A2(n709), .ZN(n711) );
  AND2_X1 U594 ( .A1(n706), .A2(n704), .ZN(n540) );
  NOR2_X2 U595 ( .A1(G2105), .A2(n543), .ZN(n907) );
  XNOR2_X1 U596 ( .A(KEYINPUT91), .B(n719), .ZN(n541) );
  AND2_X1 U597 ( .A1(n911), .A2(G114), .ZN(n542) );
  INV_X1 U598 ( .A(KEYINPUT26), .ZN(n623) );
  XNOR2_X1 U599 ( .A(n660), .B(n659), .ZN(n666) );
  XNOR2_X1 U600 ( .A(KEYINPUT31), .B(KEYINPUT97), .ZN(n676) );
  XNOR2_X1 U601 ( .A(n703), .B(KEYINPUT99), .ZN(n705) );
  NAND2_X1 U602 ( .A1(n720), .A2(n541), .ZN(n721) );
  NAND2_X1 U603 ( .A1(G160), .A2(G40), .ZN(n725) );
  AND2_X1 U604 ( .A1(G2104), .A2(G2105), .ZN(n911) );
  NOR2_X1 U605 ( .A1(G651), .A2(n611), .ZN(n803) );
  NOR2_X1 U606 ( .A1(n557), .A2(n542), .ZN(n561) );
  NAND2_X1 U607 ( .A1(n911), .A2(G113), .ZN(n547) );
  NAND2_X1 U608 ( .A1(n906), .A2(G137), .ZN(n546) );
  NAND2_X1 U609 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U610 ( .A1(n543), .A2(G2105), .ZN(n549) );
  XNOR2_X1 U611 ( .A(n549), .B(KEYINPUT65), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n517), .A2(G125), .ZN(n550) );
  NAND2_X1 U613 ( .A1(n519), .A2(n550), .ZN(n553) );
  NAND2_X1 U614 ( .A1(G101), .A2(n907), .ZN(n551) );
  XNOR2_X1 U615 ( .A(KEYINPUT23), .B(n551), .ZN(n552) );
  NAND2_X1 U616 ( .A1(G126), .A2(n517), .ZN(n556) );
  NAND2_X1 U617 ( .A1(G102), .A2(n907), .ZN(n555) );
  NAND2_X1 U618 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U619 ( .A1(G138), .A2(n516), .ZN(n559) );
  INV_X1 U620 ( .A(KEYINPUT85), .ZN(n558) );
  XNOR2_X1 U621 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U622 ( .A(KEYINPUT2), .B(KEYINPUT80), .Z(n563) );
  XOR2_X1 U623 ( .A(KEYINPUT0), .B(G543), .Z(n611) );
  INV_X1 U624 ( .A(G651), .ZN(n564) );
  NOR2_X1 U625 ( .A1(n611), .A2(n564), .ZN(n807) );
  NAND2_X1 U626 ( .A1(G73), .A2(n807), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n563), .B(n562), .ZN(n569) );
  NOR2_X1 U628 ( .A1(G543), .A2(n564), .ZN(n565) );
  XOR2_X1 U629 ( .A(KEYINPUT1), .B(n565), .Z(n802) );
  NAND2_X1 U630 ( .A1(G61), .A2(n802), .ZN(n567) );
  NOR2_X1 U631 ( .A1(G651), .A2(G543), .ZN(n806) );
  NAND2_X1 U632 ( .A1(G86), .A2(n806), .ZN(n566) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n803), .A2(G48), .ZN(n570) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(G305) );
  NAND2_X1 U637 ( .A1(G53), .A2(n803), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT70), .B(n572), .Z(n577) );
  NAND2_X1 U639 ( .A1(G91), .A2(n806), .ZN(n574) );
  NAND2_X1 U640 ( .A1(G78), .A2(n807), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U642 ( .A(KEYINPUT69), .B(n575), .Z(n576) );
  NOR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n802), .A2(G65), .ZN(n578) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(G299) );
  NAND2_X1 U646 ( .A1(G64), .A2(n802), .ZN(n581) );
  NAND2_X1 U647 ( .A1(G52), .A2(n803), .ZN(n580) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n587) );
  NAND2_X1 U649 ( .A1(n806), .A2(G90), .ZN(n582) );
  XOR2_X1 U650 ( .A(KEYINPUT67), .B(n582), .Z(n584) );
  NAND2_X1 U651 ( .A1(n807), .A2(G77), .ZN(n583) );
  NAND2_X1 U652 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U653 ( .A(KEYINPUT9), .B(n585), .Z(n586) );
  NOR2_X1 U654 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U655 ( .A(KEYINPUT68), .B(n588), .Z(G301) );
  INV_X1 U656 ( .A(G301), .ZN(G171) );
  NAND2_X1 U657 ( .A1(n806), .A2(G89), .ZN(n589) );
  XNOR2_X1 U658 ( .A(n589), .B(KEYINPUT4), .ZN(n591) );
  NAND2_X1 U659 ( .A1(G76), .A2(n807), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U661 ( .A(n592), .B(KEYINPUT5), .ZN(n598) );
  XNOR2_X1 U662 ( .A(KEYINPUT6), .B(KEYINPUT73), .ZN(n596) );
  NAND2_X1 U663 ( .A1(G63), .A2(n802), .ZN(n594) );
  NAND2_X1 U664 ( .A1(G51), .A2(n803), .ZN(n593) );
  NAND2_X1 U665 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U666 ( .A(n596), .B(n595), .ZN(n597) );
  NAND2_X1 U667 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U668 ( .A(KEYINPUT7), .B(n599), .ZN(G168) );
  NAND2_X1 U669 ( .A1(n802), .A2(G62), .ZN(n602) );
  NAND2_X1 U670 ( .A1(G75), .A2(n807), .ZN(n600) );
  XOR2_X1 U671 ( .A(KEYINPUT81), .B(n600), .Z(n601) );
  NAND2_X1 U672 ( .A1(n602), .A2(n601), .ZN(n606) );
  NAND2_X1 U673 ( .A1(G88), .A2(n806), .ZN(n604) );
  NAND2_X1 U674 ( .A1(G50), .A2(n803), .ZN(n603) );
  NAND2_X1 U675 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U676 ( .A1(n606), .A2(n605), .ZN(G166) );
  INV_X1 U677 ( .A(G166), .ZN(G303) );
  XOR2_X1 U678 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U679 ( .A1(G49), .A2(n803), .ZN(n608) );
  NAND2_X1 U680 ( .A1(G74), .A2(G651), .ZN(n607) );
  NAND2_X1 U681 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U682 ( .A(KEYINPUT79), .B(n609), .Z(n610) );
  NOR2_X1 U683 ( .A1(n802), .A2(n610), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n611), .A2(G87), .ZN(n612) );
  NAND2_X1 U685 ( .A1(n613), .A2(n612), .ZN(G288) );
  NAND2_X1 U686 ( .A1(G85), .A2(n806), .ZN(n615) );
  NAND2_X1 U687 ( .A1(G72), .A2(n807), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U689 ( .A1(G60), .A2(n802), .ZN(n617) );
  NAND2_X1 U690 ( .A1(G47), .A2(n803), .ZN(n616) );
  NAND2_X1 U691 ( .A1(n617), .A2(n616), .ZN(n618) );
  OR2_X1 U692 ( .A1(n619), .A2(n618), .ZN(G290) );
  XNOR2_X1 U693 ( .A(G1981), .B(G305), .ZN(n1017) );
  INV_X1 U694 ( .A(KEYINPUT64), .ZN(n621) );
  INV_X1 U695 ( .A(G1996), .ZN(n961) );
  XNOR2_X1 U696 ( .A(n624), .B(n623), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n669), .A2(G1341), .ZN(n625) );
  XOR2_X1 U698 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n628) );
  NAND2_X1 U699 ( .A1(G56), .A2(n802), .ZN(n627) );
  XNOR2_X1 U700 ( .A(n628), .B(n627), .ZN(n634) );
  NAND2_X1 U701 ( .A1(n806), .A2(G81), .ZN(n629) );
  XNOR2_X1 U702 ( .A(n629), .B(KEYINPUT12), .ZN(n631) );
  NAND2_X1 U703 ( .A1(G68), .A2(n807), .ZN(n630) );
  NAND2_X1 U704 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U705 ( .A(KEYINPUT13), .B(n632), .Z(n633) );
  NOR2_X1 U706 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U707 ( .A1(n803), .A2(G43), .ZN(n635) );
  NAND2_X1 U708 ( .A1(n636), .A2(n635), .ZN(n1013) );
  NAND2_X1 U709 ( .A1(G66), .A2(n802), .ZN(n638) );
  NAND2_X1 U710 ( .A1(G92), .A2(n806), .ZN(n637) );
  NAND2_X1 U711 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U712 ( .A1(G79), .A2(n807), .ZN(n640) );
  NAND2_X1 U713 ( .A1(G54), .A2(n803), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U715 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U716 ( .A(KEYINPUT15), .B(n643), .Z(n1019) );
  INV_X1 U717 ( .A(G2067), .ZN(n963) );
  NOR2_X1 U718 ( .A1(n669), .A2(n963), .ZN(n644) );
  XNOR2_X1 U719 ( .A(n644), .B(KEYINPUT95), .ZN(n646) );
  NAND2_X1 U720 ( .A1(n669), .A2(G1348), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U722 ( .A1(n662), .A2(G2072), .ZN(n648) );
  XNOR2_X1 U723 ( .A(n648), .B(KEYINPUT27), .ZN(n650) );
  INV_X1 U724 ( .A(G1956), .ZN(n934) );
  NOR2_X1 U725 ( .A1(n934), .A2(n662), .ZN(n649) );
  NOR2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n653) );
  INV_X1 U727 ( .A(G299), .ZN(n815) );
  NAND2_X1 U728 ( .A1(n653), .A2(n815), .ZN(n651) );
  NAND2_X1 U729 ( .A1(n652), .A2(n651), .ZN(n658) );
  NOR2_X1 U730 ( .A1(n653), .A2(n815), .ZN(n656) );
  XNOR2_X1 U731 ( .A(KEYINPUT28), .B(KEYINPUT94), .ZN(n654) );
  XNOR2_X1 U732 ( .A(n654), .B(KEYINPUT93), .ZN(n655) );
  XNOR2_X1 U733 ( .A(n656), .B(n655), .ZN(n657) );
  NAND2_X1 U734 ( .A1(n658), .A2(n657), .ZN(n660) );
  NOR2_X1 U735 ( .A1(n662), .A2(G1961), .ZN(n661) );
  XOR2_X1 U736 ( .A(KEYINPUT92), .B(n661), .Z(n664) );
  XNOR2_X1 U737 ( .A(KEYINPUT25), .B(G2078), .ZN(n969) );
  NAND2_X1 U738 ( .A1(n662), .A2(n969), .ZN(n663) );
  NAND2_X1 U739 ( .A1(n664), .A2(n663), .ZN(n668) );
  NAND2_X1 U740 ( .A1(G171), .A2(n668), .ZN(n665) );
  NAND2_X1 U741 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U742 ( .A(n667), .B(KEYINPUT96), .ZN(n692) );
  NOR2_X1 U743 ( .A1(G171), .A2(n668), .ZN(n675) );
  NOR2_X1 U744 ( .A1(G1966), .A2(n678), .ZN(n694) );
  INV_X1 U745 ( .A(n694), .ZN(n670) );
  NAND2_X1 U746 ( .A1(n670), .A2(G8), .ZN(n671) );
  NOR2_X1 U747 ( .A1(G2084), .A2(n669), .ZN(n693) );
  XNOR2_X1 U748 ( .A(n672), .B(KEYINPUT30), .ZN(n673) );
  NOR2_X1 U749 ( .A1(G168), .A2(n673), .ZN(n674) );
  NOR2_X1 U750 ( .A1(n675), .A2(n674), .ZN(n677) );
  XNOR2_X1 U751 ( .A(n677), .B(n676), .ZN(n691) );
  INV_X1 U752 ( .A(G8), .ZN(n683) );
  NOR2_X1 U753 ( .A1(G1971), .A2(n678), .ZN(n680) );
  NOR2_X1 U754 ( .A1(G2090), .A2(n669), .ZN(n679) );
  NOR2_X1 U755 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U756 ( .A1(n681), .A2(G303), .ZN(n682) );
  OR2_X1 U757 ( .A1(n683), .A2(n682), .ZN(n685) );
  AND2_X1 U758 ( .A1(n691), .A2(n685), .ZN(n684) );
  NAND2_X1 U759 ( .A1(n692), .A2(n684), .ZN(n689) );
  INV_X1 U760 ( .A(n685), .ZN(n687) );
  AND2_X1 U761 ( .A1(G286), .A2(G8), .ZN(n686) );
  OR2_X1 U762 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U763 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U764 ( .A(n690), .B(KEYINPUT32), .ZN(n700) );
  NAND2_X1 U765 ( .A1(n692), .A2(n691), .ZN(n697) );
  AND2_X1 U766 ( .A1(G8), .A2(n693), .ZN(n695) );
  NOR2_X1 U767 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U768 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U769 ( .A(n698), .B(KEYINPUT98), .ZN(n699) );
  NAND2_X1 U770 ( .A1(n700), .A2(n699), .ZN(n713) );
  NOR2_X1 U771 ( .A1(G1976), .A2(G288), .ZN(n707) );
  NOR2_X1 U772 ( .A1(G1971), .A2(G303), .ZN(n701) );
  NOR2_X1 U773 ( .A1(n707), .A2(n701), .ZN(n1015) );
  NAND2_X1 U774 ( .A1(n713), .A2(n1015), .ZN(n702) );
  NAND2_X1 U775 ( .A1(G1976), .A2(G288), .ZN(n1026) );
  NAND2_X1 U776 ( .A1(n702), .A2(n1026), .ZN(n703) );
  INV_X1 U777 ( .A(KEYINPUT33), .ZN(n704) );
  INV_X1 U778 ( .A(n678), .ZN(n706) );
  NAND2_X1 U779 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U780 ( .A1(n708), .A2(KEYINPUT33), .ZN(n709) );
  XNOR2_X1 U781 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U782 ( .A1(n1017), .A2(n712), .ZN(n722) );
  NOR2_X1 U783 ( .A1(G2090), .A2(G303), .ZN(n714) );
  NAND2_X1 U784 ( .A1(G8), .A2(n714), .ZN(n715) );
  NAND2_X1 U785 ( .A1(n713), .A2(n715), .ZN(n716) );
  NAND2_X1 U786 ( .A1(n716), .A2(n678), .ZN(n720) );
  NOR2_X1 U787 ( .A1(G1981), .A2(G305), .ZN(n717) );
  XOR2_X1 U788 ( .A(n717), .B(KEYINPUT24), .Z(n718) );
  NOR2_X1 U789 ( .A1(n678), .A2(n718), .ZN(n719) );
  INV_X1 U790 ( .A(n723), .ZN(n724) );
  NOR2_X1 U791 ( .A1(n725), .A2(n724), .ZN(n770) );
  XNOR2_X1 U792 ( .A(n770), .B(KEYINPUT90), .ZN(n743) );
  NAND2_X1 U793 ( .A1(G131), .A2(n516), .ZN(n727) );
  NAND2_X1 U794 ( .A1(G107), .A2(n911), .ZN(n726) );
  NAND2_X1 U795 ( .A1(n727), .A2(n726), .ZN(n730) );
  NAND2_X1 U796 ( .A1(n907), .A2(G95), .ZN(n728) );
  XOR2_X1 U797 ( .A(KEYINPUT88), .B(n728), .Z(n729) );
  NOR2_X1 U798 ( .A1(n730), .A2(n729), .ZN(n732) );
  NAND2_X1 U799 ( .A1(n517), .A2(G119), .ZN(n731) );
  NAND2_X1 U800 ( .A1(n732), .A2(n731), .ZN(n888) );
  NAND2_X1 U801 ( .A1(G1991), .A2(n888), .ZN(n742) );
  NAND2_X1 U802 ( .A1(G105), .A2(n907), .ZN(n733) );
  XOR2_X1 U803 ( .A(KEYINPUT38), .B(n733), .Z(n738) );
  NAND2_X1 U804 ( .A1(G117), .A2(n911), .ZN(n735) );
  NAND2_X1 U805 ( .A1(G129), .A2(n517), .ZN(n734) );
  NAND2_X1 U806 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U807 ( .A(KEYINPUT89), .B(n736), .Z(n737) );
  NOR2_X1 U808 ( .A1(n738), .A2(n737), .ZN(n740) );
  NAND2_X1 U809 ( .A1(n516), .A2(G141), .ZN(n739) );
  NAND2_X1 U810 ( .A1(n740), .A2(n739), .ZN(n886) );
  NAND2_X1 U811 ( .A1(G1996), .A2(n886), .ZN(n741) );
  NAND2_X1 U812 ( .A1(n742), .A2(n741), .ZN(n987) );
  NAND2_X1 U813 ( .A1(n743), .A2(n987), .ZN(n758) );
  XNOR2_X1 U814 ( .A(G1986), .B(G290), .ZN(n1021) );
  NAND2_X1 U815 ( .A1(n1021), .A2(n770), .ZN(n744) );
  XNOR2_X1 U816 ( .A(n744), .B(KEYINPUT86), .ZN(n755) );
  XNOR2_X1 U817 ( .A(G2067), .B(KEYINPUT37), .ZN(n767) );
  NAND2_X1 U818 ( .A1(G140), .A2(n516), .ZN(n746) );
  NAND2_X1 U819 ( .A1(G104), .A2(n907), .ZN(n745) );
  NAND2_X1 U820 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U821 ( .A(KEYINPUT34), .B(n747), .ZN(n753) );
  NAND2_X1 U822 ( .A1(G116), .A2(n911), .ZN(n749) );
  NAND2_X1 U823 ( .A1(G128), .A2(n517), .ZN(n748) );
  NAND2_X1 U824 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U825 ( .A(KEYINPUT35), .B(n750), .ZN(n751) );
  XNOR2_X1 U826 ( .A(KEYINPUT87), .B(n751), .ZN(n752) );
  NOR2_X1 U827 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U828 ( .A(KEYINPUT36), .B(n754), .ZN(n885) );
  NOR2_X1 U829 ( .A1(n767), .A2(n885), .ZN(n991) );
  NAND2_X1 U830 ( .A1(n770), .A2(n991), .ZN(n765) );
  AND2_X1 U831 ( .A1(n755), .A2(n765), .ZN(n756) );
  NAND2_X1 U832 ( .A1(n758), .A2(n756), .ZN(n757) );
  NOR2_X1 U833 ( .A1(G1996), .A2(n886), .ZN(n994) );
  INV_X1 U834 ( .A(n758), .ZN(n762) );
  NOR2_X1 U835 ( .A1(G1986), .A2(G290), .ZN(n759) );
  XNOR2_X1 U836 ( .A(n759), .B(KEYINPUT102), .ZN(n760) );
  NOR2_X1 U837 ( .A1(G1991), .A2(n888), .ZN(n985) );
  NOR2_X1 U838 ( .A1(n760), .A2(n985), .ZN(n761) );
  NOR2_X1 U839 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U840 ( .A1(n994), .A2(n763), .ZN(n764) );
  XNOR2_X1 U841 ( .A(n764), .B(KEYINPUT39), .ZN(n766) );
  NAND2_X1 U842 ( .A1(n766), .A2(n765), .ZN(n768) );
  NAND2_X1 U843 ( .A1(n767), .A2(n885), .ZN(n999) );
  NAND2_X1 U844 ( .A1(n768), .A2(n999), .ZN(n769) );
  NAND2_X1 U845 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U846 ( .A(n772), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U847 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U848 ( .A(G57), .ZN(G237) );
  INV_X1 U849 ( .A(G132), .ZN(G219) );
  INV_X1 U850 ( .A(G82), .ZN(G220) );
  NAND2_X1 U851 ( .A1(G7), .A2(G661), .ZN(n773) );
  XNOR2_X1 U852 ( .A(n773), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U853 ( .A(G223), .ZN(n839) );
  NAND2_X1 U854 ( .A1(n839), .A2(G567), .ZN(n774) );
  XNOR2_X1 U855 ( .A(n774), .B(KEYINPUT71), .ZN(n775) );
  XNOR2_X1 U856 ( .A(KEYINPUT11), .B(n775), .ZN(G234) );
  INV_X1 U857 ( .A(G860), .ZN(n783) );
  OR2_X1 U858 ( .A1(n1013), .A2(n783), .ZN(G153) );
  NAND2_X1 U859 ( .A1(G301), .A2(G868), .ZN(n777) );
  OR2_X1 U860 ( .A1(n1019), .A2(G868), .ZN(n776) );
  NAND2_X1 U861 ( .A1(n777), .A2(n776), .ZN(G284) );
  NOR2_X1 U862 ( .A1(G868), .A2(G299), .ZN(n778) );
  XNOR2_X1 U863 ( .A(n778), .B(KEYINPUT74), .ZN(n781) );
  INV_X1 U864 ( .A(G868), .ZN(n779) );
  NOR2_X1 U865 ( .A1(n779), .A2(G286), .ZN(n780) );
  NOR2_X1 U866 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U867 ( .A(KEYINPUT75), .B(n782), .Z(G297) );
  NAND2_X1 U868 ( .A1(n783), .A2(G559), .ZN(n784) );
  NAND2_X1 U869 ( .A1(n784), .A2(n1019), .ZN(n785) );
  XNOR2_X1 U870 ( .A(n785), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U871 ( .A1(G868), .A2(n1013), .ZN(n788) );
  NAND2_X1 U872 ( .A1(n1019), .A2(G868), .ZN(n786) );
  NOR2_X1 U873 ( .A1(G559), .A2(n786), .ZN(n787) );
  NOR2_X1 U874 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U875 ( .A(KEYINPUT76), .B(n789), .ZN(G282) );
  NAND2_X1 U876 ( .A1(G135), .A2(n516), .ZN(n791) );
  NAND2_X1 U877 ( .A1(G111), .A2(n911), .ZN(n790) );
  NAND2_X1 U878 ( .A1(n791), .A2(n790), .ZN(n797) );
  NAND2_X1 U879 ( .A1(G123), .A2(n517), .ZN(n792) );
  XNOR2_X1 U880 ( .A(n792), .B(KEYINPUT18), .ZN(n795) );
  NAND2_X1 U881 ( .A1(G99), .A2(n907), .ZN(n793) );
  XOR2_X1 U882 ( .A(KEYINPUT77), .B(n793), .Z(n794) );
  NAND2_X1 U883 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U884 ( .A1(n797), .A2(n796), .ZN(n984) );
  XNOR2_X1 U885 ( .A(n984), .B(G2096), .ZN(n798) );
  XNOR2_X1 U886 ( .A(n798), .B(KEYINPUT78), .ZN(n800) );
  INV_X1 U887 ( .A(G2100), .ZN(n799) );
  NAND2_X1 U888 ( .A1(n800), .A2(n799), .ZN(G156) );
  NAND2_X1 U889 ( .A1(G559), .A2(n1019), .ZN(n801) );
  XNOR2_X1 U890 ( .A(n801), .B(n1013), .ZN(n822) );
  NOR2_X1 U891 ( .A1(n822), .A2(G860), .ZN(n812) );
  NAND2_X1 U892 ( .A1(G67), .A2(n802), .ZN(n805) );
  NAND2_X1 U893 ( .A1(G55), .A2(n803), .ZN(n804) );
  NAND2_X1 U894 ( .A1(n805), .A2(n804), .ZN(n811) );
  NAND2_X1 U895 ( .A1(G93), .A2(n806), .ZN(n809) );
  NAND2_X1 U896 ( .A1(G80), .A2(n807), .ZN(n808) );
  NAND2_X1 U897 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U898 ( .A1(n811), .A2(n810), .ZN(n814) );
  XNOR2_X1 U899 ( .A(n812), .B(n814), .ZN(G145) );
  NOR2_X1 U900 ( .A1(G868), .A2(n814), .ZN(n813) );
  XNOR2_X1 U901 ( .A(n813), .B(KEYINPUT83), .ZN(n825) );
  XNOR2_X1 U902 ( .A(G166), .B(n814), .ZN(n820) );
  XNOR2_X1 U903 ( .A(n815), .B(G290), .ZN(n818) );
  XNOR2_X1 U904 ( .A(KEYINPUT82), .B(KEYINPUT19), .ZN(n816) );
  XNOR2_X1 U905 ( .A(n816), .B(G305), .ZN(n817) );
  XNOR2_X1 U906 ( .A(n818), .B(n817), .ZN(n819) );
  XNOR2_X1 U907 ( .A(n820), .B(n819), .ZN(n821) );
  XNOR2_X1 U908 ( .A(n821), .B(G288), .ZN(n921) );
  XNOR2_X1 U909 ( .A(n921), .B(n822), .ZN(n823) );
  NAND2_X1 U910 ( .A1(G868), .A2(n823), .ZN(n824) );
  NAND2_X1 U911 ( .A1(n825), .A2(n824), .ZN(G295) );
  NAND2_X1 U912 ( .A1(G2084), .A2(G2078), .ZN(n827) );
  XOR2_X1 U913 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n826) );
  XNOR2_X1 U914 ( .A(n827), .B(n826), .ZN(n828) );
  NAND2_X1 U915 ( .A1(G2090), .A2(n828), .ZN(n829) );
  XNOR2_X1 U916 ( .A(KEYINPUT21), .B(n829), .ZN(n830) );
  NAND2_X1 U917 ( .A1(n830), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U918 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U919 ( .A1(G220), .A2(G219), .ZN(n831) );
  XOR2_X1 U920 ( .A(KEYINPUT22), .B(n831), .Z(n832) );
  NOR2_X1 U921 ( .A1(G218), .A2(n832), .ZN(n833) );
  NAND2_X1 U922 ( .A1(G96), .A2(n833), .ZN(n843) );
  NAND2_X1 U923 ( .A1(n843), .A2(G2106), .ZN(n837) );
  NAND2_X1 U924 ( .A1(G120), .A2(G108), .ZN(n834) );
  NOR2_X1 U925 ( .A1(G237), .A2(n834), .ZN(n835) );
  NAND2_X1 U926 ( .A1(G69), .A2(n835), .ZN(n844) );
  NAND2_X1 U927 ( .A1(n844), .A2(G567), .ZN(n836) );
  NAND2_X1 U928 ( .A1(n837), .A2(n836), .ZN(n845) );
  NAND2_X1 U929 ( .A1(G483), .A2(G661), .ZN(n838) );
  NOR2_X1 U930 ( .A1(n845), .A2(n838), .ZN(n842) );
  NAND2_X1 U931 ( .A1(n842), .A2(G36), .ZN(G176) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n839), .ZN(G217) );
  AND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n840) );
  NAND2_X1 U934 ( .A1(G661), .A2(n840), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n841) );
  NAND2_X1 U936 ( .A1(n842), .A2(n841), .ZN(G188) );
  XOR2_X1 U937 ( .A(G108), .B(KEYINPUT114), .Z(G238) );
  INV_X1 U939 ( .A(G120), .ZN(G236) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  NOR2_X1 U941 ( .A1(n844), .A2(n843), .ZN(G325) );
  INV_X1 U942 ( .A(G325), .ZN(G261) );
  INV_X1 U943 ( .A(n845), .ZN(G319) );
  XNOR2_X1 U944 ( .A(G2446), .B(G2451), .ZN(n855) );
  XOR2_X1 U945 ( .A(G2430), .B(G2443), .Z(n847) );
  XNOR2_X1 U946 ( .A(G2454), .B(G2435), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U948 ( .A(G2438), .B(KEYINPUT103), .Z(n849) );
  XNOR2_X1 U949 ( .A(G1341), .B(G1348), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U951 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U952 ( .A(G2427), .B(KEYINPUT104), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n856) );
  NAND2_X1 U955 ( .A1(n856), .A2(G14), .ZN(n857) );
  XNOR2_X1 U956 ( .A(KEYINPUT105), .B(n857), .ZN(G401) );
  XOR2_X1 U957 ( .A(G2096), .B(G2678), .Z(n859) );
  XNOR2_X1 U958 ( .A(G2090), .B(KEYINPUT43), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U960 ( .A(n860), .B(KEYINPUT42), .Z(n862) );
  XNOR2_X1 U961 ( .A(G2067), .B(G2072), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U963 ( .A(KEYINPUT106), .B(G2100), .Z(n864) );
  XNOR2_X1 U964 ( .A(G2084), .B(G2078), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n866), .B(n865), .ZN(G227) );
  XOR2_X1 U967 ( .A(G1961), .B(G1966), .Z(n868) );
  XNOR2_X1 U968 ( .A(G1996), .B(G1981), .ZN(n867) );
  XNOR2_X1 U969 ( .A(n868), .B(n867), .ZN(n872) );
  XOR2_X1 U970 ( .A(G1956), .B(G1971), .Z(n870) );
  XNOR2_X1 U971 ( .A(G1986), .B(G1976), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U973 ( .A(n872), .B(n871), .Z(n874) );
  XNOR2_X1 U974 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n873) );
  XNOR2_X1 U975 ( .A(n874), .B(n873), .ZN(n876) );
  XOR2_X1 U976 ( .A(G1991), .B(G2474), .Z(n875) );
  XNOR2_X1 U977 ( .A(n876), .B(n875), .ZN(G229) );
  NAND2_X1 U978 ( .A1(G136), .A2(n516), .ZN(n878) );
  NAND2_X1 U979 ( .A1(G112), .A2(n911), .ZN(n877) );
  NAND2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n884) );
  NAND2_X1 U981 ( .A1(G124), .A2(n517), .ZN(n879) );
  XNOR2_X1 U982 ( .A(n879), .B(KEYINPUT44), .ZN(n882) );
  NAND2_X1 U983 ( .A1(G100), .A2(n907), .ZN(n880) );
  XNOR2_X1 U984 ( .A(n880), .B(KEYINPUT108), .ZN(n881) );
  NAND2_X1 U985 ( .A1(n882), .A2(n881), .ZN(n883) );
  NOR2_X1 U986 ( .A1(n884), .A2(n883), .ZN(G162) );
  XNOR2_X1 U987 ( .A(G160), .B(n885), .ZN(n887) );
  XNOR2_X1 U988 ( .A(n887), .B(n886), .ZN(n892) );
  XNOR2_X1 U989 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n888), .B(G162), .ZN(n889) );
  XNOR2_X1 U991 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U992 ( .A(n892), .B(n891), .Z(n894) );
  XNOR2_X1 U993 ( .A(n894), .B(n893), .ZN(n905) );
  NAND2_X1 U994 ( .A1(G118), .A2(n911), .ZN(n896) );
  NAND2_X1 U995 ( .A1(G130), .A2(n517), .ZN(n895) );
  NAND2_X1 U996 ( .A1(n896), .A2(n895), .ZN(n903) );
  NAND2_X1 U997 ( .A1(n516), .A2(G142), .ZN(n897) );
  XNOR2_X1 U998 ( .A(KEYINPUT110), .B(n897), .ZN(n900) );
  NAND2_X1 U999 ( .A1(n907), .A2(G106), .ZN(n898) );
  XOR2_X1 U1000 ( .A(KEYINPUT109), .B(n898), .Z(n899) );
  NAND2_X1 U1001 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U1002 ( .A(n901), .B(KEYINPUT45), .Z(n902) );
  NOR2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1004 ( .A(n905), .B(n904), .Z(n917) );
  NAND2_X1 U1005 ( .A1(G139), .A2(n516), .ZN(n909) );
  NAND2_X1 U1006 ( .A1(G103), .A2(n907), .ZN(n908) );
  NAND2_X1 U1007 ( .A1(n909), .A2(n908), .ZN(n916) );
  NAND2_X1 U1008 ( .A1(n517), .A2(G127), .ZN(n910) );
  XOR2_X1 U1009 ( .A(KEYINPUT111), .B(n910), .Z(n913) );
  NAND2_X1 U1010 ( .A1(n911), .A2(G115), .ZN(n912) );
  NAND2_X1 U1011 ( .A1(n913), .A2(n912), .ZN(n914) );
  XOR2_X1 U1012 ( .A(KEYINPUT47), .B(n914), .Z(n915) );
  NOR2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(n1001) );
  XNOR2_X1 U1014 ( .A(n917), .B(n1001), .ZN(n918) );
  NOR2_X1 U1015 ( .A1(G37), .A2(n918), .ZN(G395) );
  XNOR2_X1 U1016 ( .A(n1013), .B(KEYINPUT112), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(G301), .B(n1019), .ZN(n919) );
  XNOR2_X1 U1018 ( .A(n920), .B(n919), .ZN(n923) );
  XNOR2_X1 U1019 ( .A(G286), .B(n921), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(n923), .B(n922), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(G37), .A2(n924), .ZN(G397) );
  NOR2_X1 U1022 ( .A1(G227), .A2(G229), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(n925), .B(KEYINPUT49), .ZN(n926) );
  NOR2_X1 U1024 ( .A1(G401), .A2(n926), .ZN(n927) );
  NAND2_X1 U1025 ( .A1(G319), .A2(n927), .ZN(n928) );
  XNOR2_X1 U1026 ( .A(KEYINPUT113), .B(n928), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(G395), .A2(G397), .ZN(n929) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(G225) );
  INV_X1 U1029 ( .A(G225), .ZN(G308) );
  INV_X1 U1030 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1031 ( .A(G1981), .B(G6), .ZN(n932) );
  XNOR2_X1 U1032 ( .A(G1341), .B(G19), .ZN(n931) );
  NOR2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1034 ( .A(KEYINPUT126), .B(n933), .ZN(n936) );
  XNOR2_X1 U1035 ( .A(n934), .B(G20), .ZN(n935) );
  NAND2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n939) );
  XOR2_X1 U1037 ( .A(KEYINPUT59), .B(G1348), .Z(n937) );
  XNOR2_X1 U1038 ( .A(G4), .B(n937), .ZN(n938) );
  NOR2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(KEYINPUT60), .B(n940), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(G1966), .B(G21), .ZN(n942) );
  XNOR2_X1 U1042 ( .A(G5), .B(G1961), .ZN(n941) );
  NOR2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n952) );
  XNOR2_X1 U1045 ( .A(G1986), .B(G24), .ZN(n946) );
  XNOR2_X1 U1046 ( .A(G22), .B(G1971), .ZN(n945) );
  NOR2_X1 U1047 ( .A1(n946), .A2(n945), .ZN(n949) );
  XNOR2_X1 U1048 ( .A(G1976), .B(KEYINPUT127), .ZN(n947) );
  XNOR2_X1 U1049 ( .A(n947), .B(G23), .ZN(n948) );
  NAND2_X1 U1050 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1051 ( .A(KEYINPUT58), .B(n950), .ZN(n951) );
  NOR2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1053 ( .A(KEYINPUT61), .B(n953), .Z(n954) );
  NOR2_X1 U1054 ( .A1(G16), .A2(n954), .ZN(n983) );
  XNOR2_X1 U1055 ( .A(G29), .B(KEYINPUT123), .ZN(n980) );
  XNOR2_X1 U1056 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n1008) );
  XOR2_X1 U1057 ( .A(G2090), .B(G35), .Z(n958) );
  XNOR2_X1 U1058 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n955) );
  XNOR2_X1 U1059 ( .A(n955), .B(G34), .ZN(n956) );
  XNOR2_X1 U1060 ( .A(n956), .B(G2084), .ZN(n957) );
  NAND2_X1 U1061 ( .A1(n958), .A2(n957), .ZN(n976) );
  XNOR2_X1 U1062 ( .A(G1991), .B(G25), .ZN(n960) );
  XNOR2_X1 U1063 ( .A(G33), .B(G2072), .ZN(n959) );
  NOR2_X1 U1064 ( .A1(n960), .A2(n959), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(G32), .B(n961), .ZN(n962) );
  NAND2_X1 U1066 ( .A1(n962), .A2(G28), .ZN(n966) );
  XOR2_X1 U1067 ( .A(KEYINPUT118), .B(n963), .Z(n964) );
  XNOR2_X1 U1068 ( .A(G26), .B(n964), .ZN(n965) );
  NOR2_X1 U1069 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1070 ( .A1(n968), .A2(n967), .ZN(n972) );
  XNOR2_X1 U1071 ( .A(G27), .B(n969), .ZN(n970) );
  XNOR2_X1 U1072 ( .A(KEYINPUT119), .B(n970), .ZN(n971) );
  NOR2_X1 U1073 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1074 ( .A(KEYINPUT53), .B(n973), .ZN(n974) );
  XNOR2_X1 U1075 ( .A(KEYINPUT120), .B(n974), .ZN(n975) );
  NOR2_X1 U1076 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1077 ( .A(n1008), .B(n977), .Z(n978) );
  XNOR2_X1 U1078 ( .A(n978), .B(KEYINPUT122), .ZN(n979) );
  NAND2_X1 U1079 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1080 ( .A1(n981), .A2(G11), .ZN(n982) );
  NOR2_X1 U1081 ( .A1(n983), .A2(n982), .ZN(n1012) );
  NOR2_X1 U1082 ( .A1(n985), .A2(n984), .ZN(n989) );
  XOR2_X1 U1083 ( .A(G160), .B(G2084), .Z(n986) );
  NOR2_X1 U1084 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1085 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1086 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1087 ( .A(KEYINPUT115), .B(n992), .ZN(n997) );
  XOR2_X1 U1088 ( .A(G2090), .B(G162), .Z(n993) );
  NOR2_X1 U1089 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1090 ( .A(KEYINPUT51), .B(n995), .ZN(n996) );
  NOR2_X1 U1091 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1092 ( .A(n998), .B(KEYINPUT116), .ZN(n1000) );
  NAND2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1006) );
  XOR2_X1 U1094 ( .A(G2072), .B(n1001), .Z(n1003) );
  NOR2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1096 ( .A(KEYINPUT50), .B(n1004), .Z(n1005) );
  NOR2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1098 ( .A(KEYINPUT52), .B(n1007), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1010), .A2(G29), .ZN(n1011) );
  NAND2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1039) );
  XOR2_X1 U1102 ( .A(KEYINPUT56), .B(G16), .Z(n1037) );
  XOR2_X1 U1103 ( .A(G1341), .B(n1013), .Z(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1034) );
  XOR2_X1 U1105 ( .A(G1966), .B(G168), .Z(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1107 ( .A(KEYINPUT57), .B(n1018), .Z(n1032) );
  XNOR2_X1 U1108 ( .A(n1019), .B(G1348), .ZN(n1023) );
  AND2_X1 U1109 ( .A1(G303), .A2(G1971), .ZN(n1020) );
  NOR2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1025) );
  XNOR2_X1 U1112 ( .A(G1956), .B(G299), .ZN(n1024) );
  NOR2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1027) );
  NAND2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1030) );
  XOR2_X1 U1115 ( .A(G1961), .B(G171), .Z(n1028) );
  XNOR2_X1 U1116 ( .A(KEYINPUT124), .B(n1028), .ZN(n1029) );
  NOR2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1118 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1119 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XOR2_X1 U1120 ( .A(KEYINPUT125), .B(n1035), .Z(n1036) );
  NOR2_X1 U1121 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NOR2_X1 U1122 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XNOR2_X1 U1123 ( .A(n1040), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1124 ( .A(G311), .ZN(G150) );
endmodule

