//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 1 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n554, new_n556, new_n557, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1163, new_n1164;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT67), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND3_X1   g037(.A1(KEYINPUT68), .A2(G113), .A3(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(KEYINPUT68), .B1(G113), .B2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n462), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n466), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n473), .B1(KEYINPUT3), .B2(new_n468), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n475));
  OAI211_X1 g050(.A(G137), .B(new_n472), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G101), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n471), .B1(new_n478), .B2(new_n462), .ZN(G160));
  OAI21_X1  g054(.A(KEYINPUT69), .B1(new_n466), .B2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n467), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n481), .A2(new_n472), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n482), .A2(new_n462), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  NOR2_X1   g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(new_n462), .B2(G112), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n485), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NAND4_X1  g067(.A1(new_n481), .A2(G126), .A3(G2105), .A4(new_n472), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n481), .A2(new_n462), .A3(new_n472), .A4(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n467), .A2(new_n469), .A3(new_n462), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n494), .B1(new_n498), .B2(new_n495), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(G2104), .C1(G114), .C2(new_n462), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n493), .A2(new_n497), .A3(new_n499), .A4(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  NAND2_X1  g078(.A1(G75), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT70), .A3(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G62), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G651), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n512), .B(new_n513), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n509), .A2(new_n517), .ZN(new_n518));
  XOR2_X1   g093(.A(KEYINPUT71), .B(G88), .Z(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n517), .A2(new_n507), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n514), .A2(new_n520), .A3(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND2_X1  g099(.A1(new_n521), .A2(G51), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n506), .A2(new_n508), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n525), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n518), .A2(G89), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n530), .A2(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  NAND2_X1  g108(.A1(new_n518), .A2(G90), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  INV_X1    g110(.A(new_n521), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n509), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n537), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  NAND2_X1  g119(.A1(new_n518), .A2(G81), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT73), .B(G43), .Z(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n536), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(G651), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n526), .A2(G56), .ZN(new_n549));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(G188));
  NAND2_X1  g133(.A1(new_n521), .A2(G53), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT9), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n518), .A2(G91), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT74), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n509), .B(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n563), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n560), .B(new_n561), .C1(new_n564), .C2(new_n548), .ZN(G299));
  OAI21_X1  g140(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n566), .A2(KEYINPUT75), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n518), .A2(G87), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(KEYINPUT75), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n521), .A2(G49), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n567), .A2(new_n568), .A3(new_n569), .A4(new_n570), .ZN(G288));
  NAND3_X1  g146(.A1(new_n506), .A2(new_n508), .A3(G61), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n548), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n506), .A2(new_n508), .A3(G86), .ZN(new_n575));
  NAND2_X1  g150(.A1(G48), .A2(G543), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n517), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  XOR2_X1   g153(.A(new_n578), .B(KEYINPUT76), .Z(G305));
  NAND2_X1  g154(.A1(new_n518), .A2(G85), .ZN(new_n580));
  INV_X1    g155(.A(G47), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n581), .B2(new_n536), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n526), .A2(G60), .ZN(new_n583));
  NAND2_X1  g158(.A1(G72), .A2(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n548), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n518), .A2(G92), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n521), .A2(G54), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n563), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n591), .B(new_n592), .C1(new_n548), .C2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT77), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n595), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n588), .B1(new_n599), .B2(G868), .ZN(G284));
  XNOR2_X1  g175(.A(G284), .B(KEYINPUT78), .ZN(G321));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(G299), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n602), .B2(G168), .ZN(G297));
  OAI21_X1  g179(.A(new_n603), .B1(new_n602), .B2(G168), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G860), .ZN(G148));
  INV_X1    g182(.A(new_n552), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(new_n602), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n598), .A2(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n602), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g187(.A1(new_n462), .A2(G111), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT80), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n468), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI221_X1 g190(.A(new_n615), .B1(new_n614), .B2(new_n613), .C1(G99), .C2(G2105), .ZN(new_n616));
  INV_X1    g191(.A(G123), .ZN(new_n617));
  INV_X1    g192(.A(G135), .ZN(new_n618));
  OAI221_X1 g193(.A(new_n616), .B1(new_n483), .B2(new_n617), .C1(new_n618), .C2(new_n486), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT81), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2096), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n498), .A2(new_n468), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT13), .B(G2100), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n621), .A2(new_n626), .ZN(G156));
  XNOR2_X1  g202(.A(G2427), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2430), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT15), .B(G2435), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(KEYINPUT14), .ZN(new_n632));
  XOR2_X1   g207(.A(G2451), .B(G2454), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n634), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G1341), .B(G1348), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT82), .ZN(new_n640));
  INV_X1    g215(.A(G14), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n637), .A2(new_n638), .ZN(new_n642));
  NOR3_X1   g217(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(G401));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2067), .B(G2678), .Z(new_n646));
  NOR2_X1   g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n645), .A2(new_n646), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT17), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT18), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2072), .B(G2078), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n652), .B(new_n653), .C1(new_n651), .C2(new_n647), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n653), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2096), .B(G2100), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT83), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(G227));
  XNOR2_X1  g233(.A(G1971), .B(G1976), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  XOR2_X1   g235(.A(G1956), .B(G2474), .Z(new_n661));
  XOR2_X1   g236(.A(G1961), .B(G1966), .Z(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n665));
  INV_X1    g240(.A(new_n660), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n661), .A2(new_n662), .ZN(new_n667));
  AOI22_X1  g242(.A1(new_n664), .A2(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n669), .A2(new_n660), .A3(new_n663), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n668), .B(new_n670), .C1(new_n664), .C2(new_n665), .ZN(new_n671));
  XOR2_X1   g246(.A(G1991), .B(G1996), .Z(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT85), .B(G1986), .ZN(new_n676));
  INV_X1    g251(.A(G1981), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(G229));
  XNOR2_X1  g254(.A(KEYINPUT31), .B(G11), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT96), .Z(new_n681));
  INV_X1    g256(.A(G29), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G33), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n487), .A2(G139), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT91), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n467), .A2(new_n469), .A3(G127), .ZN(new_n686));
  INV_X1    g261(.A(G115), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n687), .B2(new_n468), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G2105), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT25), .Z(new_n691));
  NAND3_X1  g266(.A1(new_n685), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(KEYINPUT92), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT92), .ZN(new_n694));
  NAND4_X1  g269(.A1(new_n685), .A2(new_n694), .A3(new_n689), .A4(new_n691), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n683), .B1(new_n696), .B2(new_n682), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(G2072), .Z(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT30), .B(G28), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(new_n682), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT86), .B(G29), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G19), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(new_n552), .B2(new_n703), .ZN(new_n705));
  OAI221_X1 g280(.A(new_n700), .B1(new_n619), .B2(new_n702), .C1(new_n705), .C2(G1341), .ZN(new_n706));
  NOR2_X1   g281(.A1(G5), .A2(G16), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G171), .B2(G16), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(G1961), .ZN(new_n709));
  AOI211_X1 g284(.A(new_n706), .B(new_n709), .C1(G1341), .C2(new_n705), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n487), .A2(G141), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n484), .A2(G129), .ZN(new_n712));
  NAND3_X1  g287(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT94), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT93), .B(KEYINPUT26), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n711), .A2(new_n712), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G29), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G29), .B2(G32), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT27), .B(G1996), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT95), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n502), .A2(new_n701), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n702), .A2(G27), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT24), .B(G34), .ZN(new_n730));
  AOI22_X1  g305(.A1(G160), .A2(G29), .B1(new_n702), .B2(new_n730), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n729), .A2(G2078), .B1(G2084), .B2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G2078), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n721), .A2(new_n724), .B1(new_n733), .B2(new_n728), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n710), .A2(new_n725), .A3(new_n732), .A4(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(G16), .A2(G21), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G168), .B2(G16), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1966), .ZN(new_n738));
  OR2_X1    g313(.A1(G104), .A2(G2105), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n739), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n740));
  INV_X1    g315(.A(G128), .ZN(new_n741));
  INV_X1    g316(.A(G140), .ZN(new_n742));
  OAI221_X1 g317(.A(new_n740), .B1(new_n483), .B2(new_n741), .C1(new_n742), .C2(new_n486), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G29), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n702), .A2(KEYINPUT28), .A3(G26), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(KEYINPUT28), .B1(new_n702), .B2(G26), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G2067), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n731), .A2(G2084), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(KEYINPUT97), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n708), .A2(G1961), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(KEYINPUT97), .B2(new_n750), .ZN(new_n754));
  NOR4_X1   g329(.A1(new_n735), .A2(new_n738), .A3(new_n752), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n703), .A2(G4), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n599), .B2(new_n703), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(G1348), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n702), .A2(G35), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G162), .B2(new_n702), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT29), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G2090), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT98), .B(KEYINPUT23), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n703), .A2(G20), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G299), .B2(G16), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(G1956), .Z(new_n767));
  NOR2_X1   g342(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n698), .A2(new_n755), .A3(new_n758), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n484), .A2(G119), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n487), .A2(G131), .ZN(new_n771));
  NOR2_X1   g346(.A1(G95), .A2(G2105), .ZN(new_n772));
  OAI21_X1  g347(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n770), .B(new_n771), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT87), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(new_n701), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G25), .B2(new_n701), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT35), .B(G1991), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n703), .A2(G24), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n586), .B2(new_n703), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(G1986), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n781), .B2(new_n783), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n703), .A2(G23), .ZN(new_n789));
  INV_X1    g364(.A(G288), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(new_n703), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT89), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT33), .B(G1976), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n792), .B(new_n793), .Z(new_n794));
  NAND2_X1  g369(.A1(new_n703), .A2(G22), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G166), .B2(new_n703), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n796), .A2(G1971), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(G1971), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n703), .A2(G6), .ZN(new_n799));
  INV_X1    g374(.A(G305), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n703), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT32), .B(G1981), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n794), .A2(new_n797), .A3(new_n798), .A4(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT88), .B(KEYINPUT34), .ZN(new_n805));
  AOI211_X1 g380(.A(new_n784), .B(new_n788), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n786), .A2(G1986), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n792), .A2(new_n793), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n792), .A2(new_n793), .ZN(new_n810));
  AND3_X1   g385(.A1(new_n809), .A2(new_n798), .A3(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n805), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n811), .A2(new_n812), .A3(new_n797), .A4(new_n803), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n806), .A2(new_n807), .A3(new_n808), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n804), .A2(new_n805), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n784), .A2(new_n788), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n815), .A2(new_n808), .A3(new_n813), .A4(new_n816), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n817), .A2(KEYINPUT90), .A3(KEYINPUT36), .ZN(new_n818));
  AOI211_X1 g393(.A(new_n681), .B(new_n769), .C1(new_n814), .C2(new_n818), .ZN(G311));
  AOI21_X1  g394(.A(new_n769), .B1(new_n814), .B2(new_n818), .ZN(new_n820));
  INV_X1    g395(.A(new_n681), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(G150));
  NAND2_X1  g397(.A1(G80), .A2(G543), .ZN(new_n823));
  INV_X1    g398(.A(G67), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n509), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G651), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT99), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT100), .B(G93), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n518), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(G55), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n827), .B(new_n829), .C1(new_n830), .C2(new_n536), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT37), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n599), .A2(G559), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT38), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n831), .A2(new_n552), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n831), .A2(new_n552), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT39), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n835), .B(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n833), .B1(new_n841), .B2(G860), .ZN(G145));
  XNOR2_X1  g417(.A(new_n778), .B(new_n624), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n462), .A2(G118), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT104), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n468), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI221_X1 g421(.A(new_n846), .B1(new_n845), .B2(new_n844), .C1(G106), .C2(G2105), .ZN(new_n847));
  INV_X1    g422(.A(G130), .ZN(new_n848));
  INV_X1    g423(.A(G142), .ZN(new_n849));
  OAI221_X1 g424(.A(new_n847), .B1(new_n483), .B2(new_n848), .C1(new_n849), .C2(new_n486), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n843), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n497), .A2(new_n499), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT101), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n493), .A2(new_n854), .A3(new_n501), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n854), .B1(new_n493), .B2(new_n501), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n853), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n743), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n719), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n696), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT102), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n858), .B(new_n718), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n693), .A2(new_n695), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT103), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n619), .B(G160), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(G162), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n861), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n868), .B1(new_n861), .B2(new_n866), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n851), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n861), .A2(new_n866), .ZN(new_n872));
  INV_X1    g447(.A(new_n868), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n851), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n861), .A2(new_n866), .A3(new_n868), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(G37), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n871), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(KEYINPUT40), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT40), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n871), .A2(new_n877), .A3(new_n881), .A4(new_n878), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(G395));
  XNOR2_X1  g458(.A(new_n610), .B(new_n839), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n594), .A2(G299), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n594), .A2(G299), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT105), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n885), .A2(new_n886), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT41), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n887), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n889), .B1(new_n884), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT42), .ZN(new_n896));
  NAND2_X1  g471(.A1(G166), .A2(G288), .ZN(new_n897));
  NAND2_X1  g472(.A1(G303), .A2(new_n790), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(G305), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(G305), .B1(new_n897), .B2(new_n898), .ZN(new_n901));
  OAI21_X1  g476(.A(G290), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n901), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n903), .A2(new_n586), .A3(new_n899), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n889), .B(new_n906), .C1(new_n884), .C2(new_n894), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n896), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n905), .B1(new_n896), .B2(new_n907), .ZN(new_n909));
  OAI21_X1  g484(.A(G868), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n831), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n910), .B1(G868), .B2(new_n911), .ZN(G295));
  OAI21_X1  g487(.A(new_n910), .B1(G868), .B2(new_n911), .ZN(G331));
  XNOR2_X1  g488(.A(G301), .B(G286), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n838), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n915), .B1(new_n916), .B2(new_n836), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n837), .A2(new_n838), .A3(new_n914), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n918), .A3(KEYINPUT106), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n839), .A2(new_n920), .A3(new_n915), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n919), .A2(new_n893), .A3(new_n891), .A4(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n917), .A2(new_n918), .A3(new_n890), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n905), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n919), .A2(new_n921), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n891), .A2(new_n893), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n917), .A2(new_n918), .ZN(new_n927));
  AOI22_X1  g502(.A1(new_n925), .A2(new_n888), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n878), .B(new_n924), .C1(new_n928), .C2(new_n905), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT107), .B1(new_n929), .B2(KEYINPUT43), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n924), .A2(new_n878), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n905), .B1(new_n922), .B2(new_n923), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT43), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n931), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n925), .A2(new_n888), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n894), .B1(new_n917), .B2(new_n918), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n904), .B(new_n902), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n934), .A2(new_n937), .A3(new_n938), .A4(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n930), .A2(new_n933), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n939), .B1(new_n931), .B2(new_n932), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n944), .B1(new_n939), .B2(new_n929), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT44), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n946), .ZN(G397));
  XOR2_X1   g522(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n948));
  INV_X1    g523(.A(G1384), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n948), .B1(new_n857), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT109), .B1(G160), .B2(G40), .ZN(new_n951));
  AOI21_X1  g526(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n953));
  INV_X1    g528(.A(G40), .ZN(new_n954));
  NOR4_X1   g529(.A1(new_n952), .A2(new_n471), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n950), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(G1996), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n718), .B(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G2067), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n743), .B(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n779), .A2(new_n960), .A3(new_n783), .A4(new_n962), .ZN(new_n963));
  OR2_X1    g538(.A1(new_n743), .A2(G2067), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n958), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n958), .B1(new_n719), .B2(new_n962), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT126), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n957), .A2(new_n959), .ZN(new_n969));
  XOR2_X1   g544(.A(new_n969), .B(KEYINPUT46), .Z(new_n970));
  NOR2_X1   g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n971), .B(KEYINPUT47), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n960), .B(new_n962), .C1(new_n782), .C2(new_n778), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n779), .A2(new_n783), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n957), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n958), .A2(G1986), .A3(G290), .ZN(new_n976));
  XNOR2_X1  g551(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n976), .B(new_n977), .ZN(new_n978));
  AOI211_X1 g553(.A(new_n965), .B(new_n972), .C1(new_n975), .C2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(G303), .A2(G8), .ZN(new_n980));
  XOR2_X1   g555(.A(new_n980), .B(KEYINPUT55), .Z(new_n981));
  NAND3_X1  g556(.A1(new_n857), .A2(KEYINPUT45), .A3(new_n949), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n502), .A2(new_n949), .ZN(new_n983));
  INV_X1    g558(.A(new_n948), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n956), .A2(new_n982), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1971), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n493), .A2(new_n501), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT101), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n493), .A2(new_n854), .A3(new_n501), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n852), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n989), .B1(new_n993), .B2(G1384), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n857), .A2(KEYINPUT111), .A3(new_n949), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT50), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n983), .A2(KEYINPUT50), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n956), .A2(new_n997), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n996), .A2(G2090), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n988), .B1(new_n999), .B2(KEYINPUT112), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n1001));
  INV_X1    g576(.A(new_n995), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT111), .B1(new_n857), .B2(new_n949), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G2090), .ZN(new_n1005));
  INV_X1    g580(.A(new_n998), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g584(.A(G8), .B(new_n981), .C1(new_n1000), .C2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n994), .A2(new_n995), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n956), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT49), .B1(new_n578), .B2(new_n677), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT49), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1014), .B(G1981), .C1(new_n574), .C2(new_n577), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n578), .A2(new_n677), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT113), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1016), .B(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1012), .A2(new_n1019), .A3(G8), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n790), .A2(G1976), .ZN(new_n1021));
  INV_X1    g596(.A(G1976), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(G288), .B2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1012), .A2(G8), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1012), .A2(G8), .A3(new_n1021), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1020), .B(new_n1024), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n502), .A2(new_n1001), .A3(new_n949), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n956), .B(new_n1029), .C1(new_n1011), .C2(new_n1001), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n988), .B1(new_n1030), .B2(G2090), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G8), .ZN(new_n1032));
  INV_X1    g607(.A(new_n981), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n996), .A2(G2084), .A3(new_n998), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n994), .A2(new_n1036), .A3(new_n995), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n983), .A2(new_n984), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1038), .A2(new_n951), .A3(new_n955), .ZN(new_n1039));
  AOI21_X1  g614(.A(G1966), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(G8), .B1(new_n1035), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(G286), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1010), .A2(new_n1028), .A3(new_n1034), .A4(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT63), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(G8), .B1(new_n1000), .B2(new_n1009), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1044), .B1(new_n1046), .B2(new_n1033), .ZN(new_n1047));
  INV_X1    g622(.A(G8), .ZN(new_n1048));
  INV_X1    g623(.A(new_n988), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n999), .A2(KEYINPUT112), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1027), .B1(new_n1052), .B2(new_n981), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1047), .A2(new_n1053), .A3(new_n1042), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1045), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1020), .A2(new_n1022), .A3(new_n790), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n1017), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1012), .A2(KEYINPUT114), .A3(G8), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT114), .B1(new_n1012), .B2(G8), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n1010), .B2(new_n1027), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1061), .B(KEYINPUT115), .C1(new_n1010), .C2(new_n1027), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1037), .A2(new_n733), .A3(new_n1039), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT123), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT123), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1037), .A2(new_n1069), .A3(new_n733), .A4(new_n1039), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(KEYINPUT53), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1072));
  INV_X1    g647(.A(G1961), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n956), .A2(new_n982), .A3(new_n733), .A4(new_n985), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1072), .A2(new_n1073), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(G301), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  AND4_X1   g652(.A1(new_n1034), .A2(new_n1010), .A3(new_n1028), .A4(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT51), .ZN(new_n1079));
  NAND2_X1  g654(.A1(G286), .A2(G8), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G2084), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1004), .A2(new_n1084), .A3(new_n1006), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1085), .B1(new_n1086), .B2(G1966), .ZN(new_n1087));
  OAI211_X1 g662(.A(G8), .B(new_n1083), .C1(new_n1087), .C2(G286), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1041), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1087), .A2(G8), .A3(G286), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT62), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT62), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1088), .A2(new_n1089), .A3(new_n1093), .A4(new_n1090), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1078), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1055), .A2(new_n1066), .A3(new_n1095), .ZN(new_n1096));
  XOR2_X1   g671(.A(G299), .B(KEYINPUT57), .Z(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT116), .B(G1956), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1030), .A2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n1100), .B(KEYINPUT117), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n986), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1097), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1012), .A2(KEYINPUT118), .ZN(new_n1104));
  NAND2_X1  g679(.A1(G160), .A2(G40), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n953), .ZN(new_n1106));
  INV_X1    g681(.A(new_n955), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1108), .B1(new_n994), .B2(new_n995), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1104), .A2(new_n1111), .A3(new_n961), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n996), .A2(new_n998), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1115), .A2(G1348), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1104), .A2(new_n1111), .A3(KEYINPUT119), .A4(new_n961), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1099), .A2(new_n1097), .A3(new_n1102), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1103), .B1(new_n1120), .B2(new_n599), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n598), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .A4(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n598), .A2(new_n1122), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n552), .A2(KEYINPUT120), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT58), .B(G1341), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1128), .B1(new_n1104), .B2(new_n1111), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n986), .A2(G1996), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1127), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT59), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1133), .B(new_n1127), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1126), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1099), .A2(new_n1097), .A3(new_n1102), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1138), .A2(new_n1103), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT61), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1121), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1071), .A2(G301), .A3(new_n1076), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1075), .A2(new_n1074), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT53), .B1(KEYINPUT124), .B2(G2078), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n950), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1105), .B1(KEYINPUT124), .B2(G2078), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1145), .A2(new_n982), .A3(new_n1146), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1143), .B(new_n1147), .C1(new_n1115), .C2(G1961), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(G171), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1142), .A2(KEYINPUT54), .A3(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT125), .ZN(new_n1151));
  XOR2_X1   g726(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1152));
  NOR2_X1   g727(.A1(new_n1148), .A2(G171), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1152), .B1(new_n1077), .B2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1154), .A2(new_n1053), .A3(new_n1091), .A4(new_n1034), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1096), .B1(new_n1141), .B2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n586), .B(G1986), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n975), .B1(new_n958), .B2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1159), .B(KEYINPUT110), .Z(new_n1160));
  OAI21_X1  g735(.A(new_n979), .B1(new_n1157), .B2(new_n1160), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g736(.A1(G227), .A2(new_n460), .ZN(new_n1163));
  NOR2_X1   g737(.A1(G401), .A2(G229), .ZN(new_n1164));
  AND4_X1   g738(.A1(new_n879), .A2(new_n941), .A3(new_n1163), .A4(new_n1164), .ZN(G308));
  NAND4_X1  g739(.A1(new_n879), .A2(new_n941), .A3(new_n1163), .A4(new_n1164), .ZN(G225));
endmodule


