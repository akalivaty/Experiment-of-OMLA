//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT64), .B(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT65), .Z(new_n215));
  XOR2_X1   g0015(.A(KEYINPUT67), .B(G244), .Z(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT66), .B(G77), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G107), .A2(G264), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n209), .B1(new_n213), .B2(new_n215), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G87), .B(G97), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  OR2_X1    g0042(.A1(KEYINPUT68), .A2(G1), .ZN(new_n243));
  NAND2_X1  g0043(.A1(KEYINPUT68), .A2(G1), .ZN(new_n244));
  NAND4_X1  g0044(.A1(new_n243), .A2(G13), .A3(G20), .A4(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(new_n202), .ZN(new_n247));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n211), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n243), .A2(new_n244), .ZN(new_n251));
  INV_X1    g0051(.A(G20), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n247), .B1(new_n202), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G33), .A3(new_n210), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n250), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  XOR2_X1   g0061(.A(new_n261), .B(KEYINPUT9), .Z(new_n262));
  INV_X1    g0062(.A(G190), .ZN(new_n263));
  AND2_X1   g0063(.A1(G1), .A2(G13), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  XOR2_X1   g0067(.A(KEYINPUT68), .B(G1), .Z(new_n268));
  NOR2_X1   g0068(.A1(G41), .A2(G45), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n267), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G226), .ZN(new_n272));
  INV_X1    g0072(.A(G274), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(new_n264), .B2(new_n265), .ZN(new_n274));
  INV_X1    g0074(.A(G1), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(new_n275), .A3(new_n270), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n278), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G223), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(new_n282), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G222), .A3(new_n278), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n284), .B(new_n286), .C1(new_n217), .C2(new_n285), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n277), .B1(new_n267), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n262), .B1(new_n263), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G200), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  OR3_X1    g0092(.A1(new_n290), .A2(KEYINPUT10), .A3(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(KEYINPUT10), .B1(new_n290), .B2(new_n292), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n289), .A2(G179), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n288), .A2(G169), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n296), .A2(new_n297), .A3(new_n261), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G68), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n258), .A2(G50), .B1(G20), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n210), .A2(G33), .ZN(new_n303));
  INV_X1    g0103(.A(G77), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n249), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT11), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n306), .B(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n246), .A2(new_n301), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n309), .A2(KEYINPUT72), .A3(KEYINPUT12), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(KEYINPUT12), .B1(new_n309), .B2(KEYINPUT72), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT71), .ZN(new_n313));
  INV_X1    g0113(.A(new_n253), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n313), .B1(new_n314), .B2(G68), .ZN(new_n315));
  NOR3_X1   g0115(.A1(new_n253), .A2(KEYINPUT71), .A3(new_n301), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n311), .A2(new_n312), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n308), .A2(new_n317), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n266), .B(G238), .C1(new_n251), .C2(new_n269), .ZN(new_n319));
  INV_X1    g0119(.A(G97), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n280), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(G226), .A2(G1698), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n322), .B1(new_n228), .B2(G1698), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n321), .B1(new_n323), .B2(new_n285), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n319), .B(new_n276), .C1(new_n324), .C2(new_n266), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT13), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT70), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n228), .A2(G1698), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(G226), .B2(G1698), .ZN(new_n329));
  AND2_X1   g0129(.A1(KEYINPUT3), .A2(G33), .ZN(new_n330));
  NOR2_X1   g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI22_X1  g0132(.A1(new_n329), .A2(new_n332), .B1(new_n280), .B2(new_n320), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n267), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT13), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n334), .A2(new_n335), .A3(new_n319), .A4(new_n276), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n326), .A2(new_n327), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n325), .A2(KEYINPUT70), .A3(KEYINPUT13), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(G200), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n326), .A2(G190), .A3(new_n336), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n318), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n326), .A2(G179), .A3(new_n336), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n337), .A2(G169), .A3(new_n338), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT14), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n337), .A2(KEYINPUT14), .A3(G169), .A4(new_n338), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n343), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n341), .B1(new_n348), .B2(new_n318), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT74), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n253), .A2(new_n256), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n245), .A2(new_n255), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n332), .A2(new_n210), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n281), .A2(new_n252), .A3(new_n282), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT7), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n355), .A2(new_n357), .A3(G68), .ZN(new_n358));
  AND2_X1   g0158(.A1(G58), .A2(G68), .ZN(new_n359));
  OAI21_X1  g0159(.A(G20), .B1(new_n359), .B2(new_n201), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT73), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n258), .A2(new_n361), .A3(G159), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n361), .B1(new_n258), .B2(G159), .ZN(new_n364));
  OAI211_X1 g0164(.A(KEYINPUT16), .B(new_n360), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n249), .B1(new_n358), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n252), .A2(KEYINPUT64), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT64), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G20), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n281), .A2(new_n367), .A3(new_n369), .A4(new_n282), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT7), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n332), .A2(new_n354), .A3(new_n252), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(G68), .A3(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n360), .B1(new_n363), .B2(new_n364), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT16), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n353), .B1(new_n366), .B2(new_n376), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n266), .B(G232), .C1(new_n251), .C2(new_n269), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n276), .ZN(new_n379));
  OR2_X1    g0179(.A1(G223), .A2(G1698), .ZN(new_n380));
  INV_X1    g0180(.A(G226), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(G1698), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n380), .B(new_n382), .C1(new_n330), .C2(new_n331), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G33), .A2(G87), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n266), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n291), .B1(new_n379), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n383), .A2(new_n384), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n267), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n388), .A2(new_n263), .A3(new_n276), .A4(new_n378), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT17), .ZN(new_n391));
  NOR3_X1   g0191(.A1(new_n377), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n353), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n354), .B1(new_n332), .B2(new_n210), .ZN(new_n395));
  NOR4_X1   g0195(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT7), .A4(G20), .ZN(new_n396));
  NOR3_X1   g0196(.A1(new_n395), .A2(new_n396), .A3(new_n301), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n394), .B1(new_n397), .B2(new_n374), .ZN(new_n398));
  INV_X1    g0198(.A(new_n365), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n355), .A2(new_n357), .A3(G68), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n250), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n393), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n386), .A2(new_n389), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT17), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n350), .B1(new_n392), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(G169), .B1(new_n379), .B2(new_n385), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n388), .A2(G179), .A3(new_n276), .A4(new_n378), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n402), .A2(new_n408), .A3(KEYINPUT18), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT18), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n406), .A2(new_n407), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n410), .B1(new_n377), .B2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n391), .B1(new_n377), .B2(new_n390), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n402), .A2(KEYINPUT17), .A3(new_n403), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n415), .A3(KEYINPUT74), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n405), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  XOR2_X1   g0217(.A(new_n255), .B(KEYINPUT69), .Z(new_n418));
  NOR3_X1   g0218(.A1(new_n418), .A2(G20), .A3(G33), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT15), .B(G87), .ZN(new_n420));
  OAI22_X1  g0220(.A1(new_n303), .A2(new_n420), .B1(new_n217), .B2(new_n210), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n249), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n314), .A2(G77), .B1(new_n246), .B2(new_n217), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n216), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n271), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(G232), .A2(G1698), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n278), .A2(G238), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n285), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(new_n267), .C1(G107), .C2(new_n285), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n426), .A2(new_n276), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n424), .B1(G190), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n291), .B2(new_n432), .ZN(new_n434));
  INV_X1    g0234(.A(G179), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(G169), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n431), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n424), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  NOR4_X1   g0240(.A1(new_n300), .A2(new_n349), .A3(new_n417), .A4(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n245), .A2(G107), .ZN(new_n442));
  XNOR2_X1  g0242(.A(new_n442), .B(KEYINPUT25), .ZN(new_n443));
  INV_X1    g0243(.A(G107), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n243), .A2(G33), .A3(new_n244), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n245), .A2(new_n250), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n443), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n367), .B(new_n369), .C1(new_n330), .C2(new_n331), .ZN(new_n448));
  INV_X1    g0248(.A(G87), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT22), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT22), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n285), .A2(new_n210), .A3(new_n451), .A4(G87), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  OR2_X1    g0253(.A1(KEYINPUT23), .A2(G107), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT23), .B1(new_n252), .B2(G107), .ZN(new_n455));
  OAI22_X1  g0255(.A1(new_n210), .A2(new_n454), .B1(KEYINPUT76), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(KEYINPUT76), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n252), .A2(G33), .A3(G116), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n453), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT24), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT24), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n453), .A2(new_n463), .A3(new_n460), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n447), .B1(new_n465), .B2(new_n249), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n243), .A2(G45), .A3(new_n244), .ZN(new_n467));
  AND2_X1   g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(G264), .B(new_n266), .C1(new_n467), .C2(new_n470), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT5), .B(G41), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n268), .A2(new_n274), .A3(G45), .A4(new_n472), .ZN(new_n473));
  MUX2_X1   g0273(.A(G250), .B(G257), .S(G1698), .Z(new_n474));
  AOI22_X1  g0274(.A1(new_n474), .A2(new_n285), .B1(G33), .B2(G294), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n471), .B(new_n473), .C1(new_n475), .C2(new_n266), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(KEYINPUT77), .A3(G169), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n474), .A2(new_n285), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G294), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n267), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n481), .A2(G179), .A3(new_n473), .A4(new_n471), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT77), .B1(new_n476), .B2(G169), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(KEYINPUT78), .B1(new_n466), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT78), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n250), .B1(new_n462), .B2(new_n464), .ZN(new_n488));
  OAI221_X1 g0288(.A(new_n487), .B1(new_n483), .B2(new_n484), .C1(new_n488), .C2(new_n447), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT21), .ZN(new_n490));
  INV_X1    g0290(.A(G116), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n246), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n245), .A2(new_n250), .A3(new_n445), .A4(G116), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G283), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n280), .A2(G97), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n210), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n248), .A2(new_n211), .B1(G20), .B2(new_n491), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT20), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n497), .A2(KEYINPUT20), .A3(new_n498), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n494), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G303), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n266), .B1(new_n332), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(G257), .A2(G1698), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n278), .A2(G264), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n285), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(G270), .B(new_n266), .C1(new_n467), .C2(new_n470), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n508), .A2(new_n473), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G169), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n490), .B1(new_n502), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n501), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n492), .B(new_n493), .C1(new_n513), .C2(new_n499), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n514), .A2(KEYINPUT21), .A3(G169), .A4(new_n510), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n510), .A2(G200), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n508), .A2(G190), .A3(new_n473), .A4(new_n509), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n502), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n510), .A2(new_n435), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n514), .ZN(new_n520));
  AND4_X1   g0320(.A1(new_n512), .A2(new_n515), .A3(new_n518), .A4(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n486), .A2(new_n489), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n476), .A2(new_n291), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT79), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT79), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n476), .A2(new_n525), .A3(new_n291), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n524), .B(new_n526), .C1(G190), .C2(new_n476), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n466), .A2(new_n527), .ZN(new_n528));
  OR2_X1    g0328(.A1(new_n446), .A2(new_n320), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n246), .A2(new_n320), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g0331(.A(KEYINPUT75), .B(KEYINPUT6), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n532), .A2(G97), .A3(new_n444), .ZN(new_n533));
  XOR2_X1   g0333(.A(G97), .B(G107), .Z(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n367), .A2(new_n369), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n371), .A2(G107), .A3(new_n372), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n258), .A2(G77), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n531), .B1(new_n540), .B2(new_n249), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n285), .A2(G244), .A3(new_n278), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT4), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n285), .A2(KEYINPUT4), .A3(G244), .A4(new_n278), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n283), .A2(G250), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .A4(new_n495), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n267), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n467), .A2(new_n470), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n550), .A2(new_n267), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G257), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n549), .A2(new_n473), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n437), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n548), .A2(new_n267), .B1(new_n551), .B2(G257), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n555), .A2(new_n435), .A3(new_n473), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n542), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n553), .A2(G200), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n555), .A2(G190), .A3(new_n473), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n559), .A3(new_n541), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n283), .A2(G244), .B1(G33), .B2(G116), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n285), .A2(G238), .A3(new_n278), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n266), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n268), .A2(new_n274), .A3(G45), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n467), .A2(G250), .A3(new_n266), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(G200), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n285), .A2(G244), .A3(G1698), .ZN(new_n568));
  NAND2_X1  g0368(.A1(G33), .A2(G116), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n562), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n267), .ZN(new_n571));
  INV_X1    g0371(.A(new_n566), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n572), .A3(G190), .ZN(new_n573));
  NOR2_X1   g0373(.A1(G97), .A2(G107), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n449), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT19), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n576), .A2(new_n280), .A3(new_n320), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n575), .B1(new_n577), .B2(new_n536), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n367), .A2(new_n369), .A3(G33), .A4(G97), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n576), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n285), .A2(new_n210), .A3(G68), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n582), .A2(new_n249), .B1(new_n246), .B2(new_n420), .ZN(new_n583));
  OR2_X1    g0383(.A1(new_n446), .A2(new_n449), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n567), .A2(new_n573), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n582), .A2(new_n249), .ZN(new_n586));
  OR2_X1    g0386(.A1(new_n446), .A2(new_n420), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n246), .A2(new_n420), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n437), .B1(new_n563), .B2(new_n566), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n571), .A2(new_n572), .A3(new_n435), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n585), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n528), .A2(new_n557), .A3(new_n560), .A4(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n522), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n441), .A2(new_n595), .ZN(G372));
  INV_X1    g0396(.A(new_n557), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n597), .A2(KEYINPUT26), .A3(new_n593), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT26), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n585), .A2(new_n592), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n599), .B1(new_n557), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n512), .A2(new_n515), .A3(new_n520), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n466), .A2(new_n485), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n602), .B(new_n592), .C1(new_n594), .C2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n441), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n348), .A2(new_n318), .ZN(new_n609));
  INV_X1    g0409(.A(new_n439), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n609), .B1(new_n341), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n405), .A2(new_n416), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n413), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n298), .B1(new_n613), .B2(new_n295), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n608), .A2(new_n614), .ZN(G369));
  AND2_X1   g0415(.A1(new_n486), .A2(new_n489), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n210), .A2(G13), .ZN(new_n617));
  OR3_X1    g0417(.A1(new_n617), .A2(KEYINPUT27), .A3(new_n251), .ZN(new_n618));
  OAI21_X1  g0418(.A(KEYINPUT27), .B1(new_n617), .B2(new_n251), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(new_n619), .A3(G213), .ZN(new_n620));
  INV_X1    g0420(.A(G343), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n603), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n616), .A2(new_n528), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n622), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n605), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g0427(.A(new_n627), .B(KEYINPUT81), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n616), .B(new_n528), .C1(new_n466), .C2(new_n625), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n605), .A2(new_n622), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n625), .A2(new_n502), .ZN(new_n633));
  MUX2_X1   g0433(.A(new_n521), .B(new_n604), .S(new_n633), .Z(new_n634));
  XNOR2_X1  g0434(.A(KEYINPUT80), .B(G330), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n629), .A2(new_n639), .ZN(G399));
  NAND3_X1  g0440(.A1(new_n574), .A2(new_n449), .A3(new_n491), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n641), .B(KEYINPUT82), .ZN(new_n642));
  INV_X1    g0442(.A(new_n207), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(G41), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n642), .A2(new_n275), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n214), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n645), .B1(new_n646), .B2(new_n644), .ZN(new_n647));
  XOR2_X1   g0447(.A(new_n647), .B(KEYINPUT28), .Z(new_n648));
  AND2_X1   g0448(.A1(new_n607), .A2(new_n625), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n616), .A2(new_n603), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n592), .B(new_n602), .C1(new_n650), .C2(new_n594), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n625), .ZN(new_n652));
  MUX2_X1   g0452(.A(new_n649), .B(new_n652), .S(KEYINPUT29), .Z(new_n653));
  INV_X1    g0453(.A(new_n476), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n563), .A2(new_n566), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n555), .A2(new_n519), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT30), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n571), .A2(new_n572), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(new_n476), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n660), .A2(KEYINPUT30), .A3(new_n555), .A4(new_n519), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n553), .A2(new_n476), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT83), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n510), .A2(new_n435), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n664), .B1(new_n655), .B2(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n659), .A2(KEYINPUT83), .A3(new_n435), .A4(new_n510), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n663), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n622), .B1(new_n662), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT31), .ZN(new_n670));
  AOI21_X1  g0470(.A(KEYINPUT84), .B1(new_n595), .B2(new_n625), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT84), .ZN(new_n672));
  NOR4_X1   g0472(.A1(new_n522), .A2(new_n594), .A3(new_n672), .A4(new_n622), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n670), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n636), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n653), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n648), .B1(new_n677), .B2(G1), .ZN(G364));
  INV_X1    g0478(.A(new_n617), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n275), .B1(new_n679), .B2(G45), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(new_n644), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n638), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n636), .B2(new_n634), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n210), .A2(G190), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(KEYINPUT88), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n291), .A2(G179), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(KEYINPUT88), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT89), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n690), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(G179), .A2(G200), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n686), .A2(new_n688), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AOI22_X1  g0497(.A1(new_n694), .A2(G283), .B1(G329), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT90), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n687), .A2(G20), .A3(G190), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n210), .B1(G190), .B2(new_n695), .ZN(new_n701));
  INV_X1    g0501(.A(G294), .ZN(new_n702));
  OAI221_X1 g0502(.A(new_n332), .B1(new_n503), .B2(new_n700), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n435), .A2(new_n291), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n685), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  XNOR2_X1  g0506(.A(KEYINPUT33), .B(G317), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n435), .A2(G200), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n536), .A2(G190), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n706), .A2(new_n707), .B1(G322), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G326), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n536), .A2(G190), .A3(new_n704), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n685), .A2(new_n708), .ZN(new_n715));
  OR2_X1    g0515(.A1(new_n715), .A2(KEYINPUT87), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(KEYINPUT87), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI211_X1 g0518(.A(new_n703), .B(new_n714), .C1(G311), .C2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n694), .A2(G107), .ZN(new_n720));
  INV_X1    g0520(.A(new_n718), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n217), .ZN(new_n722));
  OAI221_X1 g0522(.A(new_n285), .B1(new_n449), .B2(new_n700), .C1(new_n713), .C2(new_n202), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n701), .A2(new_n320), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(G58), .ZN(new_n726));
  OAI221_X1 g0526(.A(new_n725), .B1(new_n726), .B2(new_n709), .C1(new_n705), .C2(new_n301), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n722), .A2(new_n723), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(G159), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n696), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT32), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n699), .A2(new_n719), .B1(new_n720), .B2(new_n732), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n733), .A2(KEYINPUT91), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n264), .B1(new_n252), .B2(G169), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n735), .A2(KEYINPUT86), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(KEYINPUT86), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n733), .A2(KEYINPUT91), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n734), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n682), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n241), .A2(G45), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT85), .Z(new_n743));
  NOR2_X1   g0543(.A1(new_n643), .A2(new_n285), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n743), .B(new_n744), .C1(G45), .C2(new_n215), .ZN(new_n745));
  INV_X1    g0545(.A(G355), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n285), .A2(new_n207), .ZN(new_n747));
  OAI221_X1 g0547(.A(new_n745), .B1(G116), .B2(new_n207), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n738), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n741), .B1(new_n748), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n751), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n753), .B1(new_n634), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n684), .B1(new_n740), .B2(new_n755), .ZN(G396));
  NAND2_X1  g0556(.A1(new_n424), .A2(new_n622), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n610), .B1(new_n434), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n439), .A2(new_n622), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n607), .A2(new_n760), .A3(new_n625), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n760), .B(KEYINPUT93), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n761), .B1(new_n762), .B2(new_n649), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n682), .B1(new_n763), .B2(new_n675), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n764), .B1(new_n675), .B2(new_n763), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n738), .A2(new_n749), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n682), .B1(new_n767), .B2(G77), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n694), .A2(G87), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n702), .A2(new_n709), .B1(new_n713), .B2(new_n503), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n725), .B(new_n332), .C1(new_n444), .C2(new_n700), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n705), .B(KEYINPUT92), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n770), .B(new_n771), .C1(G283), .C2(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(G311), .A2(new_n697), .B1(new_n718), .B2(G116), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n769), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n713), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G137), .A2(new_n776), .B1(new_n710), .B2(G143), .ZN(new_n777));
  INV_X1    g0577(.A(G150), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n777), .B1(new_n778), .B2(new_n705), .C1(new_n721), .C2(new_n729), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT34), .Z(new_n780));
  NAND2_X1  g0580(.A1(new_n697), .A2(G132), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n285), .B1(new_n700), .B2(new_n202), .ZN(new_n782));
  INV_X1    g0582(.A(new_n701), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n782), .B1(new_n783), .B2(G58), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n781), .B(new_n784), .C1(new_n693), .C2(new_n301), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n775), .B1(new_n780), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n768), .B1(new_n786), .B2(new_n738), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(new_n750), .B2(new_n760), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n765), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(G384));
  AOI211_X1 g0590(.A(new_n491), .B(new_n213), .C1(new_n535), .C2(KEYINPUT35), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(KEYINPUT35), .B2(new_n535), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT36), .Z(new_n793));
  OR3_X1    g0593(.A1(new_n217), .A2(new_n214), .A3(new_n359), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n202), .A2(G68), .ZN(new_n795));
  AOI211_X1 g0595(.A(G13), .B(new_n268), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n394), .B1(new_n358), .B2(new_n374), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n393), .B1(new_n798), .B2(new_n401), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n620), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n417), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT38), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n402), .A2(new_n403), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n620), .B2(new_n799), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n799), .A2(new_n408), .ZN(new_n805));
  OAI21_X1  g0605(.A(KEYINPUT37), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n377), .A2(new_n411), .ZN(new_n807));
  INV_X1    g0607(.A(new_n620), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n377), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT37), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n807), .A2(new_n803), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n802), .B1(new_n806), .B2(new_n811), .ZN(new_n812));
  AND3_X1   g0612(.A1(new_n801), .A2(new_n812), .A3(KEYINPUT98), .ZN(new_n813));
  AOI21_X1  g0613(.A(KEYINPUT98), .B1(new_n801), .B2(new_n812), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n809), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT96), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n414), .A2(new_n415), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n413), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n817), .B1(new_n414), .B2(new_n415), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n816), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n807), .A2(new_n803), .A3(new_n809), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(KEYINPUT37), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n811), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n802), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n815), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(KEYINPUT40), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n346), .A2(new_n347), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n829), .A2(new_n342), .A3(new_n341), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT94), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n318), .A2(new_n625), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n832), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n341), .B(new_n834), .C1(new_n348), .C2(new_n318), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n831), .B1(new_n830), .B2(new_n832), .ZN(new_n837));
  OAI21_X1  g0637(.A(KEYINPUT95), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n830), .A2(new_n832), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(KEYINPUT94), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT95), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n840), .A2(new_n841), .A3(new_n835), .A4(new_n833), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n843), .A2(new_n674), .A3(new_n760), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n828), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT102), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n838), .A2(new_n842), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n674), .A2(new_n760), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n801), .A2(new_n812), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n806), .A2(new_n811), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT38), .B1(new_n801), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n843), .A2(KEYINPUT102), .A3(new_n674), .A4(new_n760), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n849), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT40), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n845), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n441), .B2(new_n674), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n854), .B1(new_n844), .B2(new_n846), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT40), .B1(new_n861), .B2(new_n856), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n441), .A2(new_n674), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n862), .A2(new_n863), .A3(new_n845), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n860), .A2(new_n635), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n609), .A2(new_n625), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT100), .ZN(new_n867));
  XOR2_X1   g0667(.A(KEYINPUT97), .B(KEYINPUT39), .Z(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(new_n825), .B2(new_n802), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT98), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n850), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n801), .A2(new_n812), .A3(KEYINPUT98), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n869), .A2(KEYINPUT99), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT39), .B1(new_n851), .B2(new_n853), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT99), .B1(new_n815), .B2(new_n869), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n867), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT99), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n871), .A2(new_n872), .ZN(new_n879));
  INV_X1    g0679(.A(new_n868), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n826), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n878), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n882), .A2(KEYINPUT100), .A3(new_n874), .A4(new_n873), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n866), .B1(new_n877), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n620), .B1(new_n409), .B2(new_n412), .ZN(new_n885));
  INV_X1    g0685(.A(new_n759), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n761), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n843), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n885), .B1(new_n888), .B2(new_n854), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT101), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n653), .A2(new_n891), .A3(new_n441), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n891), .B1(new_n653), .B2(new_n441), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n614), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n890), .B(new_n894), .ZN(new_n895));
  OAI22_X1  g0695(.A1(new_n865), .A2(new_n895), .B1(new_n268), .B2(new_n679), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n865), .A2(new_n895), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n797), .B1(new_n896), .B2(new_n897), .ZN(G367));
  INV_X1    g0698(.A(new_n752), .ZN(new_n899));
  INV_X1    g0699(.A(new_n420), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n899), .B1(new_n643), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n234), .A2(new_n744), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n741), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n625), .B1(new_n583), .B2(new_n584), .ZN(new_n904));
  INV_X1    g0704(.A(new_n592), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n600), .B2(new_n904), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n701), .A2(new_n301), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(G150), .B2(new_n710), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n776), .A2(G143), .ZN(new_n910));
  INV_X1    g0710(.A(new_n700), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n332), .B1(new_n911), .B2(G58), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n909), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(G50), .B2(new_n718), .ZN(new_n914));
  AOI22_X1  g0714(.A1(G137), .A2(new_n697), .B1(new_n772), .B2(G159), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n914), .B(new_n915), .C1(new_n217), .C2(new_n693), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n694), .A2(G97), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n697), .A2(G317), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n911), .A2(G116), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT46), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n285), .B1(new_n710), .B2(G303), .ZN(new_n921));
  XNOR2_X1  g0721(.A(KEYINPUT109), .B(G311), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n776), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(G294), .B2(new_n772), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n917), .A2(new_n918), .A3(new_n925), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n718), .A2(G283), .B1(G107), .B2(new_n783), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT108), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n916), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT47), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n738), .B1(new_n929), .B2(new_n930), .ZN(new_n932));
  OAI221_X1 g0732(.A(new_n903), .B1(new_n754), .B2(new_n907), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n597), .A2(new_n622), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n557), .B(new_n560), .C1(new_n541), .C2(new_n625), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n629), .A2(KEYINPUT106), .A3(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT44), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT106), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n628), .B2(new_n936), .ZN(new_n941));
  OR3_X1    g0741(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n939), .B1(new_n938), .B2(new_n941), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n628), .A2(new_n936), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT45), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n942), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT107), .ZN(new_n947));
  INV_X1    g0747(.A(new_n639), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n624), .B1(new_n632), .B2(new_n623), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(new_n638), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n677), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n942), .A2(new_n943), .A3(new_n639), .A4(new_n945), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n949), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n947), .B1(new_n946), .B2(new_n948), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n677), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n644), .B(KEYINPUT41), .Z(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n681), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n907), .A2(KEYINPUT43), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n624), .A2(new_n936), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT42), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n557), .B1(new_n616), .B2(new_n935), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n625), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n963), .A2(KEYINPUT103), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(KEYINPUT42), .B2(new_n962), .ZN(new_n967));
  AOI21_X1  g0767(.A(KEYINPUT103), .B1(new_n963), .B2(new_n965), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n961), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n907), .A2(KEYINPUT43), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n969), .B(new_n970), .Z(new_n971));
  NAND2_X1  g0771(.A1(new_n948), .A2(new_n937), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT104), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT105), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n973), .A2(new_n974), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n971), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n933), .B1(new_n960), .B2(new_n979), .ZN(G387));
  NAND3_X1  g0780(.A1(new_n630), .A2(new_n631), .A3(new_n751), .ZN(new_n981));
  INV_X1    g0781(.A(new_n642), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n982), .A2(new_n747), .B1(G107), .B2(new_n207), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n418), .A2(G50), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT50), .ZN(new_n985));
  AOI21_X1  g0785(.A(G45), .B1(G68), .B2(G77), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n985), .A2(new_n982), .A3(new_n986), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n643), .B(new_n285), .C1(new_n231), .C2(G45), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n983), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n682), .B1(new_n989), .B2(new_n899), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n701), .A2(new_n420), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G159), .B2(new_n776), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n202), .B2(new_n709), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n705), .A2(new_n255), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n700), .A2(new_n217), .ZN(new_n995));
  NOR4_X1   g0795(.A1(new_n993), .A2(new_n332), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(G150), .A2(new_n697), .B1(new_n718), .B2(G68), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n917), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n332), .B1(new_n712), .B2(new_n696), .C1(new_n693), .C2(new_n491), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT110), .Z(new_n1000));
  INV_X1    g0800(.A(G283), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n701), .A2(new_n1001), .B1(new_n702), .B2(new_n700), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n772), .A2(new_n922), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G317), .A2(new_n710), .B1(new_n776), .B2(G322), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1003), .B(new_n1004), .C1(new_n721), .C2(new_n503), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT48), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1002), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n1006), .B2(new_n1005), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT49), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1000), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n998), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n990), .B1(new_n1012), .B2(new_n738), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n951), .A2(new_n681), .B1(new_n981), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n952), .A2(new_n644), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n677), .A2(new_n951), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(G393));
  NAND2_X1  g0817(.A1(new_n697), .A2(G322), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n285), .B1(new_n911), .B2(G283), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n720), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT111), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G311), .A2(new_n710), .B1(new_n776), .B2(G317), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT52), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n772), .A2(G303), .B1(G116), .B2(new_n783), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n702), .B2(new_n721), .ZN(new_n1025));
  NOR3_X1   g0825(.A1(new_n1021), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n701), .A2(new_n304), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n285), .B1(new_n700), .B2(new_n301), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G150), .A2(new_n776), .B1(new_n710), .B2(G159), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1027), .B(new_n1028), .C1(new_n1029), .C2(KEYINPUT51), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1029), .A2(KEYINPUT51), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G50), .B2(new_n772), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n418), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G143), .A2(new_n697), .B1(new_n718), .B2(new_n1033), .ZN(new_n1034));
  AND4_X1   g0834(.A1(new_n769), .A2(new_n1030), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n738), .B1(new_n1026), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n899), .B1(G97), .B2(new_n643), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n238), .A2(new_n744), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n741), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1036), .B(new_n1039), .C1(new_n754), .C2(new_n937), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n946), .A2(new_n948), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n954), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1040), .B1(new_n1042), .B2(new_n680), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n644), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n1042), .B2(new_n952), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1041), .A2(KEYINPUT107), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1046), .A2(new_n949), .A3(new_n953), .A4(new_n954), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1043), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(G390));
  INV_X1    g0849(.A(KEYINPUT115), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n888), .A2(new_n866), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n877), .A2(new_n883), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT113), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n886), .B1(new_n652), .B2(new_n758), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n843), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n866), .B(KEYINPUT112), .Z(new_n1056));
  NAND3_X1  g0856(.A1(new_n1055), .A2(new_n827), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1052), .A2(new_n1053), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(G330), .ZN(new_n1059));
  OR3_X1    g0859(.A1(new_n844), .A2(KEYINPUT114), .A3(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(KEYINPUT114), .B1(new_n844), .B2(new_n1059), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1058), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1053), .B1(new_n1052), .B2(new_n1057), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1050), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1052), .A2(new_n1057), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(KEYINPUT113), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1067), .A2(KEYINPUT115), .A3(new_n1062), .A4(new_n1058), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n676), .A2(new_n760), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1052), .B(new_n1057), .C1(new_n847), .C2(new_n1069), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n674), .A2(G330), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n441), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n614), .B(new_n1072), .C1(new_n892), .C2(new_n893), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1069), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1074), .A2(new_n843), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n887), .B1(new_n1062), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1054), .B1(new_n1074), .B2(new_n843), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1071), .A2(KEYINPUT116), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n762), .B1(new_n1071), .B2(KEYINPUT116), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n847), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1073), .B1(new_n1076), .B2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1065), .A2(new_n1068), .A3(new_n1070), .A4(new_n1082), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1083), .A2(new_n644), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1065), .A2(new_n1070), .A3(new_n1068), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT117), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1076), .A2(new_n1081), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1073), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AND3_X1   g0889(.A1(new_n1085), .A2(new_n1086), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1086), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1084), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n877), .A2(new_n749), .A3(new_n883), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n682), .B1(new_n767), .B2(new_n256), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n285), .B(new_n1027), .C1(G87), .C2(new_n911), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1095), .B1(new_n491), .B2(new_n709), .C1(new_n1001), .C2(new_n713), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(G294), .B2(new_n697), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G97), .A2(new_n718), .B1(new_n772), .B2(G107), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1097), .B(new_n1098), .C1(new_n301), .C2(new_n693), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n772), .A2(G137), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(KEYINPUT54), .B(G143), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1100), .B1(new_n729), .B2(new_n701), .C1(new_n721), .C2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT118), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n710), .A2(G132), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n776), .A2(G128), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n700), .A2(new_n778), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT53), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .A4(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n332), .B1(new_n697), .B2(G125), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n693), .B2(new_n202), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT119), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1099), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1094), .B1(new_n1112), .B2(new_n738), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1093), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n1085), .B2(new_n680), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1092), .A2(new_n1116), .ZN(G378));
  INV_X1    g0917(.A(new_n890), .ZN(new_n1118));
  XOR2_X1   g0918(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n261), .A2(new_n620), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT55), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n295), .A2(new_n299), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1123), .B1(new_n295), .B2(new_n299), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1120), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1126), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1128), .A2(new_n1119), .A3(new_n1124), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n859), .B2(G330), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1130), .ZN(new_n1132));
  NOR4_X1   g0932(.A1(new_n862), .A2(new_n1059), .A3(new_n845), .A4(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1118), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n857), .A2(new_n858), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n845), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(G330), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n1132), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n859), .A2(G330), .A3(new_n1130), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1138), .A2(new_n890), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT121), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1134), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1138), .A2(KEYINPUT121), .A3(new_n890), .A4(new_n1139), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n1142), .A2(KEYINPUT57), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1083), .A2(new_n1088), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1044), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1134), .A2(new_n1140), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT57), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1146), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1147), .A2(new_n681), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n682), .B1(new_n767), .B2(G50), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(G107), .A2(new_n710), .B1(new_n776), .B2(G116), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n320), .B2(new_n705), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n285), .A2(G41), .ZN(new_n1156));
  NOR4_X1   g0956(.A1(new_n1155), .A2(new_n908), .A3(new_n995), .A4(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(G283), .A2(new_n697), .B1(new_n718), .B2(new_n900), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(new_n726), .C2(new_n693), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(G41), .ZN(new_n1161));
  AOI21_X1  g0961(.A(G50), .B1(new_n280), .B2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1160), .A2(KEYINPUT58), .B1(new_n1156), .B2(new_n1162), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n706), .A2(G132), .B1(G125), .B2(new_n776), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1101), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n710), .A2(G128), .B1(new_n911), .B2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1164), .B(new_n1166), .C1(new_n778), .C2(new_n701), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G137), .B2(new_n718), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1170));
  AOI211_X1 g0970(.A(G33), .B(G41), .C1(new_n697), .C2(G124), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT59), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1171), .B1(new_n729), .B2(new_n693), .C1(new_n1168), .C2(new_n1172), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1163), .B1(KEYINPUT58), .B2(new_n1160), .C1(new_n1170), .C2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1153), .B1(new_n1174), .B2(new_n738), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n1130), .B2(new_n750), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1152), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1151), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(KEYINPUT122), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT122), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1151), .A2(new_n1180), .A3(new_n1177), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(G375));
  NOR2_X1   g0983(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1185), .A2(new_n959), .A3(new_n1089), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n847), .A2(new_n749), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT123), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n285), .B(new_n991), .C1(G97), .C2(new_n911), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n1001), .B2(new_n709), .C1(new_n702), .C2(new_n713), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G303), .B2(new_n697), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(G107), .A2(new_n718), .B1(new_n772), .B2(G116), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1191), .B(new_n1192), .C1(new_n304), .C2(new_n693), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n783), .A2(G50), .B1(new_n776), .B2(G132), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n710), .A2(G137), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n332), .B1(new_n911), .B2(G159), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n772), .B2(new_n1165), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(G128), .A2(new_n697), .B1(new_n718), .B2(G150), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(new_n693), .C2(new_n726), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1193), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n738), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n741), .B1(new_n301), .B2(new_n766), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1188), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1087), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1204), .B1(new_n1205), .B2(new_n680), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1186), .A2(new_n1207), .ZN(G381));
  OR4_X1    g1008(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n933), .B(new_n1048), .C1(new_n960), .C2(new_n979), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n1209), .A2(G378), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1182), .A2(new_n1211), .ZN(G407));
  NAND2_X1  g1012(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(KEYINPUT117), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1085), .A2(new_n1086), .A3(new_n1089), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1115), .B1(new_n1216), .B2(new_n1084), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1182), .A2(new_n1217), .ZN(new_n1218));
  OAI211_X1 g1018(.A(G213), .B(G407), .C1(new_n1218), .C2(G343), .ZN(G409));
  NAND3_X1  g1019(.A1(new_n1151), .A2(G378), .A3(new_n1177), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(KEYINPUT124), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT124), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1142), .A2(new_n1223), .A3(new_n1143), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1222), .A2(new_n681), .A3(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1145), .A2(new_n959), .A3(new_n1147), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1225), .A2(new_n1176), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n1217), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1220), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n621), .A2(G213), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1089), .A2(KEYINPUT60), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1044), .B1(new_n1233), .B2(new_n1184), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1185), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1207), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n789), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(G384), .A3(new_n1207), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1230), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(G2897), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1238), .A2(new_n1239), .A3(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1241), .ZN(new_n1243));
  AOI21_X1  g1043(.A(G384), .B1(new_n1236), .B2(new_n1207), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n789), .B(new_n1206), .C1(new_n1234), .C2(new_n1235), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1243), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1242), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT61), .B1(new_n1231), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT63), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1249), .B1(new_n1231), .B2(new_n1251), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(G393), .B(G396), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT125), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1210), .A2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n958), .B1(new_n1047), .B2(new_n677), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n976), .B(new_n978), .C1(new_n1258), .C2(new_n681), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1048), .B1(new_n1259), .B2(new_n933), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1255), .B1(new_n1257), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G387), .A2(G390), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1255), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1262), .A2(new_n1210), .A3(new_n1263), .A4(new_n1256), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1261), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1240), .B1(new_n1220), .B2(new_n1228), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(KEYINPUT63), .A3(new_n1250), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1248), .A2(new_n1252), .A3(new_n1266), .A4(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT62), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1267), .A2(new_n1270), .A3(new_n1250), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT61), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1242), .A2(new_n1246), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1272), .B1(new_n1267), .B2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1270), .B1(new_n1267), .B2(new_n1250), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(new_n1271), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1265), .B(KEYINPUT126), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1269), .B1(new_n1276), .B2(new_n1277), .ZN(G405));
  NAND2_X1  g1078(.A1(new_n1265), .A2(new_n1250), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1261), .A2(new_n1251), .A3(new_n1264), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT127), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1178), .A2(G378), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1282), .B1(new_n1218), .B2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(G378), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1283), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1285), .A2(KEYINPUT127), .A3(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1281), .B1(new_n1284), .B2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1218), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1289));
  OAI21_X1  g1089(.A(KEYINPUT127), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1289), .A2(new_n1290), .A3(new_n1280), .A4(new_n1279), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1288), .A2(new_n1291), .ZN(G402));
endmodule


