

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736;

  XNOR2_X1 U377 ( .A(n699), .B(n700), .ZN(n701) );
  NOR2_X1 U378 ( .A1(n625), .A2(n733), .ZN(n578) );
  NOR2_X1 U379 ( .A1(n637), .A2(n620), .ZN(n598) );
  BUF_X1 U380 ( .A(n560), .Z(n356) );
  NAND2_X1 U381 ( .A1(n568), .A2(n423), .ZN(n388) );
  OR2_X1 U382 ( .A1(n686), .A2(n606), .ZN(n393) );
  XNOR2_X1 U383 ( .A(n442), .B(n475), .ZN(n715) );
  XNOR2_X1 U384 ( .A(n395), .B(G116), .ZN(n458) );
  XNOR2_X1 U385 ( .A(n394), .B(KEYINPUT3), .ZN(n488) );
  INV_X1 U386 ( .A(KEYINPUT72), .ZN(n394) );
  NOR2_X4 U387 ( .A1(n570), .A2(n412), .ZN(n625) );
  NOR2_X1 U388 ( .A1(G953), .A2(G237), .ZN(n493) );
  XOR2_X1 U389 ( .A(G104), .B(G107), .Z(n505) );
  INV_X1 U390 ( .A(G953), .ZN(n710) );
  NOR2_X2 U391 ( .A1(n591), .A2(n579), .ZN(n580) );
  XNOR2_X2 U392 ( .A(n371), .B(n363), .ZN(n666) );
  XNOR2_X2 U393 ( .A(n388), .B(KEYINPUT0), .ZN(n592) );
  XNOR2_X2 U394 ( .A(n501), .B(n500), .ZN(n526) );
  NOR2_X2 U395 ( .A1(n662), .A2(n668), .ZN(n372) );
  NOR2_X1 U396 ( .A1(n502), .A2(n374), .ZN(n411) );
  INV_X1 U397 ( .A(n579), .ZN(n590) );
  INV_X1 U398 ( .A(KEYINPUT22), .ZN(n386) );
  XNOR2_X1 U399 ( .A(n583), .B(KEYINPUT35), .ZN(n584) );
  AND2_X1 U400 ( .A1(n359), .A2(n535), .ZN(n375) );
  NOR2_X1 U401 ( .A1(n576), .A2(n651), .ZN(n588) );
  XNOR2_X1 U402 ( .A(n387), .B(n386), .ZN(n576) );
  NOR2_X1 U403 ( .A1(n592), .A2(n419), .ZN(n387) );
  XNOR2_X1 U404 ( .A(n372), .B(n539), .ZN(n660) );
  XNOR2_X1 U405 ( .A(n381), .B(KEYINPUT106), .ZN(n540) );
  NAND2_X1 U406 ( .A1(n411), .A2(n590), .ZN(n410) );
  NAND2_X1 U407 ( .A1(n569), .A2(n420), .ZN(n419) );
  XNOR2_X1 U408 ( .A(n698), .B(n697), .ZN(n700) );
  XNOR2_X1 U409 ( .A(n393), .B(n361), .ZN(n554) );
  XNOR2_X1 U410 ( .A(n380), .B(n429), .ZN(n470) );
  NAND2_X1 U411 ( .A1(n391), .A2(n392), .ZN(n380) );
  XNOR2_X1 U412 ( .A(n720), .B(G101), .ZN(n487) );
  XNOR2_X1 U413 ( .A(n462), .B(n397), .ZN(n720) );
  XNOR2_X1 U414 ( .A(G113), .B(n441), .ZN(n475) );
  XOR2_X1 U415 ( .A(G902), .B(KEYINPUT15), .Z(n606) );
  XNOR2_X1 U416 ( .A(KEYINPUT10), .B(G140), .ZN(n429) );
  XNOR2_X1 U417 ( .A(KEYINPUT66), .B(KEYINPUT4), .ZN(n397) );
  XNOR2_X1 U418 ( .A(n357), .B(KEYINPUT19), .ZN(n560) );
  NOR2_X1 U419 ( .A1(n554), .A2(n374), .ZN(n357) );
  NAND2_X1 U420 ( .A1(n666), .A2(n665), .ZN(n662) );
  NOR2_X1 U421 ( .A1(n410), .A2(n409), .ZN(n408) );
  XNOR2_X1 U422 ( .A(n487), .B(n396), .ZN(n510) );
  OR2_X2 U423 ( .A1(n627), .A2(n663), .ZN(n533) );
  NOR2_X2 U424 ( .A1(n549), .A2(n634), .ZN(n663) );
  AND2_X1 U425 ( .A1(n571), .A2(n422), .ZN(n525) );
  NOR2_X2 U426 ( .A1(n645), .A2(n571), .ZN(n652) );
  NOR2_X1 U427 ( .A1(n370), .A2(n617), .ZN(n599) );
  XNOR2_X1 U428 ( .A(n470), .B(n421), .ZN(n474) );
  XNOR2_X1 U429 ( .A(n499), .B(KEYINPUT94), .ZN(n500) );
  NOR2_X1 U430 ( .A1(G902), .A2(n612), .ZN(n501) );
  XNOR2_X1 U431 ( .A(KEYINPUT71), .B(G469), .ZN(n407) );
  XNOR2_X1 U432 ( .A(KEYINPUT68), .B(G131), .ZN(n486) );
  AND2_X1 U433 ( .A1(n584), .A2(n585), .ZN(n368) );
  XNOR2_X1 U434 ( .A(n486), .B(G134), .ZN(n722) );
  XNOR2_X1 U435 ( .A(G137), .B(KEYINPUT69), .ZN(n503) );
  NAND2_X1 U436 ( .A1(n428), .A2(G146), .ZN(n391) );
  NOR2_X1 U437 ( .A1(n390), .A2(G953), .ZN(n389) );
  INV_X1 U438 ( .A(G224), .ZN(n390) );
  XNOR2_X1 U439 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n435) );
  XOR2_X1 U440 ( .A(KEYINPUT75), .B(KEYINPUT85), .Z(n436) );
  NAND2_X1 U441 ( .A1(n651), .A2(n652), .ZN(n591) );
  XNOR2_X1 U442 ( .A(n526), .B(KEYINPUT6), .ZN(n579) );
  XNOR2_X1 U443 ( .A(n510), .B(n414), .ZN(n612) );
  XNOR2_X1 U444 ( .A(n498), .B(n490), .ZN(n414) );
  XOR2_X1 U445 ( .A(G122), .B(G104), .Z(n441) );
  INV_X1 U446 ( .A(n410), .ZN(n551) );
  NAND2_X1 U447 ( .A1(n382), .A2(n528), .ZN(n381) );
  XNOR2_X1 U448 ( .A(n383), .B(n362), .ZN(n382) );
  BUF_X1 U449 ( .A(n526), .Z(n412) );
  XNOR2_X1 U450 ( .A(n482), .B(n481), .ZN(n483) );
  INV_X1 U451 ( .A(G475), .ZN(n481) );
  INV_X1 U452 ( .A(n592), .ZN(n595) );
  INV_X1 U453 ( .A(n412), .ZN(n413) );
  XNOR2_X1 U454 ( .A(n511), .B(n512), .ZN(n694) );
  NOR2_X1 U455 ( .A1(G952), .A2(n710), .ZN(n708) );
  INV_X1 U456 ( .A(KEYINPUT70), .ZN(n404) );
  INV_X1 U457 ( .A(KEYINPUT48), .ZN(n401) );
  INV_X1 U458 ( .A(G125), .ZN(n428) );
  XOR2_X1 U459 ( .A(G137), .B(G116), .Z(n489) );
  INV_X1 U460 ( .A(n645), .ZN(n420) );
  BUF_X1 U461 ( .A(n554), .Z(n371) );
  INV_X1 U462 ( .A(KEYINPUT80), .ZN(n559) );
  INV_X1 U463 ( .A(G107), .ZN(n395) );
  NAND2_X1 U464 ( .A1(n416), .A2(n400), .ZN(n600) );
  XNOR2_X1 U465 ( .A(G128), .B(KEYINPUT88), .ZN(n430) );
  XNOR2_X1 U466 ( .A(n431), .B(n366), .ZN(n432) );
  XNOR2_X1 U467 ( .A(KEYINPUT79), .B(KEYINPUT23), .ZN(n431) );
  XNOR2_X1 U468 ( .A(n367), .B(KEYINPUT24), .ZN(n366) );
  INV_X1 U469 ( .A(KEYINPUT87), .ZN(n367) );
  XNOR2_X1 U470 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n426) );
  XNOR2_X1 U471 ( .A(KEYINPUT99), .B(G134), .ZN(n464) );
  XNOR2_X1 U472 ( .A(n480), .B(n479), .ZN(n696) );
  XNOR2_X1 U473 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U474 ( .A(n474), .B(n473), .ZN(n480) );
  XNOR2_X1 U475 ( .A(n722), .B(G146), .ZN(n396) );
  XNOR2_X1 U476 ( .A(G140), .B(G110), .ZN(n504) );
  XNOR2_X1 U477 ( .A(n380), .B(n389), .ZN(n438) );
  XNOR2_X1 U478 ( .A(n619), .B(n524), .ZN(n549) );
  INV_X1 U479 ( .A(KEYINPUT101), .ZN(n524) );
  NAND2_X1 U480 ( .A1(n525), .A2(n634), .ZN(n502) );
  INV_X1 U481 ( .A(n529), .ZN(n409) );
  NOR2_X1 U482 ( .A1(n591), .A2(n413), .ZN(n657) );
  INV_X1 U483 ( .A(n371), .ZN(n529) );
  XNOR2_X1 U484 ( .A(n418), .B(n417), .ZN(n442) );
  XNOR2_X1 U485 ( .A(n440), .B(KEYINPUT16), .ZN(n417) );
  XNOR2_X1 U486 ( .A(n458), .B(n488), .ZN(n418) );
  XNOR2_X1 U487 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n373) );
  XNOR2_X1 U488 ( .A(n547), .B(n546), .ZN(n734) );
  NAND2_X1 U489 ( .A1(n595), .A2(n413), .ZN(n596) );
  NOR2_X1 U490 ( .A1(n589), .A2(n590), .ZN(n617) );
  XNOR2_X1 U491 ( .A(n692), .B(n376), .ZN(n695) );
  XNOR2_X1 U492 ( .A(n694), .B(n693), .ZN(n376) );
  INV_X1 U493 ( .A(n665), .ZN(n374) );
  AND2_X1 U494 ( .A1(n461), .A2(G221), .ZN(n358) );
  AND2_X1 U495 ( .A1(n640), .A2(n632), .ZN(n359) );
  XOR2_X1 U496 ( .A(n450), .B(n449), .Z(n360) );
  XOR2_X1 U497 ( .A(n445), .B(KEYINPUT77), .Z(n361) );
  XOR2_X1 U498 ( .A(KEYINPUT104), .B(n527), .Z(n362) );
  XOR2_X1 U499 ( .A(KEYINPUT38), .B(KEYINPUT73), .Z(n363) );
  XNOR2_X1 U500 ( .A(n470), .B(n503), .ZN(n721) );
  XOR2_X1 U501 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n364) );
  AND2_X1 U502 ( .A1(n585), .A2(KEYINPUT82), .ZN(n365) );
  XNOR2_X1 U503 ( .A(n440), .B(n430), .ZN(n433) );
  XNOR2_X2 U504 ( .A(G119), .B(G110), .ZN(n440) );
  OR2_X2 U505 ( .A1(n609), .A2(G902), .ZN(n384) );
  XNOR2_X1 U506 ( .A(n577), .B(KEYINPUT32), .ZN(n733) );
  XNOR2_X1 U507 ( .A(n541), .B(n373), .ZN(n736) );
  NOR2_X1 U508 ( .A1(n598), .A2(n663), .ZN(n370) );
  NAND2_X1 U509 ( .A1(n599), .A2(n368), .ZN(n398) );
  NAND2_X1 U510 ( .A1(n375), .A2(n536), .ZN(n379) );
  NAND2_X1 U511 ( .A1(n369), .A2(n582), .ZN(n583) );
  XNOR2_X1 U512 ( .A(n581), .B(KEYINPUT34), .ZN(n369) );
  NOR2_X2 U513 ( .A1(n694), .A2(G902), .ZN(n513) );
  NOR2_X4 U514 ( .A1(n538), .A2(n521), .ZN(n634) );
  XNOR2_X1 U515 ( .A(n434), .B(n358), .ZN(n385) );
  XNOR2_X1 U516 ( .A(n385), .B(n721), .ZN(n609) );
  XNOR2_X1 U517 ( .A(n467), .B(n468), .ZN(n704) );
  XOR2_X2 U518 ( .A(G478), .B(n469), .Z(n521) );
  XNOR2_X1 U519 ( .A(n715), .B(n443), .ZN(n686) );
  XNOR2_X1 U520 ( .A(n377), .B(n616), .ZN(G57) );
  NOR2_X2 U521 ( .A1(n615), .A2(n708), .ZN(n377) );
  XNOR2_X1 U522 ( .A(n378), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U523 ( .A1(n701), .A2(n708), .ZN(n378) );
  XNOR2_X1 U524 ( .A(n408), .B(KEYINPUT36), .ZN(n514) );
  XNOR2_X1 U525 ( .A(n379), .B(n404), .ZN(n403) );
  NAND2_X1 U526 ( .A1(n525), .A2(n526), .ZN(n383) );
  XNOR2_X2 U527 ( .A(n384), .B(n360), .ZN(n571) );
  NAND2_X1 U528 ( .A1(n427), .A2(G125), .ZN(n392) );
  XNOR2_X2 U529 ( .A(G128), .B(G143), .ZN(n462) );
  NAND2_X1 U530 ( .A1(n584), .A2(n585), .ZN(n586) );
  NAND2_X1 U531 ( .A1(n399), .A2(n398), .ZN(n400) );
  NAND2_X1 U532 ( .A1(n732), .A2(n599), .ZN(n399) );
  XNOR2_X1 U533 ( .A(n402), .B(n401), .ZN(n558) );
  NAND2_X1 U534 ( .A1(n405), .A2(n403), .ZN(n402) );
  XNOR2_X1 U535 ( .A(n406), .B(n364), .ZN(n405) );
  NAND2_X1 U536 ( .A1(n736), .A2(n734), .ZN(n406) );
  XNOR2_X2 U537 ( .A(n528), .B(KEYINPUT1), .ZN(n651) );
  XNOR2_X2 U538 ( .A(n513), .B(n407), .ZN(n528) );
  NOR2_X2 U539 ( .A1(n540), .A2(n356), .ZN(n627) );
  NOR2_X2 U540 ( .A1(n543), .A2(n542), .ZN(n545) );
  NAND2_X1 U541 ( .A1(n415), .A2(n586), .ZN(n416) );
  XNOR2_X1 U542 ( .A(n578), .B(n365), .ZN(n415) );
  XNOR2_X1 U543 ( .A(n689), .B(n424), .ZN(n690) );
  NOR2_X2 U544 ( .A1(n690), .A2(n708), .ZN(n691) );
  AND2_X1 U545 ( .A1(n493), .A2(G214), .ZN(n421) );
  NOR2_X1 U546 ( .A1(n516), .A2(n645), .ZN(n422) );
  AND2_X1 U547 ( .A1(n567), .A2(n566), .ZN(n423) );
  XOR2_X1 U548 ( .A(n688), .B(n687), .Z(n424) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U551 ( .A(n487), .B(n439), .ZN(n443) );
  INV_X1 U552 ( .A(KEYINPUT100), .ZN(n522) );
  XNOR2_X1 U553 ( .A(n704), .B(n703), .ZN(n705) );
  NAND2_X1 U554 ( .A1(G234), .A2(n710), .ZN(n425) );
  XNOR2_X1 U555 ( .A(n425), .B(n426), .ZN(n461) );
  INV_X1 U556 ( .A(G146), .ZN(n427) );
  XNOR2_X1 U557 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U558 ( .A(n436), .B(n435), .ZN(n437) );
  NOR2_X1 U559 ( .A1(G902), .A2(G237), .ZN(n444) );
  XOR2_X1 U560 ( .A(KEYINPUT74), .B(n444), .Z(n485) );
  NAND2_X1 U561 ( .A1(G210), .A2(n485), .ZN(n445) );
  XOR2_X1 U562 ( .A(KEYINPUT89), .B(KEYINPUT20), .Z(n448) );
  INV_X1 U563 ( .A(n606), .ZN(n446) );
  NAND2_X1 U564 ( .A1(G234), .A2(n446), .ZN(n447) );
  XNOR2_X1 U565 ( .A(n448), .B(n447), .ZN(n456) );
  NAND2_X1 U566 ( .A1(n456), .A2(G217), .ZN(n450) );
  XOR2_X1 U567 ( .A(KEYINPUT90), .B(KEYINPUT25), .Z(n449) );
  NAND2_X1 U568 ( .A1(G237), .A2(G234), .ZN(n451) );
  XNOR2_X1 U569 ( .A(n451), .B(KEYINPUT14), .ZN(n677) );
  OR2_X1 U570 ( .A1(n710), .A2(G902), .ZN(n452) );
  NAND2_X1 U571 ( .A1(n677), .A2(n452), .ZN(n454) );
  NOR2_X1 U572 ( .A1(G953), .A2(G952), .ZN(n453) );
  NOR2_X1 U573 ( .A1(n454), .A2(n453), .ZN(n562) );
  NAND2_X1 U574 ( .A1(G953), .A2(G900), .ZN(n455) );
  NAND2_X1 U575 ( .A1(n562), .A2(n455), .ZN(n516) );
  NAND2_X1 U576 ( .A1(n456), .A2(G221), .ZN(n457) );
  XNOR2_X1 U577 ( .A(n457), .B(KEYINPUT21), .ZN(n645) );
  XOR2_X1 U578 ( .A(n458), .B(G122), .Z(n460) );
  XNOR2_X1 U579 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n459) );
  XNOR2_X1 U580 ( .A(n460), .B(n459), .ZN(n468) );
  NAND2_X1 U581 ( .A1(n461), .A2(G217), .ZN(n466) );
  INV_X1 U582 ( .A(n462), .ZN(n463) );
  XNOR2_X1 U583 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U584 ( .A(n466), .B(n465), .ZN(n467) );
  NOR2_X1 U585 ( .A1(G902), .A2(n704), .ZN(n469) );
  XOR2_X1 U586 ( .A(KEYINPUT11), .B(KEYINPUT96), .Z(n472) );
  XNOR2_X1 U587 ( .A(G143), .B(KEYINPUT97), .ZN(n471) );
  XNOR2_X1 U588 ( .A(n472), .B(n471), .ZN(n473) );
  INV_X1 U589 ( .A(n475), .ZN(n478) );
  INV_X1 U590 ( .A(n486), .ZN(n476) );
  XNOR2_X1 U591 ( .A(n476), .B(KEYINPUT12), .ZN(n477) );
  NOR2_X1 U592 ( .A1(G902), .A2(n696), .ZN(n484) );
  XNOR2_X1 U593 ( .A(KEYINPUT13), .B(KEYINPUT98), .ZN(n482) );
  XNOR2_X2 U594 ( .A(n484), .B(n483), .ZN(n538) );
  NAND2_X1 U595 ( .A1(G214), .A2(n485), .ZN(n665) );
  XOR2_X1 U596 ( .A(KEYINPUT5), .B(KEYINPUT93), .Z(n492) );
  XNOR2_X1 U597 ( .A(G119), .B(G113), .ZN(n491) );
  XNOR2_X1 U598 ( .A(n492), .B(n491), .ZN(n497) );
  XOR2_X1 U599 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n495) );
  NAND2_X1 U600 ( .A1(G210), .A2(n493), .ZN(n494) );
  XNOR2_X1 U601 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U602 ( .A(n497), .B(n496), .ZN(n498) );
  INV_X1 U603 ( .A(G472), .ZN(n499) );
  INV_X1 U604 ( .A(n503), .ZN(n507) );
  XNOR2_X1 U605 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U606 ( .A(n507), .B(n506), .Z(n509) );
  NAND2_X1 U607 ( .A1(G227), .A2(n710), .ZN(n508) );
  XNOR2_X1 U608 ( .A(n509), .B(n508), .ZN(n512) );
  INV_X1 U609 ( .A(n510), .ZN(n511) );
  NAND2_X1 U610 ( .A1(n514), .A2(n651), .ZN(n640) );
  NAND2_X1 U611 ( .A1(n665), .A2(n526), .ZN(n515) );
  XOR2_X1 U612 ( .A(KEYINPUT30), .B(n515), .Z(n518) );
  NAND2_X1 U613 ( .A1(n528), .A2(n652), .ZN(n597) );
  NOR2_X1 U614 ( .A1(n516), .A2(n597), .ZN(n517) );
  NAND2_X1 U615 ( .A1(n518), .A2(n517), .ZN(n542) );
  INV_X1 U616 ( .A(n521), .ZN(n537) );
  NOR2_X1 U617 ( .A1(n537), .A2(n538), .ZN(n582) );
  INV_X1 U618 ( .A(n582), .ZN(n519) );
  NOR2_X1 U619 ( .A1(n542), .A2(n519), .ZN(n520) );
  NAND2_X1 U620 ( .A1(n529), .A2(n520), .ZN(n632) );
  NAND2_X1 U621 ( .A1(n521), .A2(n538), .ZN(n523) );
  XNOR2_X2 U622 ( .A(n523), .B(n522), .ZN(n619) );
  INV_X1 U623 ( .A(n663), .ZN(n530) );
  XOR2_X1 U624 ( .A(KEYINPUT28), .B(KEYINPUT105), .Z(n527) );
  NAND2_X1 U625 ( .A1(n530), .A2(n627), .ZN(n531) );
  NAND2_X1 U626 ( .A1(n531), .A2(KEYINPUT78), .ZN(n532) );
  XNOR2_X1 U627 ( .A(n532), .B(KEYINPUT47), .ZN(n536) );
  INV_X1 U628 ( .A(KEYINPUT78), .ZN(n534) );
  NAND2_X1 U629 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U630 ( .A1(n538), .A2(n537), .ZN(n668) );
  XNOR2_X1 U631 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n539) );
  NOR2_X1 U632 ( .A1(n660), .A2(n540), .ZN(n541) );
  INV_X1 U633 ( .A(n666), .ZN(n543) );
  XNOR2_X1 U634 ( .A(KEYINPUT81), .B(KEYINPUT39), .ZN(n544) );
  XNOR2_X1 U635 ( .A(n545), .B(n544), .ZN(n548) );
  NAND2_X1 U636 ( .A1(n548), .A2(n634), .ZN(n547) );
  XOR2_X1 U637 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n546) );
  NAND2_X1 U638 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U639 ( .A(KEYINPUT110), .B(n550), .Z(n735) );
  INV_X1 U640 ( .A(n651), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n551), .A2(n573), .ZN(n553) );
  XOR2_X1 U642 ( .A(KEYINPUT43), .B(KEYINPUT103), .Z(n552) );
  XNOR2_X1 U643 ( .A(n553), .B(n552), .ZN(n555) );
  NAND2_X1 U644 ( .A1(n555), .A2(n409), .ZN(n642) );
  INV_X1 U645 ( .A(n642), .ZN(n556) );
  NOR2_X1 U646 ( .A1(n735), .A2(n556), .ZN(n557) );
  AND2_X2 U647 ( .A1(n558), .A2(n557), .ZN(n602) );
  XNOR2_X2 U648 ( .A(n602), .B(n559), .ZN(n724) );
  NOR2_X1 U649 ( .A1(n724), .A2(KEYINPUT2), .ZN(n601) );
  INV_X1 U650 ( .A(n668), .ZN(n569) );
  INV_X1 U651 ( .A(n560), .ZN(n568) );
  NAND2_X1 U652 ( .A1(G953), .A2(G898), .ZN(n561) );
  NAND2_X1 U653 ( .A1(n562), .A2(n561), .ZN(n563) );
  NAND2_X1 U654 ( .A1(KEYINPUT86), .A2(n563), .ZN(n567) );
  NOR2_X1 U655 ( .A1(G898), .A2(n710), .ZN(n717) );
  NAND2_X1 U656 ( .A1(n677), .A2(n717), .ZN(n564) );
  NOR2_X1 U657 ( .A1(KEYINPUT86), .A2(n564), .ZN(n565) );
  NAND2_X1 U658 ( .A1(G902), .A2(n565), .ZN(n566) );
  NAND2_X1 U659 ( .A1(n588), .A2(n571), .ZN(n570) );
  XOR2_X1 U660 ( .A(KEYINPUT102), .B(n571), .Z(n587) );
  INV_X1 U661 ( .A(n587), .ZN(n646) );
  NAND2_X1 U662 ( .A1(n579), .A2(n646), .ZN(n572) );
  NOR2_X1 U663 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U664 ( .A(KEYINPUT76), .B(n574), .Z(n575) );
  NOR2_X1 U665 ( .A1(n576), .A2(n575), .ZN(n577) );
  INV_X1 U666 ( .A(KEYINPUT44), .ZN(n585) );
  XNOR2_X1 U667 ( .A(n580), .B(KEYINPUT33), .ZN(n672) );
  NOR2_X1 U668 ( .A1(n592), .A2(n672), .ZN(n581) );
  INV_X1 U669 ( .A(n584), .ZN(n732) );
  NAND2_X1 U670 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U671 ( .A(KEYINPUT95), .B(KEYINPUT31), .Z(n594) );
  NAND2_X1 U672 ( .A1(n657), .A2(n595), .ZN(n593) );
  XNOR2_X1 U673 ( .A(n594), .B(n593), .ZN(n637) );
  NOR2_X1 U674 ( .A1(n597), .A2(n596), .ZN(n620) );
  XNOR2_X2 U675 ( .A(n600), .B(KEYINPUT45), .ZN(n709) );
  NAND2_X1 U676 ( .A1(n601), .A2(n709), .ZN(n605) );
  NAND2_X1 U677 ( .A1(n602), .A2(n709), .ZN(n603) );
  NAND2_X1 U678 ( .A1(n603), .A2(KEYINPUT2), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n644) );
  NAND2_X1 U680 ( .A1(n644), .A2(n606), .ZN(n607) );
  XNOR2_X2 U681 ( .A(n607), .B(KEYINPUT65), .ZN(n702) );
  NAND2_X1 U682 ( .A1(n702), .A2(G217), .ZN(n608) );
  XNOR2_X1 U683 ( .A(n608), .B(n609), .ZN(n610) );
  NOR2_X2 U684 ( .A1(n610), .A2(n708), .ZN(n611) );
  XNOR2_X1 U685 ( .A(n611), .B(KEYINPUT126), .ZN(G66) );
  NAND2_X1 U686 ( .A1(n702), .A2(G472), .ZN(n614) );
  XNOR2_X1 U687 ( .A(n612), .B(KEYINPUT62), .ZN(n613) );
  XNOR2_X1 U688 ( .A(n614), .B(n613), .ZN(n615) );
  XOR2_X1 U689 ( .A(KEYINPUT63), .B(KEYINPUT84), .Z(n616) );
  XOR2_X1 U690 ( .A(G101), .B(n617), .Z(G3) );
  NAND2_X1 U691 ( .A1(n620), .A2(n634), .ZN(n618) );
  XNOR2_X1 U692 ( .A(n618), .B(G104), .ZN(G6) );
  XOR2_X1 U693 ( .A(KEYINPUT111), .B(KEYINPUT27), .Z(n622) );
  NAND2_X1 U694 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U695 ( .A(n622), .B(n621), .ZN(n624) );
  XOR2_X1 U696 ( .A(G107), .B(KEYINPUT26), .Z(n623) );
  XNOR2_X1 U697 ( .A(n624), .B(n623), .ZN(G9) );
  XOR2_X1 U698 ( .A(G110), .B(n625), .Z(n626) );
  XNOR2_X1 U699 ( .A(KEYINPUT112), .B(n626), .ZN(G12) );
  AND2_X1 U700 ( .A1(n627), .A2(n619), .ZN(n631) );
  XOR2_X1 U701 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n629) );
  XNOR2_X1 U702 ( .A(G128), .B(KEYINPUT114), .ZN(n628) );
  XNOR2_X1 U703 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U704 ( .A(n631), .B(n630), .ZN(G30) );
  XNOR2_X1 U705 ( .A(G143), .B(n632), .ZN(G45) );
  NAND2_X1 U706 ( .A1(n627), .A2(n634), .ZN(n633) );
  XNOR2_X1 U707 ( .A(n633), .B(G146), .ZN(G48) );
  XOR2_X1 U708 ( .A(G113), .B(KEYINPUT115), .Z(n636) );
  NAND2_X1 U709 ( .A1(n637), .A2(n634), .ZN(n635) );
  XNOR2_X1 U710 ( .A(n636), .B(n635), .ZN(G15) );
  NAND2_X1 U711 ( .A1(n619), .A2(n637), .ZN(n638) );
  XNOR2_X1 U712 ( .A(n638), .B(G116), .ZN(G18) );
  XOR2_X1 U713 ( .A(KEYINPUT116), .B(KEYINPUT37), .Z(n639) );
  XNOR2_X1 U714 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U715 ( .A(G125), .B(n641), .ZN(G27) );
  XNOR2_X1 U716 ( .A(G140), .B(n642), .ZN(G42) );
  XOR2_X1 U717 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n685) );
  NOR2_X1 U718 ( .A1(n660), .A2(n672), .ZN(n643) );
  NOR2_X1 U719 ( .A1(G953), .A2(n643), .ZN(n683) );
  BUF_X1 U720 ( .A(n644), .Z(n681) );
  XOR2_X1 U721 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n648) );
  NAND2_X1 U722 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U723 ( .A(n648), .B(n647), .ZN(n649) );
  NOR2_X1 U724 ( .A1(n649), .A2(n412), .ZN(n650) );
  XOR2_X1 U725 ( .A(KEYINPUT118), .B(n650), .Z(n655) );
  NOR2_X1 U726 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U727 ( .A(KEYINPUT50), .B(n653), .ZN(n654) );
  NOR2_X1 U728 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U729 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U730 ( .A(KEYINPUT51), .B(n658), .Z(n659) );
  NOR2_X1 U731 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U732 ( .A(KEYINPUT119), .B(n661), .Z(n675) );
  NOR2_X1 U733 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U734 ( .A(KEYINPUT121), .B(n664), .Z(n671) );
  NOR2_X1 U735 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U736 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U737 ( .A(KEYINPUT120), .B(n669), .ZN(n670) );
  NOR2_X1 U738 ( .A1(n671), .A2(n670), .ZN(n673) );
  NOR2_X1 U739 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U740 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U741 ( .A(KEYINPUT52), .B(n676), .ZN(n679) );
  NAND2_X1 U742 ( .A1(n677), .A2(G952), .ZN(n678) );
  NOR2_X1 U743 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U744 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U745 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U746 ( .A(n685), .B(n684), .ZN(G75) );
  NAND2_X1 U747 ( .A1(n702), .A2(G210), .ZN(n689) );
  XOR2_X1 U748 ( .A(KEYINPUT83), .B(KEYINPUT55), .Z(n688) );
  XNOR2_X1 U749 ( .A(n686), .B(KEYINPUT54), .ZN(n687) );
  XNOR2_X1 U750 ( .A(KEYINPUT56), .B(n691), .ZN(G51) );
  XOR2_X1 U751 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n693) );
  NAND2_X1 U752 ( .A1(n702), .A2(G469), .ZN(n692) );
  NOR2_X1 U753 ( .A1(n708), .A2(n695), .ZN(G54) );
  XNOR2_X1 U754 ( .A(KEYINPUT59), .B(KEYINPUT124), .ZN(n698) );
  XNOR2_X1 U755 ( .A(n696), .B(KEYINPUT123), .ZN(n697) );
  NAND2_X1 U756 ( .A1(n702), .A2(G475), .ZN(n699) );
  NAND2_X1 U757 ( .A1(n702), .A2(G478), .ZN(n706) );
  INV_X1 U758 ( .A(KEYINPUT125), .ZN(n703) );
  XNOR2_X1 U759 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U760 ( .A1(n708), .A2(n707), .ZN(G63) );
  NAND2_X1 U761 ( .A1(n710), .A2(n709), .ZN(n714) );
  NAND2_X1 U762 ( .A1(G953), .A2(G224), .ZN(n711) );
  XNOR2_X1 U763 ( .A(KEYINPUT61), .B(n711), .ZN(n712) );
  NAND2_X1 U764 ( .A1(n712), .A2(G898), .ZN(n713) );
  NAND2_X1 U765 ( .A1(n714), .A2(n713), .ZN(n719) );
  XOR2_X1 U766 ( .A(n715), .B(G101), .Z(n716) );
  NOR2_X1 U767 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U768 ( .A(n719), .B(n718), .ZN(G69) );
  XOR2_X1 U769 ( .A(n721), .B(n722), .Z(n723) );
  XNOR2_X1 U770 ( .A(n720), .B(n723), .ZN(n727) );
  XOR2_X1 U771 ( .A(n724), .B(n727), .Z(n725) );
  NOR2_X1 U772 ( .A1(G953), .A2(n725), .ZN(n726) );
  XNOR2_X1 U773 ( .A(n726), .B(KEYINPUT127), .ZN(n731) );
  XNOR2_X1 U774 ( .A(G227), .B(n727), .ZN(n728) );
  NAND2_X1 U775 ( .A1(n728), .A2(G900), .ZN(n729) );
  NAND2_X1 U776 ( .A1(n729), .A2(G953), .ZN(n730) );
  NAND2_X1 U777 ( .A1(n731), .A2(n730), .ZN(G72) );
  XNOR2_X1 U778 ( .A(n732), .B(G122), .ZN(G24) );
  XOR2_X1 U779 ( .A(G119), .B(n733), .Z(G21) );
  XNOR2_X1 U780 ( .A(n734), .B(G131), .ZN(G33) );
  XOR2_X1 U781 ( .A(G134), .B(n735), .Z(G36) );
  XNOR2_X1 U782 ( .A(n736), .B(G137), .ZN(G39) );
endmodule

