//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  INV_X1    g0012(.A(G50), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  OAI22_X1  g0016(.A1(new_n213), .A2(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT65), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n217), .B(new_n219), .C1(G77), .C2(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  INV_X1    g0022(.A(G116), .ZN(new_n223));
  INV_X1    g0023(.A(G270), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G257), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n202), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n230), .A2(new_n207), .ZN(new_n231));
  INV_X1    g0031(.A(G58), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(new_n215), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT64), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n212), .B(new_n229), .C1(new_n231), .C2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n224), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT66), .ZN(new_n248));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XOR2_X1   g0049(.A(G50), .B(G58), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  XOR2_X1   g0052(.A(KEYINPUT8), .B(G58), .Z(new_n253));
  NAND3_X1  g0053(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n230), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n258), .B1(new_n206), .B2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n256), .B1(new_n260), .B2(new_n253), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  OAI21_X1  g0063(.A(KEYINPUT76), .B1(new_n263), .B2(G33), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT77), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n265), .B1(new_n266), .B2(KEYINPUT3), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT76), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(new_n266), .A3(KEYINPUT3), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n263), .A2(KEYINPUT77), .A3(G33), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n264), .A2(new_n267), .A3(new_n269), .A4(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT7), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G20), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT3), .B(G33), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n272), .B1(new_n275), .B2(G20), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G68), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT75), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n279), .B1(new_n232), .B2(new_n215), .ZN(new_n280));
  NAND3_X1  g0080(.A1(KEYINPUT75), .A2(G58), .A3(G68), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(new_n233), .A3(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n282), .A2(G20), .B1(G159), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(KEYINPUT16), .B1(new_n278), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n263), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(KEYINPUT7), .B1(new_n288), .B2(new_n207), .ZN(new_n289));
  AOI211_X1 g0089(.A(new_n272), .B(G20), .C1(new_n286), .C2(new_n287), .ZN(new_n290));
  OAI21_X1  g0090(.A(G68), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(KEYINPUT16), .A3(new_n284), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n258), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n262), .B1(new_n285), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G41), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(G1), .A3(G13), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(G232), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT78), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G274), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT67), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  OR2_X1    g0102(.A1(G41), .A2(G45), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT67), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n303), .A2(new_n304), .A3(new_n206), .A4(G274), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n296), .A2(new_n297), .A3(KEYINPUT78), .A4(G232), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n300), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT79), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n300), .A2(new_n306), .A3(KEYINPUT79), .A4(new_n307), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OR2_X1    g0112(.A1(G223), .A2(G1698), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n214), .A2(G1698), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n286), .A2(new_n313), .A3(new_n287), .A4(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G33), .A2(G87), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n296), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n317), .A2(G179), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n308), .A2(new_n317), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n312), .A2(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n294), .A2(KEYINPUT18), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT81), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT81), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n294), .A2(new_n321), .A3(new_n324), .A4(KEYINPUT18), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT80), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n294), .A2(new_n321), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT18), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT82), .B(G190), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n315), .A2(new_n316), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n333), .B1(new_n334), .B2(new_n296), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n312), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT83), .ZN(new_n338));
  INV_X1    g0138(.A(G200), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n319), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT83), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n312), .A2(new_n341), .A3(new_n336), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n338), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n258), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n288), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n215), .B1(new_n276), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n282), .A2(G20), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n283), .A2(G159), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n344), .B1(new_n350), .B2(KEYINPUT16), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT16), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n215), .B1(new_n274), .B2(new_n276), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n352), .B1(new_n353), .B2(new_n349), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n261), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  XOR2_X1   g0155(.A(KEYINPUT84), .B(KEYINPUT17), .Z(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n343), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  AOI211_X1 g0158(.A(KEYINPUT83), .B(new_n335), .C1(new_n310), .C2(new_n311), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n341), .B1(new_n312), .B2(new_n336), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n294), .B1(new_n361), .B2(new_n340), .ZN(new_n362));
  NOR2_X1   g0162(.A1(KEYINPUT84), .A2(KEYINPUT17), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n358), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n312), .A2(new_n318), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n319), .A2(new_n320), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n329), .B1(new_n355), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT80), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(new_n323), .A3(new_n325), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n331), .A2(new_n364), .A3(new_n370), .ZN(new_n371));
  OR2_X1    g0171(.A1(KEYINPUT74), .A2(KEYINPUT14), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n266), .A2(new_n202), .ZN(new_n373));
  NOR2_X1   g0173(.A1(G226), .A2(G1698), .ZN(new_n374));
  INV_X1    g0174(.A(G232), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n374), .B1(new_n375), .B2(G1698), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n373), .B1(new_n376), .B2(new_n275), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n377), .A2(new_n296), .ZN(new_n378));
  XOR2_X1   g0178(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n296), .A2(new_n297), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G238), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n378), .A2(new_n380), .A3(new_n383), .A4(new_n306), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n383), .B(new_n306), .C1(new_n377), .C2(new_n296), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n385), .A2(KEYINPUT72), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT13), .B1(new_n385), .B2(KEYINPUT72), .ZN(new_n387));
  OAI211_X1 g0187(.A(G179), .B(new_n384), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n385), .A2(new_n379), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n390), .A2(G169), .B1(KEYINPUT74), .B2(KEYINPUT14), .ZN(new_n391));
  NAND2_X1  g0191(.A1(KEYINPUT74), .A2(KEYINPUT14), .ZN(new_n392));
  AOI211_X1 g0192(.A(new_n320), .B(new_n392), .C1(new_n384), .C2(new_n389), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n372), .B(new_n388), .C1(new_n391), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n207), .A2(G33), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n395), .B(KEYINPUT68), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n396), .A2(G77), .ZN(new_n397));
  INV_X1    g0197(.A(new_n283), .ZN(new_n398));
  OAI22_X1  g0198(.A1(new_n398), .A2(new_n213), .B1(new_n207), .B2(G68), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n258), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  XOR2_X1   g0200(.A(KEYINPUT73), .B(KEYINPUT11), .Z(new_n401));
  XNOR2_X1  g0201(.A(new_n400), .B(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n255), .A2(new_n215), .ZN(new_n403));
  XNOR2_X1  g0203(.A(new_n403), .B(KEYINPUT12), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n215), .B2(new_n260), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n394), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n390), .A2(G200), .ZN(new_n409));
  INV_X1    g0209(.A(G190), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n384), .B1(new_n386), .B2(new_n387), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n406), .B(new_n409), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n371), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n259), .A2(G50), .ZN(new_n415));
  INV_X1    g0215(.A(G150), .ZN(new_n416));
  NOR3_X1   g0216(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n416), .A2(new_n398), .B1(new_n417), .B2(new_n207), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n418), .B1(new_n396), .B2(new_n253), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n415), .B1(G50), .B2(new_n254), .C1(new_n419), .C2(new_n344), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT9), .ZN(new_n421));
  INV_X1    g0221(.A(G1698), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(G222), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G223), .A2(G1698), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n275), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n296), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n425), .B(new_n426), .C1(G77), .C2(new_n275), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n427), .B(new_n306), .C1(new_n214), .C2(new_n381), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n420), .A2(new_n421), .B1(new_n428), .B2(G200), .ZN(new_n429));
  OAI221_X1 g0229(.A(new_n429), .B1(new_n421), .B2(new_n420), .C1(new_n410), .C2(new_n428), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n430), .B(KEYINPUT10), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n428), .A2(G179), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(new_n320), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n420), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT70), .ZN(new_n435));
  NAND2_X1  g0235(.A1(G238), .A2(G1698), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n275), .B(new_n436), .C1(new_n375), .C2(G1698), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n437), .B(new_n426), .C1(G107), .C2(new_n275), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n382), .A2(G244), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(new_n306), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(G200), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n253), .A2(new_n283), .B1(G20), .B2(G77), .ZN(new_n443));
  XOR2_X1   g0243(.A(KEYINPUT15), .B(G87), .Z(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n443), .B1(new_n395), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G77), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n446), .A2(new_n258), .B1(new_n447), .B2(new_n255), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n259), .A2(G77), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT69), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n435), .B1(new_n442), .B2(new_n451), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n438), .A2(new_n306), .A3(new_n439), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G190), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n441), .A2(KEYINPUT70), .A3(new_n448), .A4(new_n450), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n452), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G179), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n440), .A2(new_n320), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(new_n451), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n431), .A2(new_n434), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n255), .A2(new_n203), .ZN(new_n464));
  XNOR2_X1  g0264(.A(new_n464), .B(KEYINPUT25), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n275), .A2(new_n207), .A3(G87), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT22), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n469));
  XNOR2_X1  g0269(.A(new_n469), .B(KEYINPUT88), .ZN(new_n470));
  NOR2_X1   g0270(.A1(KEYINPUT89), .A2(KEYINPUT23), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n207), .A2(G107), .ZN(new_n472));
  NAND2_X1  g0272(.A1(KEYINPUT89), .A2(KEYINPUT23), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR4_X1   g0274(.A1(new_n207), .A2(KEYINPUT89), .A3(KEYINPUT23), .A4(G107), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n275), .A2(KEYINPUT22), .A3(new_n207), .A4(G87), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n468), .A2(new_n470), .A3(new_n476), .A4(new_n477), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n478), .B(KEYINPUT24), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n465), .B1(new_n479), .B2(new_n258), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n222), .A2(new_n422), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n226), .A2(G1698), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n275), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  OR2_X1    g0283(.A1(KEYINPUT90), .A2(G294), .ZN(new_n484));
  NAND2_X1  g0284(.A1(KEYINPUT90), .A2(G294), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n484), .A2(G33), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n296), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(G45), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(G1), .ZN(new_n489));
  AND2_X1   g0289(.A1(KEYINPUT5), .A2(G41), .ZN(new_n490));
  NOR2_X1   g0290(.A1(KEYINPUT5), .A2(G41), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n492), .A2(G264), .A3(new_n296), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n489), .B(G274), .C1(new_n491), .C2(new_n490), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n487), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(new_n339), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(G190), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n206), .A2(G33), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n254), .A2(new_n500), .A3(new_n230), .A4(new_n257), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G107), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n480), .A2(new_n498), .A3(new_n499), .A4(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n444), .A2(new_n254), .ZN(new_n505));
  OAI221_X1 g0305(.A(KEYINPUT19), .B1(new_n204), .B2(G87), .C1(new_n373), .C2(G20), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n266), .A2(new_n202), .A3(G20), .ZN(new_n507));
  OR2_X1    g0307(.A1(new_n507), .A2(KEYINPUT19), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n275), .A2(new_n207), .A3(G68), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n505), .B1(new_n510), .B2(new_n258), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n445), .B2(new_n501), .ZN(new_n512));
  NOR2_X1   g0312(.A1(G238), .A2(G1698), .ZN(new_n513));
  INV_X1    g0313(.A(G244), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(G1698), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n515), .A2(new_n275), .B1(G33), .B2(G116), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(new_n296), .ZN(new_n517));
  OAI21_X1  g0317(.A(G250), .B1(new_n488), .B2(G1), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n489), .A2(G274), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n426), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n457), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n512), .B(new_n522), .C1(G169), .C2(new_n521), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n501), .A2(new_n221), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT86), .ZN(new_n525));
  XNOR2_X1  g0325(.A(new_n524), .B(new_n525), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n511), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(G200), .B1(new_n517), .B2(new_n520), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n521), .A2(G190), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n523), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n422), .A2(G257), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G264), .A2(G1698), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n275), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n534), .B(new_n426), .C1(G303), .C2(new_n275), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n492), .A2(G270), .A3(new_n296), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n535), .A2(new_n536), .A3(new_n494), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n502), .A2(G116), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n255), .A2(new_n223), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n257), .A2(new_n230), .B1(G20), .B2(new_n223), .ZN(new_n540));
  AOI21_X1  g0340(.A(G20), .B1(G33), .B2(G283), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(G33), .B2(new_n202), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n540), .A2(new_n542), .A3(KEYINPUT20), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT20), .B1(new_n540), .B2(new_n542), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n538), .B(new_n539), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n537), .A2(new_n545), .A3(G169), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT21), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT87), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT87), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n546), .A2(new_n550), .A3(new_n547), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n537), .A2(KEYINPUT21), .A3(G169), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n536), .A2(new_n494), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n553), .A2(G179), .A3(new_n535), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n549), .A2(new_n551), .B1(new_n555), .B2(new_n545), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n537), .A2(G200), .ZN(new_n557));
  INV_X1    g0357(.A(new_n545), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n557), .B(new_n558), .C1(new_n333), .C2(new_n537), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n504), .A2(new_n531), .A3(new_n556), .A4(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n501), .A2(new_n202), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n254), .A2(G97), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n277), .A2(G107), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n203), .A2(KEYINPUT6), .A3(G97), .ZN(new_n564));
  XOR2_X1   g0364(.A(G97), .B(G107), .Z(new_n565));
  OAI21_X1  g0365(.A(new_n564), .B1(new_n565), .B2(KEYINPUT6), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n566), .A2(G20), .B1(G77), .B2(new_n283), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  AOI211_X1 g0368(.A(new_n561), .B(new_n562), .C1(new_n568), .C2(new_n258), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n492), .A2(G257), .A3(new_n296), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n286), .A2(new_n287), .A3(G244), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT4), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n572), .A2(new_n573), .B1(G33), .B2(G283), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n275), .A2(KEYINPUT4), .A3(G244), .A4(new_n422), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n573), .B1(new_n275), .B2(G250), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n574), .B(new_n575), .C1(new_n422), .C2(new_n576), .ZN(new_n577));
  AOI211_X1 g0377(.A(new_n495), .B(new_n571), .C1(new_n577), .C2(new_n426), .ZN(new_n578));
  OAI21_X1  g0378(.A(KEYINPUT85), .B1(new_n578), .B2(new_n339), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n571), .B1(new_n577), .B2(new_n426), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n494), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT85), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n582), .A3(G200), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n578), .A2(G190), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n569), .A2(new_n579), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n562), .B1(new_n568), .B2(new_n258), .ZN(new_n586));
  INV_X1    g0386(.A(new_n561), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n578), .A2(new_n457), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n581), .A2(new_n320), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n468), .A2(new_n477), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n592), .A2(KEYINPUT24), .A3(new_n470), .A4(new_n476), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT24), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n478), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n258), .A3(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n465), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(new_n503), .A3(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n496), .A2(G169), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n457), .B2(new_n496), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n585), .A2(new_n591), .A3(new_n601), .ZN(new_n602));
  NOR4_X1   g0402(.A1(new_n414), .A2(new_n463), .A3(new_n560), .A4(new_n602), .ZN(G372));
  NOR2_X1   g0403(.A1(new_n414), .A2(new_n463), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n556), .A2(new_n601), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT92), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n585), .A2(new_n591), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n596), .A2(new_n499), .A3(new_n503), .A4(new_n597), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n608), .A2(new_n497), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n515), .A2(new_n275), .ZN(new_n610));
  NAND2_X1  g0410(.A1(G33), .A2(G116), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(KEYINPUT91), .A3(new_n426), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT91), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n516), .B2(new_n296), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n520), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n527), .B(new_n529), .C1(new_n339), .C2(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n512), .B(new_n522), .C1(G169), .C2(new_n616), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n609), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT92), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n556), .A2(new_n621), .A3(new_n601), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n606), .A2(new_n607), .A3(new_n620), .A4(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n523), .A2(new_n530), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT26), .B1(new_n591), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n618), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n619), .A2(new_n591), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT26), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n623), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n604), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n434), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n368), .A2(new_n322), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n460), .B(KEYINPUT93), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n635), .A2(new_n412), .B1(new_n407), .B2(new_n394), .ZN(new_n636));
  INV_X1    g0436(.A(new_n364), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n633), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n632), .B1(new_n638), .B2(new_n431), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n631), .A2(new_n639), .ZN(G369));
  INV_X1    g0440(.A(G13), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n641), .A2(G1), .A3(G20), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT27), .ZN(new_n643));
  OR3_X1    g0443(.A1(new_n642), .A2(KEYINPUT94), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(G213), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n645), .B1(new_n642), .B2(new_n643), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT94), .B1(new_n642), .B2(new_n643), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n644), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n648), .A2(KEYINPUT95), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(KEYINPUT95), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(G343), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n601), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n556), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n653), .A2(new_n558), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n555), .A2(new_n545), .ZN(new_n660));
  INV_X1    g0460(.A(new_n551), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n550), .B1(new_n546), .B2(new_n547), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n660), .B(new_n559), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n659), .B1(new_n663), .B2(new_n658), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n664), .A2(G330), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n556), .A2(new_n654), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n653), .B1(new_n480), .B2(new_n503), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n601), .B1(new_n668), .B2(new_n609), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n656), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n656), .B1(new_n667), .B2(new_n670), .ZN(G399));
  INV_X1    g0471(.A(new_n210), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(G41), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n204), .A2(G87), .A3(G116), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G1), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n234), .B2(new_n674), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT28), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n607), .A2(new_n605), .ZN(new_n679));
  INV_X1    g0479(.A(new_n620), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT96), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(KEYINPUT26), .B1(new_n619), .B2(new_n591), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT96), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n607), .A2(new_n620), .A3(new_n683), .A4(new_n605), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n591), .A2(new_n624), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n626), .B1(new_n685), .B2(new_n628), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n681), .A2(new_n682), .A3(new_n684), .A4(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n687), .A2(KEYINPUT29), .A3(new_n653), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n630), .A2(new_n653), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT29), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n663), .A2(new_n609), .A3(new_n624), .ZN(new_n692));
  INV_X1    g0492(.A(new_n602), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(new_n693), .A3(new_n653), .ZN(new_n694));
  INV_X1    g0494(.A(new_n496), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(new_n554), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n696), .A2(KEYINPUT30), .A3(new_n521), .A4(new_n580), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n616), .A2(G179), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n698), .A2(new_n581), .A3(new_n537), .A4(new_n695), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT30), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n580), .A2(new_n521), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n496), .A2(G179), .A3(new_n553), .A4(new_n535), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n697), .A2(new_n699), .A3(new_n703), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n704), .A2(KEYINPUT31), .A3(new_n654), .ZN(new_n705));
  AOI21_X1  g0505(.A(KEYINPUT31), .B1(new_n704), .B2(new_n654), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n694), .A2(new_n707), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n688), .A2(new_n691), .B1(G330), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n678), .B1(new_n709), .B2(G1), .ZN(G364));
  NAND2_X1  g0510(.A1(new_n457), .A2(new_n339), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT99), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n712), .A2(G20), .A3(new_n410), .ZN(new_n713));
  INV_X1    g0513(.A(G159), .ZN(new_n714));
  OAI21_X1  g0514(.A(KEYINPUT32), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n207), .A2(new_n457), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n332), .A2(new_n339), .A3(new_n716), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n712), .A2(G190), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n718), .A2(new_n207), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  OAI221_X1 g0520(.A(new_n715), .B1(new_n232), .B2(new_n717), .C1(new_n720), .C2(new_n202), .ZN(new_n721));
  INV_X1    g0521(.A(new_n716), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n722), .A2(new_n339), .A3(G190), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n721), .B1(G68), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n207), .A2(G179), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(G190), .A3(G200), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G87), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n725), .A2(new_n410), .A3(G200), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n203), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n713), .A2(KEYINPUT32), .A3(new_n714), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n332), .A2(G200), .A3(new_n716), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT98), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI211_X1 g0536(.A(new_n730), .B(new_n731), .C1(G50), .C2(new_n736), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n722), .A2(G190), .A3(G200), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n288), .B1(new_n738), .B2(G77), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n724), .A2(new_n728), .A3(new_n737), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n738), .A2(G311), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n484), .A2(new_n485), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n741), .B1(new_n720), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n743), .B1(G326), .B2(new_n736), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT100), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n275), .B1(new_n727), .B2(G303), .ZN(new_n746));
  INV_X1    g0546(.A(new_n729), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G283), .ZN(new_n748));
  INV_X1    g0548(.A(new_n713), .ZN(new_n749));
  INV_X1    g0549(.A(new_n717), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n749), .A2(G329), .B1(G322), .B2(new_n750), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n745), .A2(new_n746), .A3(new_n748), .A4(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n723), .ZN(new_n753));
  XOR2_X1   g0553(.A(KEYINPUT33), .B(G317), .Z(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n740), .B1(new_n752), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n230), .B1(G20), .B2(new_n320), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n757), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n251), .A2(G45), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n235), .A2(new_n488), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n672), .A2(new_n275), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G355), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n210), .A2(new_n275), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n765), .B1(G116), .B2(new_n210), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n756), .A2(new_n757), .B1(new_n761), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n641), .A2(G20), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G45), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n674), .A2(G1), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT97), .ZN(new_n773));
  INV_X1    g0573(.A(new_n760), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n769), .B(new_n773), .C1(new_n664), .C2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n772), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n665), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(G330), .B2(new_n664), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n775), .A2(new_n778), .ZN(G396));
  AOI22_X1  g0579(.A1(new_n736), .A2(G137), .B1(G159), .B2(new_n738), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(new_n416), .B2(new_n753), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(G143), .B2(new_n750), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT34), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(G50), .B2(new_n727), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n729), .A2(new_n215), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n288), .ZN(new_n786));
  INV_X1    g0586(.A(G132), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n784), .B(new_n786), .C1(new_n787), .C2(new_n713), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(G58), .B2(new_n719), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n719), .A2(G97), .B1(G116), .B2(new_n738), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n729), .A2(new_n221), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(new_n750), .B2(G294), .ZN(new_n792));
  INV_X1    g0592(.A(G283), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n792), .B1(new_n793), .B2(new_n753), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(G311), .B2(new_n749), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n275), .B1(new_n727), .B2(G107), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n790), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(G303), .B2(new_n736), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n757), .B1(new_n789), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n799), .A2(new_n773), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n757), .A2(new_n758), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n653), .B1(new_n448), .B2(new_n450), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n461), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n634), .A2(new_n803), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n800), .B1(G77), .B2(new_n802), .C1(new_n759), .C2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n689), .A2(new_n807), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n630), .A2(new_n462), .A3(new_n653), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n708), .A2(G330), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n814), .A2(new_n772), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n809), .A2(new_n816), .ZN(G384));
  OAI21_X1  g0617(.A(new_n352), .B1(new_n346), .B2(new_n349), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n261), .B1(new_n351), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n651), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n371), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n819), .B1(new_n367), .B2(new_n651), .ZN(new_n822));
  OAI21_X1  g0622(.A(KEYINPUT37), .B1(new_n362), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n343), .A2(new_n355), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT37), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n294), .A2(new_n652), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n824), .A2(new_n825), .A3(new_n328), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n821), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT38), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT104), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n371), .A2(new_n820), .B1(new_n827), .B2(new_n823), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(KEYINPUT38), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n831), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n833), .A2(KEYINPUT104), .A3(KEYINPUT38), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n835), .A2(KEYINPUT39), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n364), .A2(new_n633), .ZN(new_n838));
  INV_X1    g0638(.A(new_n826), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n824), .A2(new_n328), .A3(new_n826), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(KEYINPUT37), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n827), .ZN(new_n843));
  AOI21_X1  g0643(.A(KEYINPUT38), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(KEYINPUT38), .B2(new_n833), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT39), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n837), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n408), .A2(new_n654), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n633), .A2(new_n652), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n654), .A2(new_n460), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n811), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n394), .A2(new_n407), .A3(new_n654), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT102), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n394), .A2(KEYINPUT102), .A3(new_n407), .A4(new_n654), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n408), .B(new_n412), .C1(new_n406), .C2(new_n653), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n855), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT103), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n855), .A2(KEYINPUT103), .A3(new_n862), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n865), .A2(new_n836), .A3(new_n835), .A4(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n850), .A2(new_n852), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n688), .A2(new_n691), .A3(new_n604), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n639), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n868), .B(new_n870), .Z(new_n871));
  INV_X1    g0671(.A(KEYINPUT40), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n807), .B1(new_n860), .B2(new_n861), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n560), .A2(new_n602), .A3(new_n654), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n704), .A2(new_n654), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT31), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n704), .A2(KEYINPUT31), .A3(new_n654), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n874), .A2(new_n879), .A3(KEYINPUT105), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT105), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(new_n694), .B2(new_n707), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n873), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  NOR3_X1   g0683(.A1(new_n845), .A2(new_n872), .A3(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n883), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n835), .A2(new_n885), .A3(new_n836), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n884), .B1(new_n886), .B2(new_n872), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n604), .B1(new_n882), .B2(new_n880), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n887), .B(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(G330), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n871), .B(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n206), .B2(new_n770), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n566), .B(KEYINPUT101), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n223), .B1(new_n893), .B2(KEYINPUT35), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n894), .B(new_n231), .C1(KEYINPUT35), .C2(new_n893), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT36), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n280), .A2(new_n281), .ZN(new_n897));
  NOR3_X1   g0697(.A1(new_n897), .A2(new_n447), .A3(new_n234), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n215), .A2(G50), .ZN(new_n899));
  OAI211_X1 g0699(.A(G1), .B(new_n641), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n892), .A2(new_n896), .A3(new_n900), .ZN(G367));
  INV_X1    g0701(.A(G317), .ZN(new_n902));
  OAI22_X1  g0702(.A1(new_n720), .A2(new_n203), .B1(new_n902), .B2(new_n713), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(G311), .B2(new_n736), .ZN(new_n904));
  OAI22_X1  g0704(.A1(new_n753), .A2(new_n742), .B1(new_n729), .B2(new_n202), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n727), .A2(KEYINPUT46), .A3(G116), .ZN(new_n906));
  INV_X1    g0706(.A(new_n738), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n906), .B1(new_n907), .B2(new_n793), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n905), .A2(new_n908), .A3(new_n275), .ZN(new_n909));
  INV_X1    g0709(.A(G303), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n904), .B(new_n909), .C1(new_n910), .C2(new_n717), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT46), .B1(new_n727), .B2(G116), .ZN(new_n912));
  INV_X1    g0712(.A(G137), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n713), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n747), .A2(G77), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n416), .B2(new_n717), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n726), .A2(new_n232), .ZN(new_n917));
  AOI211_X1 g0717(.A(new_n916), .B(new_n917), .C1(new_n719), .C2(G68), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n738), .A2(G50), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n736), .A2(G143), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n288), .B1(new_n723), .B2(G159), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n918), .A2(new_n919), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n911), .A2(new_n912), .B1(new_n914), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT47), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n757), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n653), .A2(new_n527), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n626), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n619), .B2(new_n926), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n928), .A2(new_n774), .ZN(new_n929));
  INV_X1    g0729(.A(new_n764), .ZN(new_n930));
  OAI221_X1 g0730(.A(new_n761), .B1(new_n210), .B2(new_n445), .C1(new_n243), .C2(new_n930), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n925), .A2(new_n773), .A3(new_n929), .A4(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n670), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n933), .A2(new_n607), .A3(new_n605), .A4(new_n666), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n654), .A2(new_n588), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n607), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n591), .B1(new_n936), .B2(new_n601), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n934), .A2(KEYINPUT42), .B1(new_n653), .B2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT106), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n934), .B2(KEYINPUT42), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n928), .A2(KEYINPUT43), .ZN(new_n941));
  INV_X1    g0741(.A(new_n666), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n670), .A2(new_n679), .A3(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT42), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n943), .A2(KEYINPUT106), .A3(new_n944), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n938), .A2(new_n940), .A3(new_n941), .A4(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT107), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n943), .A2(KEYINPUT106), .A3(new_n944), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT106), .B1(new_n943), .B2(new_n944), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n951), .A2(KEYINPUT107), .A3(new_n941), .A4(new_n938), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n941), .B1(new_n951), .B2(new_n938), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n928), .A2(KEYINPUT43), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n665), .A2(new_n933), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n591), .A2(new_n653), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(new_n607), .B2(new_n935), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n953), .A2(new_n956), .A3(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n962), .B1(new_n953), .B2(new_n956), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n771), .A2(G1), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n667), .B(new_n933), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n709), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n655), .B1(new_n669), .B2(new_n666), .ZN(new_n970));
  AND3_X1   g0770(.A1(new_n960), .A2(KEYINPUT45), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT45), .B1(new_n960), .B2(new_n970), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n970), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT44), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n974), .A2(new_n975), .A3(new_n959), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT44), .B1(new_n960), .B2(new_n970), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n973), .A2(new_n978), .A3(new_n957), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n709), .B1(new_n969), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n673), .B(KEYINPUT41), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n967), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(KEYINPUT108), .B1(new_n966), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n953), .A2(new_n956), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n961), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n963), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT108), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n987), .A2(new_n988), .A3(new_n982), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n932), .B1(new_n984), .B2(new_n989), .ZN(G387));
  NAND2_X1  g0790(.A1(new_n968), .A2(new_n967), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n713), .A2(new_n416), .B1(new_n202), .B2(new_n729), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n726), .A2(new_n447), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n992), .A2(new_n288), .A3(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT109), .ZN(new_n995));
  INV_X1    g0795(.A(new_n736), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n996), .A2(new_n714), .B1(new_n213), .B2(new_n717), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n738), .A2(G68), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n719), .A2(new_n444), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n723), .A2(new_n253), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n736), .A2(G322), .B1(G311), .B2(new_n723), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n910), .B2(new_n907), .C1(new_n902), .C2(new_n717), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT48), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n793), .B2(new_n720), .C1(new_n742), .C2(new_n726), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT49), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n749), .A2(G326), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n747), .A2(G116), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1008), .A2(new_n288), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1002), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n1013), .A2(new_n757), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n761), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n764), .B1(new_n240), .B2(new_n488), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n675), .B2(new_n767), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n253), .A2(new_n213), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT50), .Z(new_n1019));
  NAND2_X1  g0819(.A1(G68), .A2(G77), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1019), .A2(new_n488), .A3(new_n1020), .A4(new_n675), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1017), .A2(new_n1021), .B1(new_n203), .B2(new_n672), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n773), .B1(new_n1015), .B2(new_n1022), .C1(new_n933), .C2(new_n774), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n673), .B(KEYINPUT110), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n969), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n709), .A2(new_n968), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n991), .B1(new_n1014), .B2(new_n1023), .C1(new_n1026), .C2(new_n1027), .ZN(G393));
  INV_X1    g0828(.A(new_n979), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n957), .B1(new_n973), .B2(new_n978), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n969), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1029), .A2(new_n709), .A3(new_n968), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1032), .A2(new_n1033), .A3(new_n1025), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1029), .A2(new_n967), .A3(new_n1030), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n736), .A2(G317), .B1(G311), .B2(new_n750), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT52), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n723), .A2(G303), .B1(G283), .B2(new_n727), .ZN(new_n1038));
  INV_X1    g0838(.A(G294), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1038), .B1(new_n1039), .B2(new_n907), .ZN(new_n1040));
  NOR4_X1   g0840(.A1(new_n1037), .A2(new_n275), .A3(new_n730), .A4(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n749), .A2(G322), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(new_n223), .C2(new_n720), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT111), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n720), .A2(new_n447), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n736), .A2(G150), .B1(G159), .B2(new_n750), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT51), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1045), .B(new_n1047), .C1(G50), .C2(new_n723), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n288), .B(new_n791), .C1(new_n749), .C2(G143), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(new_n215), .C2(new_n726), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n253), .B2(new_n738), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n757), .B1(new_n1044), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n959), .A2(new_n760), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n764), .A2(new_n247), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1054), .B(new_n761), .C1(new_n202), .C2(new_n210), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1052), .A2(new_n773), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1035), .A2(new_n1056), .ZN(new_n1057));
  AND3_X1   g0857(.A1(new_n1034), .A2(KEYINPUT112), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(KEYINPUT112), .B1(new_n1034), .B2(new_n1057), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(G390));
  INV_X1    g0861(.A(KEYINPUT114), .ZN(new_n1062));
  INV_X1    g0862(.A(G330), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n807), .A2(new_n1063), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n708), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1065), .A2(KEYINPUT113), .A3(new_n862), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT113), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n708), .A2(new_n1064), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n860), .A2(new_n861), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1064), .B1(new_n880), .B2(new_n882), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1066), .A2(new_n1070), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n687), .A2(new_n653), .A3(new_n808), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1073), .A2(new_n854), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n862), .B(new_n1064), .C1(new_n880), .C2(new_n882), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n862), .B2(new_n1065), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n855), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n869), .B(new_n639), .C1(new_n888), .C2(new_n1063), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n849), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n863), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n837), .A2(new_n1084), .A3(new_n847), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n845), .A2(new_n849), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n1074), .B2(new_n1069), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1066), .A2(new_n1070), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1076), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1062), .B(new_n1082), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1076), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1072), .A2(new_n1074), .B1(new_n855), .B2(new_n1077), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1062), .B1(new_n1095), .B2(new_n1080), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1094), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1091), .A2(new_n1025), .A3(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n837), .A2(new_n758), .A3(new_n847), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n773), .B1(new_n253), .B2(new_n802), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n736), .A2(G128), .B1(G50), .B2(new_n747), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n749), .A2(G125), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1103), .B(new_n1104), .C1(new_n787), .C2(new_n717), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n720), .A2(new_n714), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(KEYINPUT54), .B(G143), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n907), .A2(new_n1107), .ZN(new_n1108));
  NOR4_X1   g0908(.A1(new_n1105), .A2(new_n1106), .A3(new_n288), .A4(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n726), .A2(new_n416), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT53), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1109), .B(new_n1111), .C1(new_n913), .C2(new_n753), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT115), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n785), .B(new_n1045), .C1(G107), .C2(new_n723), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n728), .B1(new_n223), .B2(new_n717), .C1(new_n907), .C2(new_n202), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n275), .B(new_n1115), .C1(G294), .C2(new_n749), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1114), .B(new_n1116), .C1(new_n793), .C2(new_n996), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1102), .B1(new_n1118), .B2(new_n757), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1100), .A2(new_n967), .B1(new_n1101), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1099), .A2(new_n1120), .ZN(G378));
  NAND3_X1  g0921(.A1(new_n1094), .A2(new_n1097), .A3(new_n1079), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n1081), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n868), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n431), .A2(new_n434), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(KEYINPUT55), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT55), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n431), .A2(new_n1127), .A3(new_n434), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1129), .A2(new_n420), .A3(new_n652), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n652), .A2(new_n420), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1126), .A2(new_n1128), .A3(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1130), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1133), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n887), .A2(G330), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n886), .A2(new_n872), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n884), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1138), .A2(G330), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1136), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1124), .A2(new_n1137), .A3(new_n1142), .ZN(new_n1143));
  AND4_X1   g0943(.A1(G330), .A2(new_n1138), .A3(new_n1139), .A4(new_n1136), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1136), .B1(new_n887), .B2(G330), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n868), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1123), .A2(new_n1143), .A3(KEYINPUT57), .A4(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT118), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1142), .A2(new_n1148), .A3(new_n1137), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n1124), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n868), .A2(new_n1142), .A3(new_n1148), .A4(new_n1137), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1150), .A2(new_n1151), .B1(new_n1081), .B2(new_n1122), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1025), .B(new_n1147), .C1(new_n1152), .C2(KEYINPUT57), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1136), .A2(new_n758), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n719), .A2(G68), .B1(G116), .B2(new_n736), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT116), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n993), .B(new_n1156), .C1(G107), .C2(new_n750), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n275), .A2(G41), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1158), .B1(new_n729), .B2(new_n232), .C1(new_n445), .C2(new_n907), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G97), .B2(new_n723), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1157), .B(new_n1160), .C1(new_n793), .C2(new_n713), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT58), .Z(new_n1162));
  NOR2_X1   g0962(.A1(G33), .A2(G41), .ZN(new_n1163));
  OR3_X1    g0963(.A1(new_n1158), .A2(G50), .A3(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n753), .A2(new_n787), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n907), .A2(new_n913), .B1(new_n726), .B2(new_n1107), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1165), .B(new_n1166), .C1(new_n736), .C2(G125), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n416), .B2(new_n720), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(G128), .B2(new_n750), .ZN(new_n1169));
  XOR2_X1   g0969(.A(new_n1169), .B(KEYINPUT59), .Z(new_n1170));
  INV_X1    g0970(.A(G124), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1163), .B1(new_n714), .B2(new_n729), .C1(new_n713), .C2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1164), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n757), .B1(new_n1162), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n772), .B1(new_n213), .B2(new_n801), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1154), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1177), .B1(new_n1178), .B2(new_n967), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1153), .A2(new_n1179), .ZN(G375));
  NOR2_X1   g0980(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1182), .A2(new_n981), .A3(new_n1082), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n773), .B1(G68), .B2(new_n802), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1000), .B1(new_n793), .B2(new_n717), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT119), .Z(new_n1186));
  OAI221_X1 g0986(.A(new_n1186), .B1(new_n202), .B2(new_n726), .C1(new_n910), .C2(new_n713), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n915), .B1(new_n753), .B2(new_n223), .C1(new_n203), .C2(new_n907), .ZN(new_n1188));
  NOR3_X1   g0988(.A1(new_n1187), .A2(new_n275), .A3(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n1039), .B2(new_n996), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n719), .A2(G50), .B1(G150), .B2(new_n738), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT120), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1192), .B(new_n275), .C1(new_n787), .C2(new_n996), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G128), .B2(new_n749), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n727), .A2(G159), .B1(new_n747), .B2(G58), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1194), .B(new_n1195), .C1(new_n753), .C2(new_n1107), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n717), .A2(new_n913), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1190), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1184), .B1(new_n1198), .B2(new_n757), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT121), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1199), .B(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1069), .A2(new_n758), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1201), .A2(new_n1202), .B1(new_n967), .B2(new_n1079), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1183), .A2(new_n1203), .ZN(G381));
  INV_X1    g1004(.A(G384), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1205), .A2(new_n1183), .A3(new_n1203), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n868), .B1(new_n1207), .B2(new_n1148), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1151), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n967), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n1176), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1147), .A2(new_n1025), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1178), .A2(new_n1123), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT57), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1211), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(G378), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1060), .B(new_n932), .C1(new_n984), .C2(new_n989), .ZN(new_n1219));
  OR2_X1    g1019(.A1(G393), .A2(G396), .ZN(new_n1220));
  OR4_X1    g1020(.A1(new_n1206), .A2(new_n1218), .A3(new_n1219), .A4(new_n1220), .ZN(G407));
  OAI211_X1 g1021(.A(G407), .B(G213), .C1(G343), .C2(new_n1218), .ZN(G409));
  NOR2_X1   g1022(.A1(new_n645), .A2(G343), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G375), .B2(G378), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1095), .A2(KEYINPUT60), .A3(new_n1080), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n1025), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1082), .A2(KEYINPUT60), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1226), .B1(new_n1227), .B2(new_n1182), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n967), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1229), .B1(new_n1230), .B2(new_n1095), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1205), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1181), .B1(KEYINPUT60), .B2(new_n1082), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G384), .B(new_n1203), .C1(new_n1233), .C2(new_n1226), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n981), .B(new_n1123), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1143), .A2(new_n1146), .A3(new_n967), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1217), .A2(new_n1237), .A3(new_n1176), .A4(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1224), .A2(new_n1236), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(KEYINPUT62), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT61), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1223), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1243), .B(new_n1239), .C1(new_n1216), .C2(new_n1217), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1223), .A2(G2897), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n1235), .B2(KEYINPUT122), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1235), .A2(KEYINPUT122), .A3(new_n1245), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT122), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1247), .A2(new_n1248), .B1(new_n1236), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1244), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT62), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1224), .A2(new_n1252), .A3(new_n1236), .A4(new_n1239), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1241), .A2(new_n1242), .A3(new_n1251), .A4(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(G387), .A2(G390), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT124), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1255), .A2(new_n1256), .A3(new_n1219), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(G393), .B(G396), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT123), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1258), .B(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1257), .A2(new_n1261), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1260), .A2(new_n1256), .A3(new_n1255), .A4(new_n1219), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1262), .A2(KEYINPUT126), .A3(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT126), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1254), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT63), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(new_n1251), .B2(new_n1240), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1262), .A2(new_n1242), .A3(new_n1263), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1217), .B1(new_n1153), .B2(new_n1179), .ZN(new_n1271));
  AND4_X1   g1071(.A1(new_n1217), .A2(new_n1237), .A3(new_n1176), .A4(new_n1238), .ZN(new_n1272));
  NOR4_X1   g1072(.A1(new_n1271), .A2(new_n1272), .A3(new_n1235), .A4(new_n1223), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1270), .B1(new_n1273), .B2(KEYINPUT63), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1269), .A2(new_n1274), .A3(KEYINPUT125), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT125), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1245), .ZN(new_n1277));
  AOI211_X1 g1077(.A(new_n1249), .B(new_n1277), .C1(new_n1232), .C2(new_n1234), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n1246), .A2(new_n1278), .B1(KEYINPUT122), .B2(new_n1235), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(new_n1224), .B2(new_n1239), .ZN(new_n1280));
  OAI21_X1  g1080(.A(KEYINPUT63), .B1(new_n1280), .B2(new_n1273), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1262), .A2(new_n1242), .A3(new_n1263), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(new_n1240), .B2(new_n1268), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1276), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1267), .B1(new_n1275), .B2(new_n1284), .ZN(G405));
  OAI211_X1 g1085(.A(KEYINPUT127), .B(new_n1236), .C1(new_n1264), .C2(new_n1265), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1265), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1262), .A2(KEYINPUT126), .A3(new_n1263), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1236), .A2(KEYINPUT127), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1287), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1271), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1218), .A2(new_n1291), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1286), .A2(new_n1290), .A3(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1292), .B1(new_n1286), .B2(new_n1290), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(G402));
endmodule


