//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 1 0 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1334, new_n1335, new_n1336, new_n1337, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1412,
    new_n1413, new_n1415, new_n1416, new_n1417;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  AND2_X1   g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n202), .A2(G50), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G107), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n205), .B1(new_n217), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n208), .B1(new_n210), .B2(new_n211), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XOR2_X1   g0026(.A(G238), .B(G244), .Z(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT64), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  NAND3_X1  g0043(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(G1), .A2(G13), .ZN(new_n245));
  AND3_X1   g0045(.A1(new_n244), .A2(KEYINPUT67), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g0046(.A(KEYINPUT67), .B1(new_n244), .B2(new_n245), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT8), .B(G58), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(G20), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G150), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  OAI22_X1  g0055(.A1(new_n249), .A2(new_n252), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G20), .ZN(new_n257));
  INV_X1    g0057(.A(G50), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n257), .B1(new_n201), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n248), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n258), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n248), .A2(new_n263), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n261), .A2(G20), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(G50), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT9), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n271), .B1(new_n209), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n209), .A2(new_n272), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n274), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n277), .B1(G226), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT3), .B(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G222), .ZN(new_n285));
  OAI22_X1  g0085(.A1(new_n284), .A2(new_n285), .B1(new_n219), .B2(new_n282), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT3), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OR3_X1    g0090(.A1(new_n290), .A2(KEYINPUT66), .A3(new_n283), .ZN(new_n291));
  OAI21_X1  g0091(.A(KEYINPUT66), .B1(new_n290), .B2(new_n283), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n286), .B1(new_n293), .B2(G223), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n281), .B1(new_n294), .B2(new_n278), .ZN(new_n295));
  INV_X1    g0095(.A(G190), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(G200), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n270), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT10), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n270), .A2(new_n301), .A3(new_n297), .A4(new_n298), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n295), .A2(G179), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n295), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n304), .A2(new_n269), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(G20), .A2(G77), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT15), .B(G87), .ZN(new_n310));
  OAI221_X1 g0110(.A(new_n309), .B1(new_n249), .B2(new_n255), .C1(new_n252), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n248), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(G77), .B2(new_n262), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n266), .A2(G77), .A3(new_n267), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT69), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT69), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n266), .A2(new_n316), .A3(G77), .A4(new_n267), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n313), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n278), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n214), .B1(new_n291), .B2(new_n292), .ZN(new_n321));
  INV_X1    g0121(.A(G232), .ZN(new_n322));
  OAI22_X1  g0122(.A1(new_n284), .A2(new_n322), .B1(new_n221), .B2(new_n282), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n320), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G179), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n277), .B1(G244), .B2(new_n280), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n324), .A2(new_n326), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n305), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n319), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n324), .A2(G190), .A3(new_n326), .ZN(new_n331));
  INV_X1    g0131(.A(G200), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(new_n324), .B2(new_n326), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT68), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n331), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n324), .A2(KEYINPUT68), .A3(G190), .A4(new_n326), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n318), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n330), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n308), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n266), .A2(G68), .A3(new_n267), .ZN(new_n341));
  XOR2_X1   g0141(.A(new_n341), .B(KEYINPUT73), .Z(new_n342));
  OAI22_X1  g0142(.A1(new_n252), .A2(new_n219), .B1(new_n257), .B2(G68), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT72), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n343), .A2(new_n344), .B1(new_n258), .B2(new_n255), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n343), .A2(new_n344), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n248), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT11), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n263), .A2(new_n213), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT12), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n347), .A2(new_n348), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n342), .A2(new_n349), .A3(new_n351), .A4(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n276), .B1(new_n279), .B2(new_n214), .ZN(new_n355));
  NAND2_X1  g0155(.A1(G33), .A2(G97), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(G226), .A2(G1698), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n358), .B1(new_n322), .B2(G1698), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n357), .B1(new_n359), .B2(new_n282), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT70), .B1(new_n360), .B2(new_n278), .ZN(new_n361));
  INV_X1    g0161(.A(G226), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n283), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n322), .A2(G1698), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n288), .A2(new_n363), .A3(new_n289), .A4(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n356), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT70), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n367), .A3(new_n320), .ZN(new_n368));
  AOI211_X1 g0168(.A(KEYINPUT13), .B(new_n355), .C1(new_n361), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT71), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n361), .A2(new_n368), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT13), .ZN(new_n372));
  INV_X1    g0172(.A(new_n355), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT71), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n367), .B1(new_n366), .B2(new_n320), .ZN(new_n377));
  AOI211_X1 g0177(.A(KEYINPUT70), .B(new_n278), .C1(new_n365), .C2(new_n356), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n373), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT13), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n370), .A2(new_n376), .A3(G179), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n374), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT14), .B1(new_n382), .B2(G169), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT14), .ZN(new_n384));
  AOI211_X1 g0184(.A(new_n384), .B(new_n305), .C1(new_n380), .C2(new_n374), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n381), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT74), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g0188(.A(KEYINPUT74), .B(new_n381), .C1(new_n383), .C2(new_n385), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n354), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n370), .A2(new_n376), .A3(G190), .A4(new_n380), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n382), .A2(G200), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n354), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G58), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n396), .A2(new_n213), .ZN(new_n397));
  OAI21_X1  g0197(.A(G20), .B1(new_n397), .B2(new_n201), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n254), .A2(G159), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT75), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n287), .B2(G33), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n250), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(new_n288), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT7), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(new_n257), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G68), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n406), .B1(new_n405), .B2(new_n257), .ZN(new_n409));
  OAI211_X1 g0209(.A(KEYINPUT16), .B(new_n401), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT16), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n406), .B1(new_n282), .B2(G20), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n290), .A2(KEYINPUT7), .A3(new_n257), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n213), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n411), .B1(new_n414), .B2(new_n400), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n410), .A2(new_n415), .A3(new_n248), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G87), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n362), .A2(G1698), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(G223), .B2(G1698), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n417), .B1(new_n405), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n320), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n278), .A2(G232), .A3(new_n274), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n276), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(new_n296), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n276), .A2(new_n422), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n320), .B2(new_n420), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n424), .B1(new_n426), .B2(G200), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n249), .B1(new_n261), .B2(G20), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n266), .A2(new_n428), .B1(new_n263), .B2(new_n249), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n416), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT17), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT78), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n416), .A2(new_n427), .A3(KEYINPUT78), .A4(new_n429), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n432), .B1(new_n436), .B2(KEYINPUT17), .ZN(new_n437));
  NOR2_X1   g0237(.A1(G223), .A2(G1698), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n438), .B1(new_n362), .B2(G1698), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n439), .A2(new_n288), .A3(new_n403), .A4(new_n404), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n278), .B1(new_n440), .B2(new_n417), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n305), .B1(new_n441), .B2(new_n425), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT76), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n421), .A2(new_n443), .A3(new_n423), .A4(new_n325), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n443), .B1(new_n426), .B2(new_n325), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n416), .A2(new_n429), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT18), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT77), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT77), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n447), .A2(new_n448), .A3(new_n451), .A4(KEYINPUT18), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n447), .A2(new_n448), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT18), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n450), .A2(new_n452), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n437), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n340), .A2(new_n395), .A3(new_n458), .ZN(new_n459));
  XNOR2_X1  g0259(.A(G97), .B(G107), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT6), .ZN(new_n461));
  INV_X1    g0261(.A(G97), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n460), .A2(new_n461), .B1(new_n221), .B2(new_n463), .ZN(new_n464));
  OAI22_X1  g0264(.A1(new_n464), .A2(new_n257), .B1(new_n219), .B2(new_n255), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n221), .B1(new_n412), .B2(new_n413), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n248), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n261), .A2(G33), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n262), .B(new_n468), .C1(new_n246), .C2(new_n247), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G97), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n263), .A2(new_n462), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n467), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n220), .A2(G1698), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n403), .A2(new_n404), .A3(new_n474), .A4(new_n288), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT4), .ZN(new_n476));
  AND2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n288), .A2(new_n289), .A3(G250), .A4(G1698), .ZN(new_n478));
  AND2_X1   g0278(.A1(KEYINPUT4), .A2(G244), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n288), .A2(new_n289), .A3(new_n479), .A4(new_n283), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G283), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n320), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n261), .A2(G45), .ZN(new_n484));
  NOR2_X1   g0284(.A1(KEYINPUT5), .A2(G41), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n273), .ZN(new_n489));
  INV_X1    g0289(.A(G45), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(G1), .ZN(new_n491));
  INV_X1    g0291(.A(new_n487), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n491), .B1(new_n492), .B2(new_n485), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n278), .ZN(new_n494));
  INV_X1    g0294(.A(G257), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n489), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n483), .A2(new_n497), .A3(new_n325), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n475), .A2(new_n476), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n278), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n305), .B1(new_n501), .B2(new_n496), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n473), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT79), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT79), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n473), .A2(new_n505), .A3(new_n498), .A4(new_n502), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n467), .A2(new_n472), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n483), .A2(new_n497), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G200), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n499), .A2(new_n500), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n496), .B1(new_n510), .B2(new_n320), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G190), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n507), .A2(new_n509), .A3(new_n512), .A4(new_n471), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n504), .A2(new_n506), .A3(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n491), .A2(new_n216), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n278), .A2(new_n515), .B1(new_n273), .B2(new_n491), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G116), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n220), .A2(G1698), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(G238), .B2(G1698), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n518), .B1(new_n405), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n278), .B1(new_n521), .B2(KEYINPUT80), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT80), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n523), .B(new_n518), .C1(new_n405), .C2(new_n520), .ZN(new_n524));
  AOI211_X1 g0324(.A(G179), .B(new_n517), .C1(new_n522), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n521), .A2(KEYINPUT80), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n526), .A2(new_n320), .A3(new_n524), .ZN(new_n527));
  AOI21_X1  g0327(.A(G169), .B1(new_n527), .B2(new_n516), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT19), .ZN(new_n530));
  NOR2_X1   g0330(.A1(G97), .A2(G107), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n215), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n356), .A2(new_n257), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR4_X1   g0334(.A1(new_n250), .A2(new_n462), .A3(KEYINPUT19), .A4(G20), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n403), .A2(new_n404), .A3(new_n257), .A4(new_n288), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n534), .A2(new_n535), .B1(new_n536), .B2(new_n213), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n248), .ZN(new_n538));
  INV_X1    g0338(.A(new_n310), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(new_n262), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT81), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT81), .ZN(new_n543));
  AOI211_X1 g0343(.A(new_n543), .B(new_n540), .C1(new_n537), .C2(new_n248), .ZN(new_n544));
  OAI22_X1  g0344(.A1(new_n542), .A2(new_n544), .B1(new_n310), .B2(new_n469), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n529), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT82), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n470), .A2(G87), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n542), .B2(new_n544), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n517), .B1(new_n522), .B2(new_n524), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n550), .A2(new_n332), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n547), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n247), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n244), .A2(KEYINPUT67), .A3(new_n245), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n404), .A2(new_n288), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n556), .A2(new_n257), .A3(G68), .A4(new_n403), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n251), .A2(new_n530), .A3(G97), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n531), .A2(new_n215), .B1(new_n356), .B2(new_n257), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(new_n559), .B2(new_n530), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n555), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n543), .B1(new_n561), .B2(new_n540), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n538), .A2(KEYINPUT81), .A3(new_n541), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n562), .A2(new_n563), .B1(G87), .B2(new_n470), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n527), .A2(new_n516), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G200), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(KEYINPUT82), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n527), .A2(G190), .A3(new_n516), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n552), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n514), .A2(new_n546), .A3(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n288), .A2(new_n289), .A3(new_n257), .A4(G87), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT22), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n571), .A2(new_n572), .B1(G116), .B2(new_n251), .ZN(new_n573));
  OAI21_X1  g0373(.A(KEYINPUT85), .B1(new_n257), .B2(G107), .ZN(new_n574));
  XNOR2_X1  g0374(.A(new_n574), .B(KEYINPUT23), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n536), .A2(new_n572), .A3(new_n215), .ZN(new_n577));
  OAI21_X1  g0377(.A(KEYINPUT24), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n405), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n579), .A2(KEYINPUT22), .A3(new_n257), .A4(G87), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT24), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n580), .A2(new_n581), .A3(new_n575), .A4(new_n573), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n248), .ZN(new_n584));
  NAND2_X1  g0384(.A1(G33), .A2(G294), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n495), .A2(G1698), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(G250), .B2(G1698), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n585), .B1(new_n405), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT86), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT86), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n590), .B(new_n585), .C1(new_n405), .C2(new_n587), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n591), .A3(new_n320), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n494), .A2(new_n222), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n489), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G200), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n263), .A2(new_n221), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n597), .B(KEYINPUT25), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n469), .A2(new_n221), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n278), .B1(new_n588), .B2(KEYINPUT86), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n593), .B1(new_n601), .B2(new_n591), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(G190), .A3(new_n489), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n584), .A2(new_n596), .A3(new_n600), .A4(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n592), .A2(G179), .A3(new_n489), .A4(new_n594), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT87), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n305), .B1(new_n602), .B2(new_n489), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n555), .B1(new_n578), .B2(new_n582), .ZN(new_n609));
  INV_X1    g0409(.A(new_n600), .ZN(new_n610));
  OAI22_X1  g0410(.A1(new_n609), .A2(new_n610), .B1(new_n605), .B2(KEYINPUT87), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n604), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n493), .A2(G270), .A3(new_n278), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n489), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n222), .A2(G1698), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(G257), .B2(G1698), .ZN(new_n616));
  INV_X1    g0416(.A(G303), .ZN(new_n617));
  OAI22_X1  g0417(.A1(new_n405), .A2(new_n616), .B1(new_n617), .B2(new_n282), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n320), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G200), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n263), .A2(G116), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n469), .B2(G116), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n481), .B(new_n257), .C1(G33), .C2(new_n462), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT83), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT20), .ZN(new_n626));
  INV_X1    g0426(.A(G116), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n625), .A2(new_n626), .B1(new_n627), .B2(G20), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n244), .A2(new_n245), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n624), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(KEYINPUT83), .A2(KEYINPUT20), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n624), .A2(new_n628), .A3(new_n629), .A4(new_n631), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n623), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n614), .A2(new_n619), .A3(G190), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n621), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT84), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT84), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n621), .A2(new_n640), .A3(new_n636), .A4(new_n637), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT21), .ZN(new_n643));
  NOR2_X1   g0443(.A1(G257), .A2(G1698), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n644), .B1(new_n222), .B2(G1698), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n645), .A2(new_n288), .A3(new_n403), .A4(new_n404), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n290), .A2(G303), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n278), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n489), .A2(new_n613), .ZN(new_n649));
  OAI21_X1  g0449(.A(G169), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n643), .B1(new_n636), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n469), .A2(G116), .ZN(new_n652));
  INV_X1    g0452(.A(new_n622), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n633), .A2(new_n634), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n305), .B1(new_n614), .B2(new_n619), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(KEYINPUT21), .A3(new_n657), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n648), .A2(new_n649), .A3(new_n325), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n651), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n642), .A2(new_n661), .ZN(new_n662));
  NOR4_X1   g0462(.A1(new_n459), .A2(new_n570), .A3(new_n612), .A4(new_n662), .ZN(G372));
  INV_X1    g0463(.A(new_n459), .ZN(new_n664));
  INV_X1    g0464(.A(new_n546), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT88), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n565), .A2(new_n666), .A3(G200), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT88), .B1(new_n550), .B2(new_n332), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n564), .A2(new_n667), .A3(new_n668), .A4(new_n568), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n604), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n504), .A2(new_n506), .A3(new_n513), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n584), .A2(new_n600), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n605), .A2(KEYINPUT87), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n673), .B(new_n674), .C1(new_n607), .C2(new_n606), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n661), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n665), .B1(new_n672), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n504), .A2(new_n506), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n569), .A2(KEYINPUT26), .A3(new_n678), .A4(new_n546), .ZN(new_n679));
  INV_X1    g0479(.A(new_n503), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n669), .A2(new_n546), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT26), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n677), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n664), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n307), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n394), .A2(new_n330), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n437), .B1(new_n688), .B2(new_n390), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n455), .A2(new_n449), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n687), .B1(new_n691), .B2(new_n303), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n686), .A2(new_n692), .ZN(G369));
  OR2_X1    g0493(.A1(new_n662), .A2(KEYINPUT89), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n261), .A2(new_n257), .A3(G13), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n695), .A2(KEYINPUT27), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(KEYINPUT27), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G213), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(G343), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n636), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n662), .B2(KEYINPUT89), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n651), .A2(new_n658), .A3(new_n660), .ZN(new_n704));
  AOI22_X1  g0504(.A1(new_n694), .A2(new_n703), .B1(new_n704), .B2(new_n702), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT90), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n673), .A2(new_n700), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n675), .A2(new_n604), .A3(new_n707), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n708), .A2(KEYINPUT91), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(KEYINPUT91), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n675), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n700), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n706), .A2(G330), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n661), .A2(new_n700), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n709), .A2(new_n710), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n712), .A2(new_n701), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n715), .A2(new_n720), .ZN(G399));
  INV_X1    g0521(.A(new_n206), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G41), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n532), .A2(G116), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(G1), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n211), .B2(new_n724), .ZN(new_n727));
  XOR2_X1   g0527(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n728));
  XNOR2_X1  g0528(.A(new_n727), .B(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(G330), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n595), .A2(KEYINPUT94), .A3(new_n508), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT94), .B1(new_n595), .B2(new_n508), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n565), .A2(new_n325), .A3(new_n620), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n550), .A2(new_n602), .A3(new_n511), .A4(new_n659), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT93), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(KEYINPUT30), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n614), .A2(new_n619), .A3(G179), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n508), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n737), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n740), .A2(new_n550), .A3(new_n602), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  OAI211_X1 g0543(.A(KEYINPUT31), .B(new_n700), .C1(new_n734), .C2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n620), .A2(new_n325), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n550), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n511), .B1(new_n602), .B2(new_n489), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n747), .B1(new_n748), .B2(KEYINPUT94), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n742), .B(new_n738), .C1(new_n749), .C2(new_n731), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT31), .B1(new_n750), .B2(new_n700), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n745), .A2(new_n751), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n569), .A2(new_n546), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n612), .A2(new_n662), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n753), .A2(new_n754), .A3(new_n514), .A4(new_n701), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n730), .B1(new_n752), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n569), .A2(new_n678), .A3(new_n546), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n682), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n666), .B1(new_n565), .B2(G200), .ZN(new_n759));
  AOI211_X1 g0559(.A(KEYINPUT88), .B(new_n332), .C1(new_n527), .C2(new_n516), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n562), .A2(new_n563), .ZN(new_n762));
  AND3_X1   g0562(.A1(new_n762), .A2(new_n548), .A3(new_n568), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n761), .A2(new_n763), .B1(new_n545), .B2(new_n529), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT95), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n764), .A2(new_n765), .A3(KEYINPUT26), .A4(new_n680), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n669), .A2(new_n546), .A3(KEYINPUT26), .A4(new_n680), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(KEYINPUT95), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n758), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n700), .B1(new_n769), .B2(new_n677), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT96), .ZN(new_n771));
  AND3_X1   g0571(.A1(new_n770), .A2(new_n771), .A3(KEYINPUT29), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n771), .B1(new_n770), .B2(KEYINPUT29), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n685), .A2(new_n701), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT29), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n756), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n729), .B1(new_n778), .B2(G1), .ZN(G364));
  AND2_X1   g0579(.A1(new_n257), .A2(G13), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n261), .B1(new_n780), .B2(G45), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n724), .A2(KEYINPUT97), .A3(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT97), .ZN(new_n783));
  INV_X1    g0583(.A(new_n781), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n783), .B1(new_n784), .B2(new_n723), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n722), .A2(new_n290), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G355), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(G116), .B2(new_n206), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n239), .A2(G45), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n579), .A2(new_n722), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n211), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n793), .B1(new_n490), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n790), .B1(new_n791), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n209), .B1(new_n257), .B2(G169), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n797), .A2(KEYINPUT98), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(KEYINPUT98), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G13), .A2(G33), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n787), .B1(new_n796), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(G20), .A2(G179), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n807), .A2(new_n296), .A3(G200), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G322), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n325), .A2(new_n332), .A3(G190), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n811), .A2(G20), .ZN(new_n812));
  INV_X1    g0612(.A(G294), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n290), .B1(new_n809), .B2(new_n810), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(KEYINPUT100), .B1(new_n296), .B2(G20), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(G179), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n296), .A2(KEYINPUT100), .A3(G20), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(G200), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(G329), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n818), .A2(new_n332), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(G283), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n820), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n807), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(G200), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(G190), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(KEYINPUT33), .B(G317), .Z(new_n829));
  NOR2_X1   g0629(.A1(new_n826), .A2(new_n296), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G326), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n828), .A2(new_n829), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NOR3_X1   g0633(.A1(new_n807), .A2(G190), .A3(G200), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n834), .A2(KEYINPUT99), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n834), .A2(KEYINPUT99), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G311), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n325), .A2(G20), .A3(G190), .A4(G200), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT101), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n837), .A2(new_n838), .B1(new_n617), .B2(new_n840), .ZN(new_n841));
  OR4_X1    g0641(.A1(new_n814), .A2(new_n824), .A3(new_n833), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n819), .A2(G159), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT32), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n831), .A2(new_n258), .B1(new_n462), .B2(new_n812), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(G68), .B2(new_n827), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n821), .A2(G107), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n282), .B1(new_n215), .B2(new_n839), .C1(new_n809), .C2(new_n396), .ZN(new_n848));
  INV_X1    g0648(.A(new_n837), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n848), .B1(new_n849), .B2(G77), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n846), .A2(new_n847), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n842), .B1(new_n844), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n806), .B1(new_n852), .B2(new_n800), .ZN(new_n853));
  INV_X1    g0653(.A(new_n803), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n853), .B1(new_n706), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n706), .A2(G330), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n786), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n706), .A2(G330), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT102), .ZN(G396));
  AND3_X1   g0660(.A1(new_n319), .A2(new_n327), .A3(new_n329), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n701), .ZN(new_n862));
  INV_X1    g0662(.A(new_n338), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n863), .A2(new_n335), .B1(new_n319), .B2(new_n700), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n862), .B1(new_n864), .B2(new_n861), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n775), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n865), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n685), .A2(new_n701), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n866), .A2(new_n756), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n756), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n867), .B1(new_n685), .B2(new_n701), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n700), .B(new_n865), .C1(new_n677), .C2(new_n684), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n869), .A2(new_n873), .A3(new_n786), .ZN(new_n874));
  INV_X1    g0674(.A(new_n800), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n802), .ZN(new_n876));
  OAI22_X1  g0676(.A1(new_n837), .A2(new_n627), .B1(new_n221), .B2(new_n840), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n828), .A2(new_n823), .B1(new_n831), .B2(new_n617), .ZN(new_n878));
  OAI221_X1 g0678(.A(new_n290), .B1(new_n809), .B2(new_n813), .C1(new_n812), .C2(new_n462), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n819), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n880), .B1(new_n215), .B2(new_n822), .C1(new_n838), .C2(new_n881), .ZN(new_n882));
  XOR2_X1   g0682(.A(KEYINPUT103), .B(G143), .Z(new_n883));
  AOI22_X1  g0683(.A1(new_n830), .A2(G137), .B1(new_n808), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(G159), .ZN(new_n885));
  OAI221_X1 g0685(.A(new_n884), .B1(new_n253), .B2(new_n828), .C1(new_n837), .C2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT34), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  OAI221_X1 g0689(.A(new_n579), .B1(new_n396), .B2(new_n812), .C1(new_n840), .C2(new_n258), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(G132), .B2(new_n819), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n821), .A2(G68), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n889), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n882), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n894), .A2(KEYINPUT104), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n800), .B1(new_n894), .B2(KEYINPUT104), .ZN(new_n896));
  OAI221_X1 g0696(.A(new_n787), .B1(G77), .B2(new_n876), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT105), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n802), .B2(new_n867), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n874), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT106), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n874), .A2(new_n899), .A3(KEYINPUT106), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(G384));
  INV_X1    g0705(.A(new_n464), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT35), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n210), .A2(new_n627), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n906), .B2(KEYINPUT35), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT107), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n910), .B2(new_n909), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT36), .ZN(new_n913));
  OR3_X1    g0713(.A1(new_n211), .A2(new_n219), .A3(new_n397), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n258), .A2(G68), .ZN(new_n915));
  AOI211_X1 g0715(.A(new_n261), .B(G13), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n664), .B(new_n777), .C1(new_n772), .C2(new_n773), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n692), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n330), .A2(new_n700), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT108), .ZN(new_n921));
  INV_X1    g0721(.A(new_n389), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n372), .B1(new_n371), .B2(new_n373), .ZN(new_n923));
  OAI21_X1  g0723(.A(G169), .B1(new_n923), .B2(new_n369), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n384), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n382), .A2(KEYINPUT14), .A3(G169), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT74), .B1(new_n927), .B2(new_n381), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n353), .B1(new_n922), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n354), .A2(new_n701), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n929), .A2(new_n393), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n388), .A2(new_n389), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n353), .B(new_n700), .C1(new_n933), .C2(new_n394), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n868), .A2(new_n921), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n410), .A2(new_n248), .ZN(new_n936));
  INV_X1    g0736(.A(new_n409), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(G68), .A3(new_n407), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT16), .B1(new_n938), .B2(new_n401), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n429), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n698), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n457), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n448), .A2(new_n941), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT37), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n453), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n436), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n940), .B1(new_n447), .B2(new_n941), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n951), .A2(new_n434), .A3(new_n435), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT37), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n944), .A2(KEYINPUT38), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT38), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n942), .B1(new_n437), .B2(new_n456), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n949), .A2(new_n948), .B1(new_n952), .B2(KEYINPUT37), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n935), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT39), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n437), .A2(new_n690), .ZN(new_n963));
  INV_X1    g0763(.A(new_n945), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n453), .A2(new_n945), .A3(new_n430), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(KEYINPUT37), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(KEYINPUT109), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT109), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n966), .A2(new_n969), .A3(KEYINPUT37), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n968), .A2(new_n950), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT38), .B1(new_n965), .B2(new_n971), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n957), .A2(new_n958), .A3(new_n956), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n962), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n929), .A2(new_n700), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n955), .A2(new_n959), .A3(KEYINPUT39), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n455), .A2(new_n449), .A3(new_n698), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n961), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n919), .B(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n865), .B1(new_n752), .B2(new_n755), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n931), .B1(new_n929), .B2(new_n393), .ZN(new_n982));
  NOR3_X1   g0782(.A1(new_n390), .A2(new_n394), .A3(new_n930), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n972), .A2(new_n973), .ZN(new_n985));
  OAI21_X1  g0785(.A(KEYINPUT40), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n932), .A2(new_n934), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT40), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n960), .A2(new_n987), .A3(new_n988), .A4(new_n981), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n459), .B1(new_n755), .B2(new_n752), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n730), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n991), .B2(new_n990), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n980), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n261), .B2(new_n780), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n980), .A2(new_n993), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n917), .B1(new_n995), .B2(new_n996), .ZN(G367));
  OAI21_X1  g0797(.A(new_n804), .B1(new_n206), .B2(new_n310), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n793), .A2(new_n234), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n787), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n821), .A2(G97), .ZN(new_n1001));
  INV_X1    g0801(.A(G317), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1001), .B1(new_n881), .B2(new_n1002), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n828), .A2(new_n813), .B1(new_n831), .B2(new_n838), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n812), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1004), .B1(G107), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n579), .B1(G303), .B2(new_n808), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1006), .B(new_n1007), .C1(new_n823), .C2(new_n837), .ZN(new_n1008));
  OAI21_X1  g0808(.A(KEYINPUT46), .B1(new_n840), .B2(new_n627), .ZN(new_n1009));
  OR3_X1    g0809(.A1(new_n839), .A2(KEYINPUT46), .A3(new_n627), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1003), .B(new_n1008), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n822), .A2(new_n219), .ZN(new_n1012));
  INV_X1    g0812(.A(G137), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n881), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n837), .A2(new_n258), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n282), .B1(new_n396), .B2(new_n839), .C1(new_n828), .C2(new_n885), .ZN(new_n1016));
  NOR4_X1   g0816(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n830), .A2(new_n883), .B1(G150), .B2(new_n808), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1005), .A2(G68), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT114), .Z(new_n1021));
  AOI21_X1  g0821(.A(new_n1011), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1022), .A2(KEYINPUT47), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n875), .B1(new_n1022), .B2(KEYINPUT47), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1000), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n764), .B1(new_n564), .B2(new_n701), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n665), .A2(new_n549), .A3(new_n700), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1026), .A2(new_n803), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n473), .A2(new_n700), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n514), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n680), .A2(new_n700), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n719), .A2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1035), .B(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT113), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT44), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1034), .B1(KEYINPUT113), .B2(KEYINPUT44), .ZN(new_n1041));
  NOR3_X1   g0841(.A1(new_n720), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1040), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1041), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1043), .B1(new_n1044), .B2(new_n719), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n715), .B1(new_n1037), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1037), .A2(new_n1046), .A3(new_n715), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n717), .B1(new_n714), .B2(new_n716), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n856), .B(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n778), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n723), .B(KEYINPUT41), .Z(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n784), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT110), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n718), .A2(KEYINPUT42), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n719), .A2(new_n1033), .A3(new_n1058), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n709), .A2(new_n710), .A3(new_n1033), .A4(new_n716), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1060), .A2(KEYINPUT42), .B1(new_n678), .B2(new_n701), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1057), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1059), .A2(new_n1057), .A3(new_n1061), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT43), .Z(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(KEYINPUT111), .A3(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1066), .A2(KEYINPUT43), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1063), .A2(new_n1064), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(KEYINPUT111), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n1071), .A2(new_n1072), .B1(new_n715), .B2(new_n1034), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1072), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n715), .A2(new_n1034), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1074), .A2(new_n1075), .A3(new_n1070), .A4(new_n1068), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1029), .B1(new_n1056), .B2(new_n1077), .ZN(G387));
  NAND2_X1  g0878(.A1(new_n774), .A2(new_n777), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n870), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n1052), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1052), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n778), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n723), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n725), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1085), .A2(new_n788), .B1(new_n221), .B2(new_n722), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n231), .A2(new_n490), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n249), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n258), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT50), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n725), .B(new_n490), .C1(new_n213), .C2(new_n219), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n792), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1086), .B1(new_n1087), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n786), .B1(new_n1093), .B2(new_n804), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n812), .A2(new_n310), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(G159), .B2(new_n830), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n839), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G77), .A2(new_n1097), .B1(new_n808), .B2(G50), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1096), .A2(new_n1001), .A3(new_n579), .A4(new_n1098), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n837), .A2(new_n213), .B1(new_n249), .B2(new_n828), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT115), .Z(new_n1101));
  AOI211_X1 g0901(.A(new_n1099), .B(new_n1101), .C1(G150), .C2(new_n819), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n822), .A2(new_n627), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n405), .B1(new_n881), .B2(new_n832), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n827), .A2(G311), .B1(G317), .B2(new_n808), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1105), .B1(new_n810), .B2(new_n831), .C1(new_n837), .C2(new_n617), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT48), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1005), .A2(G283), .B1(G294), .B2(new_n1097), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n1103), .B(new_n1104), .C1(new_n1112), .C2(KEYINPUT49), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n1112), .A2(KEYINPUT49), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1102), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1094), .B1(new_n875), .B2(new_n1115), .C1(new_n714), .C2(new_n854), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1084), .B(new_n1116), .C1(new_n781), .C2(new_n1052), .ZN(G393));
  INV_X1    g0917(.A(KEYINPUT117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1049), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1119), .A2(new_n1047), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1080), .A2(new_n1052), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1118), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1050), .A2(KEYINPUT117), .A3(new_n1083), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n724), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1120), .A2(new_n784), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n804), .B1(new_n462), .B2(new_n206), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n242), .A2(new_n792), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n787), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n282), .B1(new_n1097), .B2(G283), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n847), .B(new_n1131), .C1(new_n881), .C2(new_n810), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT116), .Z(new_n1133));
  AOI22_X1  g0933(.A1(new_n830), .A2(G317), .B1(G311), .B2(new_n808), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT52), .Z(new_n1135));
  NAND2_X1  g0935(.A1(new_n849), .A2(G294), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1005), .A2(G116), .B1(new_n827), .B2(G303), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n830), .A2(G150), .B1(G159), .B2(new_n808), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT51), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n812), .A2(new_n219), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n579), .B1(new_n213), .B2(new_n839), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(G50), .C2(new_n827), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(G87), .A2(new_n821), .B1(new_n819), .B2(new_n883), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(new_n249), .C2(new_n837), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n1133), .A2(new_n1138), .B1(new_n1140), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1130), .B1(new_n1146), .B2(new_n800), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n1033), .B2(new_n854), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1127), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1126), .A2(new_n1150), .ZN(G390));
  NAND2_X1  g0951(.A1(new_n664), .A2(new_n756), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n918), .A2(new_n692), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n987), .A2(new_n756), .A3(new_n867), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n864), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n330), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n920), .B1(new_n770), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n700), .B1(new_n734), .B2(new_n743), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT31), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n744), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n704), .B1(new_n639), .B2(new_n641), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1162), .A2(new_n675), .A3(new_n604), .A4(new_n701), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n570), .A2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g0964(.A(G330), .B(new_n867), .C1(new_n1161), .C2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1165), .A2(new_n932), .A3(new_n934), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n1154), .A2(new_n1157), .A3(new_n1166), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1154), .A2(new_n1166), .B1(new_n868), .B2(new_n921), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1153), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1154), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n921), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n987), .B1(new_n872), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n975), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1173), .A2(new_n1174), .B1(new_n974), .B2(new_n976), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1174), .B1(new_n972), .B2(new_n973), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n757), .A2(new_n682), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n766), .A2(new_n768), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n677), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(new_n701), .A3(new_n1156), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n862), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1176), .B1(new_n1181), .B2(new_n987), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1171), .B1(new_n1175), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n970), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n969), .B1(new_n966), .B2(KEYINPUT37), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n947), .A2(new_n436), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n945), .B1(new_n437), .B2(new_n690), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n956), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT39), .B1(new_n1189), .B2(new_n955), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n955), .A2(KEYINPUT39), .A3(new_n959), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n935), .A2(new_n975), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n975), .B1(new_n1189), .B2(new_n955), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n987), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1193), .B1(new_n1157), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1192), .A2(new_n1195), .A3(new_n1154), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1183), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n724), .B1(new_n1170), .B2(new_n1197), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1192), .A2(new_n1195), .A3(new_n1154), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1154), .B1(new_n1192), .B2(new_n1195), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n918), .A2(new_n692), .A3(new_n1152), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1201), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1198), .A2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n801), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n787), .B1(new_n876), .B2(new_n1088), .ZN(new_n1208));
  INV_X1    g1008(.A(G132), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n282), .B1(new_n809), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(G128), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n828), .A2(new_n1013), .B1(new_n831), .B2(new_n1211), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1210), .B(new_n1212), .C1(G159), .C2(new_n1005), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(KEYINPUT54), .B(G143), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1097), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT53), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n839), .B2(new_n253), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n849), .A2(new_n1215), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n821), .A2(G50), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n819), .A2(G125), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1213), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n892), .B1(new_n881), .B2(new_n813), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT118), .Z(new_n1224));
  OAI22_X1  g1024(.A1(new_n837), .A2(new_n462), .B1(new_n215), .B2(new_n840), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n290), .B1(new_n809), .B2(new_n627), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n828), .A2(new_n221), .B1(new_n831), .B2(new_n823), .ZN(new_n1227));
  OR4_X1    g1027(.A1(new_n1141), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1222), .B1(new_n1224), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1208), .B1(new_n1229), .B2(new_n800), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1207), .A2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n1197), .B2(new_n781), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1206), .A2(new_n1233), .ZN(G378));
  NAND2_X1  g1034(.A1(new_n269), .A2(new_n941), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT55), .Z(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n303), .B2(new_n307), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  XOR2_X1   g1039(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n1240));
  NAND3_X1  g1040(.A1(new_n303), .A2(new_n307), .A3(new_n1237), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1240), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1236), .B(new_n687), .C1(new_n300), .C2(new_n302), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1243), .B1(new_n1238), .B2(new_n1244), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n990), .B2(G330), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n730), .B(new_n1246), .C1(new_n986), .C2(new_n989), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n979), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n867), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n932), .B2(new_n934), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1189), .A2(new_n955), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n988), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  AND4_X1   g1054(.A1(new_n988), .A2(new_n960), .A3(new_n987), .A4(new_n981), .ZN(new_n1255));
  OAI21_X1  g1055(.A(G330), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1246), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n979), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n990), .A2(G330), .A3(new_n1247), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1250), .A2(new_n1260), .A3(new_n784), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n787), .B1(new_n876), .B2(G50), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n396), .A2(new_n822), .B1(new_n881), .B2(new_n823), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n827), .A2(G97), .B1(new_n830), .B2(G116), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(new_n405), .A3(new_n1019), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n837), .A2(new_n310), .ZN(new_n1266));
  INV_X1    g1066(.A(G41), .ZN(new_n1267));
  OAI221_X1 g1067(.A(new_n1267), .B1(new_n219), .B2(new_n839), .C1(new_n809), .C2(new_n221), .ZN(new_n1268));
  NOR4_X1   g1068(.A1(new_n1263), .A2(new_n1265), .A3(new_n1266), .A4(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1267), .B1(new_n405), .B2(new_n250), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1269), .A2(KEYINPUT58), .B1(new_n258), .B2(new_n1270), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n1215), .A2(new_n1097), .B1(G128), .B2(new_n808), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n828), .B2(new_n1209), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1005), .A2(G150), .B1(new_n830), .B2(G125), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1274), .B(new_n1275), .C1(new_n1013), .C2(new_n837), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(KEYINPUT59), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n250), .B(new_n1267), .C1(new_n822), .C2(new_n885), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(G124), .B2(new_n819), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1276), .A2(KEYINPUT59), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  OAI221_X1 g1081(.A(new_n1271), .B1(KEYINPUT58), .B2(new_n1269), .C1(new_n1277), .C2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1262), .B1(new_n1282), .B2(new_n800), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n1246), .B2(new_n802), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1261), .A2(new_n1284), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1250), .A2(new_n1260), .A3(KEYINPUT57), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1153), .B1(new_n1197), .B2(new_n1203), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n724), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT57), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1202), .B1(new_n1201), .B2(new_n1204), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1250), .A2(new_n1260), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1289), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1285), .B1(new_n1288), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT120), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1285), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1250), .A2(new_n1260), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT57), .B1(new_n1297), .B2(new_n1287), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1250), .A2(new_n1260), .A3(KEYINPUT57), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n723), .B1(new_n1299), .B2(new_n1290), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1296), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(KEYINPUT120), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1295), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(G375));
  NAND2_X1  g1104(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT121), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1305), .B(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1307), .A2(new_n1055), .A3(new_n1170), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1194), .A2(new_n801), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n787), .B1(new_n876), .B2(G68), .ZN(new_n1310));
  OAI22_X1  g1110(.A1(new_n837), .A2(new_n221), .B1(new_n462), .B2(new_n840), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n290), .B1(new_n809), .B2(new_n823), .ZN(new_n1312));
  OAI22_X1  g1112(.A1(new_n828), .A2(new_n627), .B1(new_n831), .B2(new_n813), .ZN(new_n1313));
  OR4_X1    g1113(.A1(new_n1095), .A2(new_n1311), .A3(new_n1312), .A4(new_n1313), .ZN(new_n1314));
  OAI22_X1  g1114(.A1(new_n219), .A2(new_n822), .B1(new_n881), .B2(new_n617), .ZN(new_n1315));
  OAI22_X1  g1115(.A1(new_n828), .A2(new_n1214), .B1(new_n258), .B2(new_n812), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n831), .A2(new_n1209), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  OAI221_X1 g1118(.A(new_n1318), .B1(new_n396), .B2(new_n822), .C1(new_n1211), .C2(new_n881), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n405), .B1(G137), .B2(new_n808), .ZN(new_n1320));
  OAI221_X1 g1120(.A(new_n1320), .B1(new_n885), .B2(new_n840), .C1(new_n837), .C2(new_n253), .ZN(new_n1321));
  OAI22_X1  g1121(.A1(new_n1314), .A2(new_n1315), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1310), .B1(new_n1322), .B2(new_n800), .ZN(new_n1323));
  AOI22_X1  g1123(.A1(new_n1169), .A2(new_n784), .B1(new_n1309), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1308), .A2(new_n1324), .ZN(G381));
  INV_X1    g1125(.A(new_n1077), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1080), .B1(new_n1120), .B2(new_n1082), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n781), .B1(new_n1327), .B2(new_n1054), .ZN(new_n1328));
  AOI22_X1  g1128(.A1(new_n1326), .A2(new_n1328), .B1(new_n1028), .B2(new_n1025), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1149), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1330));
  NOR3_X1   g1130(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1329), .A2(new_n1330), .A3(new_n1331), .ZN(new_n1332));
  OR4_X1    g1132(.A1(G378), .A2(G375), .A3(new_n1332), .A4(G381), .ZN(G407));
  AOI21_X1  g1133(.A(new_n1232), .B1(new_n1198), .B2(new_n1205), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n699), .A2(G213), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1303), .A2(new_n1334), .A3(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(G407), .A2(G213), .A3(new_n1337), .ZN(G409));
  NAND4_X1  g1138(.A1(new_n1287), .A2(new_n1055), .A3(new_n1260), .A4(new_n1250), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1339), .A2(new_n1261), .A3(new_n1284), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT123), .ZN(new_n1341));
  AND3_X1   g1141(.A1(new_n1340), .A2(new_n1341), .A3(new_n1334), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1341), .B1(new_n1340), .B2(new_n1334), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  AOI21_X1  g1144(.A(KEYINPUT122), .B1(new_n1293), .B2(G378), .ZN(new_n1345));
  OAI211_X1 g1145(.A(G378), .B(new_n1296), .C1(new_n1298), .C2(new_n1300), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT122), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1344), .B1(new_n1345), .B2(new_n1348), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n904), .A2(KEYINPUT125), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT60), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n723), .B1(new_n1305), .B2(new_n1351), .ZN(new_n1352));
  XOR2_X1   g1152(.A(KEYINPUT124), .B(KEYINPUT60), .Z(new_n1353));
  OAI21_X1  g1153(.A(new_n1353), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1352), .B1(new_n1307), .B2(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n902), .A2(KEYINPUT125), .A3(new_n903), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1324), .A2(new_n1356), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1350), .B1(new_n1355), .B2(new_n1357), .ZN(new_n1358));
  AND2_X1   g1158(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1359), .A2(new_n1306), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1305), .A2(KEYINPUT121), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1360), .A2(new_n1361), .A3(new_n1354), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1352), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1362), .A2(new_n1363), .ZN(new_n1364));
  INV_X1    g1164(.A(new_n1357), .ZN(new_n1365));
  INV_X1    g1165(.A(new_n1350), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1364), .A2(new_n1365), .A3(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1358), .A2(new_n1367), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(new_n1349), .A2(new_n1335), .A3(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1369), .A2(KEYINPUT62), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1293), .A2(KEYINPUT122), .A3(G378), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1371), .A2(new_n1372), .ZN(new_n1373));
  AOI21_X1  g1173(.A(new_n1336), .B1(new_n1373), .B2(new_n1344), .ZN(new_n1374));
  INV_X1    g1174(.A(KEYINPUT62), .ZN(new_n1375));
  NAND3_X1  g1175(.A1(new_n1374), .A2(new_n1375), .A3(new_n1368), .ZN(new_n1376));
  XOR2_X1   g1176(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1377));
  AOI21_X1  g1177(.A(new_n1366), .B1(new_n1364), .B2(new_n1365), .ZN(new_n1378));
  AOI211_X1 g1178(.A(new_n1357), .B(new_n1350), .C1(new_n1362), .C2(new_n1363), .ZN(new_n1379));
  INV_X1    g1179(.A(G2897), .ZN(new_n1380));
  NOR2_X1   g1180(.A1(new_n1335), .A2(new_n1380), .ZN(new_n1381));
  NOR3_X1   g1181(.A1(new_n1378), .A2(new_n1379), .A3(new_n1381), .ZN(new_n1382));
  INV_X1    g1182(.A(new_n1381), .ZN(new_n1383));
  AOI21_X1  g1183(.A(new_n1383), .B1(new_n1358), .B2(new_n1367), .ZN(new_n1384));
  NOR2_X1   g1184(.A1(new_n1382), .A2(new_n1384), .ZN(new_n1385));
  INV_X1    g1185(.A(new_n1385), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1340), .A2(new_n1334), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1387), .A2(KEYINPUT123), .ZN(new_n1388));
  NAND3_X1  g1188(.A1(new_n1340), .A2(new_n1341), .A3(new_n1334), .ZN(new_n1389));
  NAND2_X1  g1189(.A1(new_n1388), .A2(new_n1389), .ZN(new_n1390));
  AOI21_X1  g1190(.A(new_n1390), .B1(new_n1372), .B2(new_n1371), .ZN(new_n1391));
  OAI21_X1  g1191(.A(new_n1386), .B1(new_n1391), .B2(new_n1336), .ZN(new_n1392));
  NAND4_X1  g1192(.A1(new_n1370), .A2(new_n1376), .A3(new_n1377), .A4(new_n1392), .ZN(new_n1393));
  XNOR2_X1  g1193(.A(G393), .B(G396), .ZN(new_n1394));
  NOR2_X1   g1194(.A1(new_n1329), .A2(G390), .ZN(new_n1395));
  NOR2_X1   g1195(.A1(G387), .A2(new_n1330), .ZN(new_n1396));
  OAI21_X1  g1196(.A(new_n1394), .B1(new_n1395), .B2(new_n1396), .ZN(new_n1397));
  INV_X1    g1197(.A(new_n1394), .ZN(new_n1398));
  NAND2_X1  g1198(.A1(new_n1329), .A2(G390), .ZN(new_n1399));
  NAND2_X1  g1199(.A1(G387), .A2(new_n1330), .ZN(new_n1400));
  NAND3_X1  g1200(.A1(new_n1398), .A2(new_n1399), .A3(new_n1400), .ZN(new_n1401));
  NAND2_X1  g1201(.A1(new_n1397), .A2(new_n1401), .ZN(new_n1402));
  NAND2_X1  g1202(.A1(new_n1393), .A2(new_n1402), .ZN(new_n1403));
  INV_X1    g1203(.A(KEYINPUT61), .ZN(new_n1404));
  NAND3_X1  g1204(.A1(new_n1397), .A2(new_n1404), .A3(new_n1401), .ZN(new_n1405));
  AOI21_X1  g1205(.A(new_n1385), .B1(new_n1349), .B2(new_n1335), .ZN(new_n1406));
  INV_X1    g1206(.A(KEYINPUT126), .ZN(new_n1407));
  AOI21_X1  g1207(.A(new_n1405), .B1(new_n1406), .B2(new_n1407), .ZN(new_n1408));
  NAND2_X1  g1208(.A1(new_n1392), .A2(KEYINPUT126), .ZN(new_n1409));
  INV_X1    g1209(.A(KEYINPUT63), .ZN(new_n1410));
  NAND2_X1  g1210(.A1(new_n1369), .A2(new_n1410), .ZN(new_n1411));
  NAND3_X1  g1211(.A1(new_n1374), .A2(KEYINPUT63), .A3(new_n1368), .ZN(new_n1412));
  NAND4_X1  g1212(.A1(new_n1408), .A2(new_n1409), .A3(new_n1411), .A4(new_n1412), .ZN(new_n1413));
  NAND2_X1  g1213(.A1(new_n1403), .A2(new_n1413), .ZN(G405));
  NAND3_X1  g1214(.A1(new_n1295), .A2(new_n1334), .A3(new_n1302), .ZN(new_n1415));
  NAND2_X1  g1215(.A1(new_n1415), .A2(new_n1373), .ZN(new_n1416));
  XNOR2_X1  g1216(.A(new_n1416), .B(new_n1368), .ZN(new_n1417));
  XNOR2_X1  g1217(.A(new_n1417), .B(new_n1402), .ZN(G402));
endmodule


