//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n550,
    new_n552, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1222, new_n1223;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT66), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n460), .A2(G2105), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(G160));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  OR2_X1    g048(.A1(new_n473), .A2(G112), .ZN(new_n474));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n465), .A2(G136), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n478));
  NAND4_X1  g053(.A1(new_n461), .A2(new_n463), .A3(G124), .A4(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(KEYINPUT67), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G2104), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n481), .A2(new_n482), .A3(G124), .A4(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n477), .A2(new_n478), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n478), .B1(new_n477), .B2(new_n484), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(G162));
  NAND3_X1  g062(.A1(new_n481), .A2(G138), .A3(new_n473), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT4), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n461), .A2(new_n463), .A3(G126), .A4(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n489), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  XNOR2_X1  g070(.A(KEYINPUT5), .B(G543), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n496), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n497));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n496), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n499), .A2(new_n504), .ZN(G166));
  OR2_X1    g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(KEYINPUT69), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n509), .B1(new_n501), .B2(new_n502), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n508), .A2(new_n510), .A3(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT70), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n508), .A2(new_n510), .A3(new_n513), .A4(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n515), .A2(G51), .ZN(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT6), .B(G651), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n519), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n518), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n516), .A2(new_n524), .ZN(G168));
  NAND2_X1  g100(.A1(new_n515), .A2(G52), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n496), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n527), .A2(new_n498), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n522), .A2(new_n521), .B1(new_n501), .B2(new_n502), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G90), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n526), .A2(new_n528), .A3(new_n531), .ZN(G301));
  INV_X1    g107(.A(G301), .ZN(G171));
  INV_X1    g108(.A(G543), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n534), .B1(new_n519), .B2(new_n509), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n513), .B1(new_n535), .B2(new_n508), .ZN(new_n536));
  AND4_X1   g111(.A1(new_n513), .A2(new_n508), .A3(new_n510), .A4(G543), .ZN(new_n537));
  OAI21_X1  g112(.A(G43), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AND3_X1   g113(.A1(new_n496), .A2(new_n519), .A3(G81), .ZN(new_n539));
  OAI21_X1  g114(.A(G56), .B1(new_n521), .B2(new_n522), .ZN(new_n540));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT71), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n498), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n540), .A2(KEYINPUT71), .A3(new_n541), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n539), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n538), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT72), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n550), .A2(new_n554), .ZN(G188));
  NAND4_X1  g130(.A1(new_n508), .A2(new_n510), .A3(G53), .A4(G543), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT73), .ZN(new_n559));
  INV_X1    g134(.A(G91), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n529), .B2(new_n560), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n496), .A2(new_n519), .A3(KEYINPUT73), .A4(G91), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n564));
  AND2_X1   g139(.A1(G78), .A2(G543), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n565), .B1(new_n496), .B2(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n564), .B1(new_n566), .B2(new_n498), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n523), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g144(.A(KEYINPUT74), .B(G651), .C1(new_n569), .C2(new_n565), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n563), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n558), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G299));
  INV_X1    g148(.A(G168), .ZN(G286));
  INV_X1    g149(.A(G166), .ZN(G303));
  NAND3_X1  g150(.A1(new_n535), .A2(G49), .A3(new_n508), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n530), .A2(G87), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n496), .B2(G74), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G288));
  NAND3_X1  g154(.A1(new_n519), .A2(G48), .A3(G543), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n496), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n581), .B2(new_n498), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n530), .A2(G86), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G305));
  INV_X1    g160(.A(KEYINPUT75), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n515), .A2(G47), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n496), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G85), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n588), .A2(new_n498), .B1(new_n589), .B2(new_n529), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n586), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n590), .B1(new_n515), .B2(G47), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(KEYINPUT75), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n593), .ZN(G290));
  OAI21_X1  g169(.A(G54), .B1(new_n536), .B2(new_n537), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n529), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n496), .A2(new_n519), .A3(KEYINPUT10), .A4(G92), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n523), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n598), .A2(new_n599), .B1(G651), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n595), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G171), .B2(new_n605), .ZN(G284));
  OAI21_X1  g182(.A(new_n606), .B1(G171), .B2(new_n605), .ZN(G321));
  NAND2_X1  g183(.A1(G299), .A2(new_n605), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(new_n605), .B2(G168), .ZN(G280));
  XOR2_X1   g185(.A(G280), .B(KEYINPUT76), .Z(G297));
  INV_X1    g186(.A(new_n604), .ZN(new_n612));
  XNOR2_X1  g187(.A(KEYINPUT77), .B(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(G860), .B2(new_n613), .ZN(G148));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n548), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT78), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g194(.A1(new_n464), .A2(new_n473), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G123), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT80), .Z(new_n622));
  OR2_X1    g197(.A1(new_n473), .A2(G111), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  AOI22_X1  g200(.A1(new_n465), .A2(G135), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n465), .A2(G2104), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(G2100), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(G2100), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n628), .A2(new_n633), .A3(new_n634), .ZN(G156));
  XOR2_X1   g210(.A(KEYINPUT15), .B(G2435), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2427), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT81), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n637), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(KEYINPUT14), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n642), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(G14), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n647), .A2(new_n648), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT82), .Z(G401));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  AOI21_X1  g233(.A(KEYINPUT18), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  AOI21_X1  g235(.A(new_n660), .B1(new_n656), .B2(KEYINPUT18), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n659), .B(new_n661), .Z(new_n662));
  XOR2_X1   g237(.A(G2096), .B(G2100), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G227));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT19), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  AND2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT20), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n668), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n668), .B2(new_n674), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G229));
  INV_X1    g258(.A(G290), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G16), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G16), .B2(G24), .ZN(new_n686));
  INV_X1    g261(.A(G1986), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  INV_X1    g264(.A(G107), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n460), .B1(new_n690), .B2(G2105), .ZN(new_n691));
  INV_X1    g266(.A(G95), .ZN(new_n692));
  AND3_X1   g267(.A1(new_n692), .A2(new_n473), .A3(KEYINPUT83), .ZN(new_n693));
  AOI21_X1  g268(.A(KEYINPUT83), .B1(new_n692), .B2(new_n473), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n691), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n481), .A2(G131), .A3(new_n473), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n481), .A2(G119), .A3(G2105), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G25), .B(new_n698), .S(G29), .Z(new_n699));
  XOR2_X1   g274(.A(KEYINPUT35), .B(G1991), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n688), .A2(new_n689), .A3(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G6), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(new_n584), .B2(new_n703), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT84), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT32), .B(G1981), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(G16), .A2(G23), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT85), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G288), .B2(new_n703), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT33), .B(G1976), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n711), .B(new_n712), .Z(new_n713));
  NOR2_X1   g288(.A1(G16), .A2(G22), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G166), .B2(G16), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT86), .B(G1971), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n715), .B(new_n716), .Z(new_n717));
  NAND3_X1  g292(.A1(new_n708), .A2(new_n713), .A3(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(KEYINPUT34), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n702), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT87), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n718), .A2(KEYINPUT34), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT88), .B(KEYINPUT36), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n722), .A2(new_n724), .A3(new_n726), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT31), .B(G11), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT30), .B(G28), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n731), .B(new_n734), .C1(new_n627), .C2(new_n733), .ZN(new_n735));
  NOR2_X1   g310(.A1(G168), .A2(new_n703), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n703), .B2(G21), .ZN(new_n737));
  INV_X1    g312(.A(G1966), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n735), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G1961), .ZN(new_n740));
  NOR2_X1   g315(.A1(G171), .A2(new_n703), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G5), .B2(new_n703), .ZN(new_n742));
  OAI221_X1 g317(.A(new_n739), .B1(new_n740), .B2(new_n742), .C1(new_n738), .C2(new_n737), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT94), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n465), .A2(G139), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT89), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT25), .Z(new_n748));
  AOI22_X1  g323(.A1(new_n481), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(new_n473), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n751), .A2(new_n733), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n733), .B2(G33), .ZN(new_n753));
  INV_X1    g328(.A(G2072), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n733), .A2(G26), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT28), .Z(new_n757));
  NAND3_X1  g332(.A1(new_n481), .A2(G140), .A3(new_n473), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n481), .A2(G128), .A3(G2105), .ZN(new_n759));
  OR2_X1    g334(.A1(G104), .A2(G2105), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n760), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n757), .B1(new_n762), .B2(G29), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G2067), .ZN(new_n764));
  NOR2_X1   g339(.A1(G164), .A2(new_n733), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G27), .B2(new_n733), .ZN(new_n766));
  INV_X1    g341(.A(G2078), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n764), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n755), .B(new_n768), .C1(new_n767), .C2(new_n766), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n733), .A2(G35), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G162), .B2(new_n733), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT29), .B(G2090), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n753), .A2(new_n754), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT24), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n733), .B1(new_n775), .B2(G34), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n776), .A2(KEYINPUT90), .B1(new_n775), .B2(G34), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(KEYINPUT90), .B2(new_n776), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT91), .Z(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G29), .B2(G160), .ZN(new_n780));
  INV_X1    g355(.A(G2084), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n769), .A2(new_n773), .A3(new_n774), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G29), .A2(G32), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n481), .A2(G141), .A3(new_n473), .ZN(new_n785));
  NAND3_X1  g360(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT26), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n481), .A2(G129), .A3(G2105), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n466), .A2(G105), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n785), .A2(new_n788), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT92), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT93), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n793), .A2(KEYINPUT93), .A3(new_n794), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n784), .B1(new_n800), .B2(G29), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT27), .B(G1996), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n703), .A2(G19), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n548), .B2(new_n703), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(G1341), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n703), .A2(G4), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n612), .B2(new_n703), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(G1348), .ZN(new_n809));
  AOI211_X1 g384(.A(new_n806), .B(new_n809), .C1(new_n742), .C2(new_n740), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n703), .A2(G20), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT23), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n572), .B2(new_n703), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n808), .A2(G1348), .B1(new_n813), .B2(G1956), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n813), .A2(G1956), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G1341), .B2(new_n805), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n810), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  NOR4_X1   g392(.A1(new_n744), .A2(new_n783), .A3(new_n803), .A4(new_n817), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n730), .A2(new_n818), .ZN(G311));
  NAND2_X1  g394(.A1(new_n730), .A2(new_n818), .ZN(G150));
  OAI21_X1  g395(.A(G55), .B1(new_n536), .B2(new_n537), .ZN(new_n821));
  NAND2_X1  g396(.A1(G80), .A2(G543), .ZN(new_n822));
  INV_X1    g397(.A(G67), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n523), .B2(new_n823), .ZN(new_n824));
  AOI22_X1  g399(.A1(G651), .A2(new_n824), .B1(new_n530), .B2(G93), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G860), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT37), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n612), .A2(G559), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT38), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n542), .A2(new_n543), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n831), .A2(G651), .A3(new_n545), .ZN(new_n832));
  INV_X1    g407(.A(new_n539), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(G43), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n512), .B2(new_n514), .ZN(new_n836));
  INV_X1    g411(.A(G55), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n512), .B2(new_n514), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n824), .A2(G651), .ZN(new_n839));
  INV_X1    g414(.A(G93), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n840), .B2(new_n529), .ZN(new_n841));
  OAI22_X1  g416(.A1(new_n834), .A2(new_n836), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n538), .A2(new_n821), .A3(new_n546), .A4(new_n825), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n830), .B(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT39), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(KEYINPUT95), .ZN(new_n848));
  INV_X1    g423(.A(G860), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n848), .B(new_n849), .C1(new_n846), .C2(new_n845), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n847), .A2(KEYINPUT95), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n828), .B1(new_n850), .B2(new_n851), .ZN(G145));
  NOR2_X1   g427(.A1(new_n751), .A2(new_n795), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n799), .B2(new_n751), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n490), .A2(new_n493), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT97), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n490), .A2(new_n493), .A3(KEYINPUT97), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n489), .A2(new_n859), .A3(new_n762), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n762), .B1(new_n489), .B2(new_n859), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n631), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n698), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n465), .A2(G142), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n620), .A2(G130), .ZN(new_n867));
  OR2_X1    g442(.A1(G106), .A2(G2105), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n868), .B(G2104), .C1(G118), .C2(new_n473), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n695), .A2(new_n696), .A3(new_n697), .A4(KEYINPUT98), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n865), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n870), .B1(new_n865), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n489), .A2(new_n859), .ZN(new_n875));
  INV_X1    g450(.A(new_n762), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n631), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n877), .A2(new_n878), .A3(new_n860), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n863), .A2(new_n874), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n874), .B1(new_n863), .B2(new_n879), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n854), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NOR3_X1   g457(.A1(new_n861), .A2(new_n862), .A3(new_n631), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n878), .B1(new_n877), .B2(new_n860), .ZN(new_n884));
  OAI22_X1  g459(.A1(new_n883), .A2(new_n884), .B1(new_n873), .B2(new_n872), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n793), .A2(KEYINPUT93), .A3(new_n794), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT93), .B1(new_n793), .B2(new_n794), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n751), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n751), .A2(new_n795), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n863), .A2(new_n874), .A3(new_n879), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n885), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n882), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n467), .A2(new_n471), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(new_n485), .B2(new_n486), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n477), .A2(new_n484), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(KEYINPUT68), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n477), .A2(new_n478), .A3(new_n484), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(G160), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT96), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n895), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n900), .B1(new_n895), .B2(new_n899), .ZN(new_n903));
  NOR3_X1   g478(.A1(new_n902), .A2(new_n903), .A3(new_n627), .ZN(new_n904));
  INV_X1    g479(.A(new_n627), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n895), .A2(new_n899), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT96), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n905), .B1(new_n907), .B2(new_n901), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT99), .B1(new_n904), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n627), .B1(new_n902), .B2(new_n903), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n907), .A2(new_n905), .A3(new_n901), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT99), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n893), .A2(new_n909), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT100), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n893), .A2(new_n909), .A3(KEYINPUT100), .A4(new_n913), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n910), .A2(new_n911), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n919), .A2(new_n882), .A3(new_n892), .ZN(new_n920));
  INV_X1    g495(.A(G37), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n918), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT101), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT101), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n918), .A2(new_n926), .A3(new_n923), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g504(.A1(new_n826), .A2(G868), .ZN(new_n930));
  XNOR2_X1  g505(.A(G290), .B(G305), .ZN(new_n931));
  INV_X1    g506(.A(G288), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(G166), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n931), .B(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT42), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n556), .B(KEYINPUT9), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n563), .A2(new_n570), .A3(new_n567), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n604), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n595), .B(new_n603), .C1(new_n558), .C2(new_n571), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(new_n940), .A3(KEYINPUT41), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT103), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n939), .A2(new_n940), .A3(new_n943), .A4(KEYINPUT41), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n939), .A2(new_n940), .A3(KEYINPUT102), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT41), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT102), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n572), .A2(new_n948), .A3(new_n604), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n945), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n939), .A2(new_n940), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n844), .B(new_n615), .ZN(new_n953));
  MUX2_X1   g528(.A(new_n951), .B(new_n952), .S(new_n953), .Z(new_n954));
  OAI21_X1  g529(.A(KEYINPUT104), .B1(new_n936), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n936), .A2(new_n954), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n955), .B(new_n956), .Z(new_n957));
  AOI21_X1  g532(.A(new_n930), .B1(new_n957), .B2(G868), .ZN(G295));
  AOI21_X1  g533(.A(new_n930), .B1(new_n957), .B2(G868), .ZN(G331));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n842), .A2(new_n843), .A3(G301), .ZN(new_n961));
  AOI21_X1  g536(.A(G301), .B1(new_n842), .B2(new_n843), .ZN(new_n962));
  OAI21_X1  g537(.A(G286), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AND4_X1   g538(.A1(new_n538), .A2(new_n821), .A3(new_n546), .A4(new_n825), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n538), .A2(new_n546), .B1(new_n821), .B2(new_n825), .ZN(new_n965));
  OAI21_X1  g540(.A(G171), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n842), .A2(new_n843), .A3(G301), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(G168), .A3(new_n967), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n963), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n951), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT106), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n931), .B(new_n933), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT106), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n969), .A2(new_n951), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n963), .A2(new_n968), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n952), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n971), .A2(new_n972), .A3(new_n974), .A4(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n971), .A2(new_n974), .A3(new_n976), .ZN(new_n979));
  AOI21_X1  g554(.A(G37), .B1(new_n979), .B2(new_n935), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT107), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n974), .A2(new_n976), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n973), .B1(new_n969), .B2(new_n951), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n935), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n981), .B1(new_n986), .B2(new_n921), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n982), .A2(new_n983), .A3(new_n988), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n946), .A2(new_n949), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n975), .A2(new_n947), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n972), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n991), .A2(new_n952), .ZN(new_n993));
  AOI21_X1  g568(.A(G37), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n977), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT43), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n960), .B1(new_n989), .B2(new_n996), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n994), .A2(new_n977), .A3(new_n983), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n982), .A2(new_n988), .ZN(new_n999));
  INV_X1    g574(.A(new_n983), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n997), .B1(new_n960), .B2(new_n1001), .ZN(G397));
  AOI21_X1  g577(.A(G1384), .B1(new_n489), .B2(new_n859), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT45), .B1(new_n1004), .B2(KEYINPUT108), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(KEYINPUT108), .B2(new_n1004), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n467), .A2(G40), .A3(new_n471), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1007), .B(KEYINPUT109), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(G290), .A2(G1986), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1012), .A2(KEYINPUT48), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n762), .B(G2067), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n795), .B2(G1996), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(new_n799), .B2(G1996), .ZN(new_n1016));
  XOR2_X1   g591(.A(new_n698), .B(new_n700), .Z(new_n1017));
  OAI21_X1  g592(.A(new_n1010), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1019), .B1(KEYINPUT48), .B2(new_n1012), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n795), .A2(new_n1014), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT46), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1010), .A2(new_n1021), .B1(KEYINPUT126), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G1996), .ZN(new_n1024));
  AOI211_X1 g599(.A(KEYINPUT126), .B(new_n1022), .C1(new_n1010), .C2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1022), .A2(KEYINPUT126), .ZN(new_n1026));
  NOR4_X1   g601(.A1(new_n1006), .A2(G1996), .A3(new_n1009), .A4(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1023), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g603(.A(new_n1028), .B(KEYINPUT47), .Z(new_n1029));
  NAND4_X1  g604(.A1(new_n695), .A2(new_n696), .A3(new_n697), .A4(new_n700), .ZN(new_n1030));
  OAI22_X1  g605(.A1(new_n1016), .A2(new_n1030), .B1(G2067), .B2(new_n762), .ZN(new_n1031));
  AOI211_X1 g606(.A(new_n1020), .B(new_n1029), .C1(new_n1010), .C2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G8), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1033), .B1(new_n1008), .B2(new_n1003), .ZN(new_n1034));
  INV_X1    g609(.A(G1981), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n584), .A2(new_n1035), .ZN(new_n1036));
  XOR2_X1   g611(.A(KEYINPUT113), .B(G86), .Z(new_n1037));
  NOR2_X1   g612(.A1(new_n529), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(G1981), .B1(new_n582), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT49), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1036), .A2(KEYINPUT49), .A3(new_n1039), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1034), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n1044), .A2(KEYINPUT114), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(KEYINPUT114), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(G288), .A2(G1976), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1047), .A2(new_n1048), .B1(new_n1035), .B2(new_n584), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1034), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1008), .A2(new_n1003), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n932), .A2(G1976), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(G8), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT52), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  OR3_X1    g631(.A1(new_n932), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n1047), .ZN(new_n1061));
  NAND2_X1  g636(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n1063));
  NOR2_X1   g638(.A1(G166), .A2(new_n1033), .ZN(new_n1064));
  MUX2_X1   g639(.A(new_n1062), .B(new_n1063), .S(new_n1064), .Z(new_n1065));
  NAND2_X1  g640(.A1(new_n1003), .A2(KEYINPUT45), .ZN(new_n1066));
  INV_X1    g641(.A(G1384), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n494), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT45), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1008), .A2(new_n1066), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G1971), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT50), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1003), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1068), .A2(KEYINPUT50), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1008), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(G2090), .ZN(new_n1079));
  OAI211_X1 g654(.A(G8), .B(new_n1065), .C1(new_n1074), .C2(new_n1079), .ZN(new_n1080));
  OAI22_X1  g655(.A1(new_n1049), .A2(new_n1050), .B1(new_n1061), .B2(new_n1080), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1058), .A2(new_n1059), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1007), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT109), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n494), .A2(KEYINPUT45), .A3(new_n1067), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT109), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1007), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1003), .A2(KEYINPUT45), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n738), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1008), .A2(new_n1077), .A3(new_n781), .A4(new_n1076), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1033), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(G286), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1065), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1084), .B(new_n1087), .C1(new_n1068), .C2(KEYINPUT50), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1003), .A2(new_n1075), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G2090), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1100), .A2(new_n1073), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1095), .B1(new_n1101), .B2(new_n1033), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1082), .A2(new_n1094), .A3(new_n1102), .A4(new_n1080), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT63), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n1093), .A2(new_n1104), .A3(G286), .ZN(new_n1106));
  OAI21_X1  g681(.A(G8), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n1095), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1082), .A2(new_n1106), .A3(new_n1080), .A4(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1081), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(G168), .A2(new_n1033), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT123), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1114), .B(KEYINPUT51), .C1(new_n1092), .C2(new_n1112), .ZN(new_n1115));
  OR3_X1    g690(.A1(new_n1092), .A2(new_n1112), .A3(KEYINPUT51), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1117), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT62), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT124), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(new_n1124), .A3(new_n1118), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1060), .A2(new_n1047), .A3(new_n1080), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1102), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT125), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1082), .A2(new_n1102), .A3(new_n1130), .A4(new_n1080), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT117), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1078), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1078), .A2(new_n1132), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1133), .A2(new_n740), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT53), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1071), .B2(G2078), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n767), .A2(KEYINPUT53), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1135), .B(new_n1137), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1129), .A2(new_n1131), .A3(G171), .A4(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1110), .B1(new_n1126), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1123), .A2(new_n1118), .ZN(new_n1143));
  XNOR2_X1  g718(.A(G301), .B(KEYINPUT54), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1145));
  AOI211_X1 g720(.A(new_n1139), .B(new_n1083), .C1(KEYINPUT45), .C2(new_n1003), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1144), .B1(new_n1006), .B2(new_n1146), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1140), .A2(new_n1144), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1143), .A2(new_n1129), .A3(new_n1131), .A4(new_n1148), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n937), .A2(KEYINPUT115), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n571), .B1(KEYINPUT115), .B2(new_n937), .ZN(new_n1151));
  AOI21_X1  g726(.A(KEYINPUT57), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n1152), .A2(KEYINPUT116), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1152), .A2(KEYINPUT116), .B1(KEYINPUT57), .B2(new_n572), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(KEYINPUT56), .B(G2072), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1008), .A2(new_n1070), .A3(new_n1066), .A4(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1098), .B2(G1956), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(G1348), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1133), .A2(new_n1161), .A3(new_n1134), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n1051), .A2(G2067), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n604), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT118), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1167), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1160), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  XOR2_X1   g744(.A(KEYINPUT58), .B(G1341), .Z(new_n1170));
  NAND2_X1  g745(.A1(new_n1051), .A2(new_n1170), .ZN(new_n1171));
  XOR2_X1   g746(.A(KEYINPUT119), .B(G1996), .Z(new_n1172));
  NAND4_X1  g747(.A1(new_n1008), .A2(new_n1070), .A3(new_n1066), .A4(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n547), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT120), .ZN(new_n1175));
  OR2_X1    g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1176), .A2(KEYINPUT59), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT121), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT59), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1179), .B1(new_n1174), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1178), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1160), .A2(KEYINPUT61), .A3(new_n1167), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1167), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1184), .B1(new_n1185), .B2(new_n1159), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1176), .A2(new_n1179), .A3(KEYINPUT59), .A4(new_n1177), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1182), .A2(new_n1183), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1162), .A2(new_n612), .A3(new_n1163), .ZN(new_n1189));
  OR2_X1    g764(.A1(new_n1189), .A2(KEYINPUT60), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n612), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1189), .A2(KEYINPUT60), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1190), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1169), .B1(new_n1188), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1149), .B1(new_n1194), .B2(KEYINPUT122), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT122), .ZN(new_n1196));
  OAI211_X1 g771(.A(new_n1196), .B(new_n1169), .C1(new_n1188), .C2(new_n1193), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1142), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n684), .A2(new_n687), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1010), .B1(new_n1200), .B2(KEYINPUT110), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT110), .ZN(new_n1202));
  NOR3_X1   g777(.A1(new_n1199), .A2(new_n1202), .A3(new_n1011), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1018), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1032), .B1(new_n1198), .B2(new_n1204), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g780(.A1(new_n986), .A2(new_n981), .A3(new_n921), .ZN(new_n1207));
  NAND2_X1  g781(.A1(new_n1207), .A2(new_n977), .ZN(new_n1208));
  OAI21_X1  g782(.A(new_n1000), .B1(new_n1208), .B2(new_n987), .ZN(new_n1209));
  NAND3_X1  g783(.A1(new_n994), .A2(new_n977), .A3(new_n983), .ZN(new_n1210));
  NAND2_X1  g784(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g785(.A1(new_n664), .A2(G319), .ZN(new_n1212));
  NOR3_X1   g786(.A1(G229), .A2(new_n652), .A3(new_n1212), .ZN(new_n1213));
  AOI21_X1  g787(.A(new_n926), .B1(new_n918), .B2(new_n923), .ZN(new_n1214));
  AOI211_X1 g788(.A(KEYINPUT101), .B(new_n922), .C1(new_n916), .C2(new_n917), .ZN(new_n1215));
  OAI21_X1  g789(.A(new_n1213), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g790(.A(new_n1216), .ZN(new_n1217));
  AOI21_X1  g791(.A(KEYINPUT127), .B1(new_n1211), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g792(.A(KEYINPUT127), .ZN(new_n1219));
  AOI211_X1 g793(.A(new_n1219), .B(new_n1216), .C1(new_n1209), .C2(new_n1210), .ZN(new_n1220));
  NOR2_X1   g794(.A1(new_n1218), .A2(new_n1220), .ZN(G308));
  OAI21_X1  g795(.A(new_n1219), .B1(new_n1001), .B2(new_n1216), .ZN(new_n1222));
  NAND3_X1  g796(.A1(new_n1211), .A2(new_n1217), .A3(KEYINPUT127), .ZN(new_n1223));
  NAND2_X1  g797(.A1(new_n1222), .A2(new_n1223), .ZN(G225));
endmodule


