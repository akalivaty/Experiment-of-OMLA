//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n631, new_n634, new_n635, new_n637, new_n638, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND3_X1   g036(.A1(KEYINPUT68), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(KEYINPUT3), .B1(KEYINPUT68), .B2(G2104), .ZN(new_n463));
  OR2_X1    g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT69), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n462), .A2(new_n463), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(new_n471), .A3(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT67), .ZN(new_n477));
  OR2_X1    g052(.A1(new_n476), .A2(KEYINPUT67), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n475), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n465), .A2(G2104), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT70), .Z(new_n481));
  AOI22_X1  g056(.A1(G2105), .A2(new_n479), .B1(new_n481), .B2(G101), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n473), .A2(new_n482), .ZN(G160));
  NAND2_X1  g058(.A1(new_n470), .A2(G136), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n486));
  INV_X1    g061(.A(G124), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n464), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n484), .B(new_n486), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND3_X1  g065(.A1(new_n464), .A2(G126), .A3(G2105), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n465), .C1(new_n462), .C2(new_n463), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n498), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n474), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n495), .A2(KEYINPUT71), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n496), .A2(KEYINPUT4), .B1(new_n474), .B2(new_n499), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n494), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n502), .A2(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT72), .B1(new_n507), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT73), .B1(new_n510), .B2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(new_n507), .A3(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n512), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT74), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n512), .A2(new_n516), .A3(KEYINPUT74), .A4(new_n517), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G88), .ZN(new_n524));
  NAND2_X1  g099(.A1(G75), .A2(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n512), .A2(new_n516), .ZN(new_n526));
  INV_X1    g101(.A(G62), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n517), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n528), .A2(G651), .B1(G50), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n524), .A2(new_n531), .ZN(G303));
  INV_X1    g107(.A(G303), .ZN(G166));
  INV_X1    g108(.A(KEYINPUT75), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n512), .A2(new_n516), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n534), .B1(new_n512), .B2(new_n516), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n537), .A2(G63), .A3(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n520), .A2(G89), .A3(new_n521), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XOR2_X1   g115(.A(new_n540), .B(KEYINPUT7), .Z(new_n541));
  INV_X1    g116(.A(KEYINPUT76), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n529), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n517), .A2(KEYINPUT76), .A3(G543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n541), .B1(new_n545), .B2(G51), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n538), .A2(new_n539), .A3(new_n546), .ZN(G286));
  INV_X1    g122(.A(G286), .ZN(G168));
  INV_X1    g123(.A(G651), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n526), .A2(KEYINPUT75), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n512), .A2(new_n516), .A3(new_n534), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n550), .A2(G64), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(G77), .A2(G543), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n549), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g129(.A(KEYINPUT77), .B(G90), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n520), .A2(new_n521), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n545), .A2(G52), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n554), .A2(new_n558), .ZN(G171));
  NAND3_X1  g134(.A1(new_n520), .A2(G81), .A3(new_n521), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n545), .A2(G43), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(G68), .A2(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n550), .A2(new_n551), .ZN(new_n564));
  INV_X1    g139(.A(G56), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n562), .B1(G651), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  NAND2_X1  g147(.A1(KEYINPUT78), .A2(KEYINPUT9), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n530), .A2(G53), .A3(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  OAI211_X1 g150(.A(KEYINPUT78), .B(KEYINPUT9), .C1(new_n529), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(G91), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n522), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(G65), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n526), .A2(KEYINPUT79), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n512), .A2(new_n516), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n581), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(G78), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n580), .A2(new_n588), .ZN(G299));
  INV_X1    g164(.A(G171), .ZN(G301));
  NAND2_X1  g165(.A1(new_n523), .A2(G87), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n530), .A2(G49), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(G74), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n549), .B1(new_n564), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n593), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G288));
  NAND2_X1  g175(.A1(new_n523), .A2(G86), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n530), .A2(G48), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n512), .A2(new_n516), .A3(G61), .ZN(new_n603));
  NAND2_X1  g178(.A1(G73), .A2(G543), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n549), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n605), .A2(KEYINPUT81), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(KEYINPUT81), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n601), .A2(new_n602), .A3(new_n606), .A4(new_n607), .ZN(G305));
  NAND2_X1  g183(.A1(new_n537), .A2(G60), .ZN(new_n609));
  NAND2_X1  g184(.A1(G72), .A2(G543), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n549), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n545), .A2(G47), .ZN(new_n612));
  INV_X1    g187(.A(G85), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n522), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(G290));
  NAND2_X1  g191(.A1(G301), .A2(G868), .ZN(new_n617));
  AND3_X1   g192(.A1(new_n520), .A2(G92), .A3(new_n521), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT10), .ZN(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(new_n582), .B2(new_n584), .ZN(new_n621));
  AND2_X1   g196(.A1(G79), .A2(G543), .ZN(new_n622));
  OAI21_X1  g197(.A(G651), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n545), .A2(G54), .ZN(new_n624));
  AND2_X1   g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n619), .A2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n617), .B1(new_n627), .B2(G868), .ZN(G284));
  OAI21_X1  g203(.A(new_n617), .B1(new_n627), .B2(G868), .ZN(G321));
  NAND2_X1  g204(.A1(G286), .A2(G868), .ZN(new_n630));
  INV_X1    g205(.A(G299), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(G297));
  OAI21_X1  g207(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(G280));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n627), .B1(new_n634), .B2(G860), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT82), .ZN(G148));
  NAND2_X1  g211(.A1(new_n627), .A2(new_n634), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G868), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(G868), .B2(new_n567), .ZN(G323));
  XNOR2_X1  g214(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n640));
  XNOR2_X1  g215(.A(G323), .B(new_n640), .ZN(G282));
  NAND2_X1  g216(.A1(new_n481), .A2(new_n474), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT12), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT13), .Z(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(G2100), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(G2100), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n470), .A2(G135), .ZN(new_n647));
  INV_X1    g222(.A(G123), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n465), .A2(G111), .ZN(new_n649));
  OAI21_X1  g224(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n650));
  OAI221_X1 g225(.A(new_n647), .B1(new_n488), .B2(new_n648), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(G2096), .Z(new_n652));
  NAND3_X1  g227(.A1(new_n645), .A2(new_n646), .A3(new_n652), .ZN(G156));
  XNOR2_X1  g228(.A(G2427), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n658), .A3(KEYINPUT14), .ZN(new_n659));
  XOR2_X1   g234(.A(G1341), .B(G1348), .Z(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2443), .B(G2446), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT85), .ZN(new_n665));
  XOR2_X1   g240(.A(G2451), .B(G2454), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n663), .A2(new_n667), .ZN(new_n669));
  AND3_X1   g244(.A1(new_n668), .A2(G14), .A3(new_n669), .ZN(G401));
  INV_X1    g245(.A(KEYINPUT18), .ZN(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(KEYINPUT17), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n671), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2100), .ZN(new_n678));
  XOR2_X1   g253(.A(G2072), .B(G2078), .Z(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n674), .B2(KEYINPUT18), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G2096), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n678), .B(new_n681), .ZN(G227));
  XOR2_X1   g257(.A(G1971), .B(G1976), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1956), .B(G2474), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1961), .B(G1966), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n684), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n684), .A2(new_n687), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT20), .Z(new_n691));
  AOI211_X1 g266(.A(new_n689), .B(new_n691), .C1(new_n684), .C2(new_n688), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT86), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT87), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1981), .B(G1986), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(G229));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G20), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT23), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(new_n631), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1956), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT31), .B(G11), .Z(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT30), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(G28), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n709), .A2(KEYINPUT95), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n708), .B2(G28), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(KEYINPUT95), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n706), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT88), .B(G29), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n651), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n707), .A2(G33), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT25), .ZN(new_n718));
  AOI22_X1  g293(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n719), .A2(new_n465), .ZN(new_n720));
  AOI211_X1 g295(.A(new_n718), .B(new_n720), .C1(G139), .C2(new_n470), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n716), .B1(new_n721), .B2(new_n707), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n715), .B1(new_n722), .B2(G2072), .ZN(new_n723));
  INV_X1    g298(.A(new_n488), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G129), .ZN(new_n725));
  NAND3_X1  g300(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT26), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n481), .B2(G105), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n470), .A2(G141), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n725), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n731), .A2(new_n707), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n707), .B2(G32), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT27), .B(G1996), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  OAI221_X1 g311(.A(new_n723), .B1(G2072), .B2(new_n722), .C1(new_n734), .C2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n714), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(G35), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G162), .B2(new_n738), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT29), .B(G2090), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n714), .A2(G26), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT28), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n724), .A2(G128), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n470), .A2(G140), .ZN(new_n746));
  OR2_X1    g321(.A1(G104), .A2(G2105), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n747), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n744), .B1(new_n750), .B2(new_n707), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G2067), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n737), .A2(new_n742), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n701), .A2(G21), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G168), .B2(new_n701), .ZN(new_n755));
  INV_X1    g330(.A(G1966), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n738), .A2(G27), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G164), .B2(new_n738), .ZN(new_n759));
  INV_X1    g334(.A(G2078), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n753), .B(new_n757), .C1(KEYINPUT97), .C2(new_n761), .ZN(new_n762));
  AOI211_X1 g337(.A(new_n705), .B(new_n762), .C1(KEYINPUT97), .C2(new_n761), .ZN(new_n763));
  NOR2_X1   g338(.A1(G4), .A2(G16), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n627), .B2(G16), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT93), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT92), .B(G1348), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(G160), .A2(G29), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT24), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n770), .A2(G34), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(G34), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n714), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G2084), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n734), .A2(new_n736), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G171), .A2(new_n701), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G5), .B2(new_n701), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n776), .B1(new_n779), .B2(G1961), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n781), .A2(KEYINPUT96), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n781), .A2(KEYINPUT96), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n774), .A2(new_n775), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT94), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n701), .A2(G19), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n567), .B2(new_n701), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(G1341), .Z(new_n788));
  INV_X1    g363(.A(G1961), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n785), .B(new_n788), .C1(new_n789), .C2(new_n778), .ZN(new_n790));
  NOR3_X1   g365(.A1(new_n782), .A2(new_n783), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n763), .A2(new_n768), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n701), .A2(G23), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n599), .B2(new_n701), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT91), .Z(new_n795));
  XOR2_X1   g370(.A(KEYINPUT33), .B(G1976), .Z(new_n796));
  OR2_X1    g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n701), .A2(G22), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G166), .B2(new_n701), .ZN(new_n800));
  INV_X1    g375(.A(G1971), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT32), .B(G1981), .Z(new_n803));
  AND2_X1   g378(.A1(new_n701), .A2(G6), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G305), .B2(G16), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n802), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n803), .B2(new_n805), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n797), .A2(new_n798), .A3(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n738), .A2(G25), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n724), .A2(G119), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT89), .ZN(new_n813));
  OR2_X1    g388(.A1(G95), .A2(G2105), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n814), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT90), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G131), .B2(new_n470), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n811), .B1(new_n819), .B2(new_n738), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT35), .B(G1991), .Z(new_n821));
  XOR2_X1   g396(.A(new_n820), .B(new_n821), .Z(new_n822));
  NOR2_X1   g397(.A1(new_n615), .A2(new_n701), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n701), .B2(G24), .ZN(new_n824));
  INV_X1    g399(.A(G1986), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n822), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n809), .A2(new_n810), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(KEYINPUT36), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT36), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n809), .A2(new_n831), .A3(new_n810), .A4(new_n828), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n792), .B1(new_n830), .B2(new_n832), .ZN(G311));
  INV_X1    g408(.A(G311), .ZN(G150));
  NAND3_X1  g409(.A1(new_n520), .A2(G93), .A3(new_n521), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n545), .A2(G55), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(G67), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n535), .A2(new_n536), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(G80), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(new_n510), .ZN(new_n842));
  OAI21_X1  g417(.A(G651), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n838), .A2(new_n843), .A3(KEYINPUT98), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n550), .A2(G67), .A3(new_n551), .ZN(new_n846));
  INV_X1    g421(.A(new_n842), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n549), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n845), .B1(new_n848), .B2(new_n837), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n567), .B1(new_n844), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n566), .A2(G651), .ZN(new_n851));
  INV_X1    g426(.A(new_n562), .ZN(new_n852));
  AND4_X1   g427(.A1(new_n851), .A2(new_n852), .A3(new_n838), .A4(new_n843), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT38), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n626), .A2(new_n634), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT39), .ZN(new_n858));
  AOI21_X1  g433(.A(G860), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(new_n858), .B2(new_n857), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT99), .ZN(new_n861));
  AOI21_X1  g436(.A(KEYINPUT98), .B1(new_n838), .B2(new_n843), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n848), .A2(new_n837), .A3(new_n845), .ZN(new_n863));
  OAI21_X1  g438(.A(G860), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT37), .Z(new_n865));
  NAND2_X1  g440(.A1(new_n861), .A2(new_n865), .ZN(G145));
  XNOR2_X1  g441(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(G162), .B(new_n651), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(G160), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n501), .A2(KEYINPUT100), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n504), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n494), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n749), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n874), .A2(new_n749), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n730), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n877), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n879), .A2(new_n731), .A3(new_n875), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  OR3_X1    g456(.A1(new_n881), .A2(KEYINPUT102), .A3(new_n721), .ZN(new_n882));
  OAI21_X1  g457(.A(KEYINPUT102), .B1(new_n881), .B2(new_n721), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n721), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n881), .A2(KEYINPUT101), .A3(new_n721), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n818), .B(new_n643), .ZN(new_n891));
  OR2_X1    g466(.A1(G106), .A2(G2105), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n892), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n893));
  INV_X1    g468(.A(G130), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n893), .B1(new_n488), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n895), .B1(G142), .B2(new_n470), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n891), .B(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n890), .A2(new_n898), .ZN(new_n899));
  AOI22_X1  g474(.A1(new_n883), .A2(new_n882), .B1(new_n887), .B2(new_n888), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n900), .A2(new_n897), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n870), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(KEYINPUT103), .B1(new_n900), .B2(new_n897), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n870), .B1(new_n900), .B2(new_n897), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n890), .A2(new_n905), .A3(new_n898), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(G37), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n902), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n909), .A2(new_n910), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n868), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n909), .A2(new_n910), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(new_n911), .A3(new_n867), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(G395));
  NAND2_X1  g492(.A1(new_n851), .A2(new_n852), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(new_n862), .B2(new_n863), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n567), .A2(new_n843), .A3(new_n838), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n637), .B(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n626), .A2(KEYINPUT106), .A3(G299), .ZN(new_n923));
  INV_X1    g498(.A(new_n588), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT106), .B1(new_n924), .B2(new_n579), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n580), .A2(new_n926), .A3(new_n588), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n925), .A2(new_n927), .A3(new_n619), .A4(new_n625), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n923), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n922), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT41), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n923), .A2(new_n928), .A3(KEYINPUT41), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n930), .B1(new_n922), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT42), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n599), .B(G305), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n615), .B(G303), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n938), .B(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n941), .A2(KEYINPUT107), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT42), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n930), .B(new_n943), .C1(new_n922), .C2(new_n935), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n937), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n942), .B1(new_n937), .B2(new_n944), .ZN(new_n946));
  OAI21_X1  g521(.A(G868), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G868), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n862), .B2(new_n863), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(G295));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n947), .A2(new_n951), .A3(new_n949), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n951), .B1(new_n947), .B2(new_n949), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(G331));
  INV_X1    g529(.A(KEYINPUT110), .ZN(new_n955));
  OAI211_X1 g530(.A(G286), .B(new_n955), .C1(new_n554), .C2(new_n558), .ZN(new_n956));
  INV_X1    g531(.A(G64), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n535), .A2(new_n536), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n553), .ZN(new_n959));
  OAI21_X1  g534(.A(G651), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n960), .A2(KEYINPUT110), .A3(new_n557), .A4(new_n556), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n955), .B1(new_n554), .B2(new_n558), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(new_n962), .A3(G168), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n919), .A2(new_n920), .A3(new_n956), .A4(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n963), .A2(new_n956), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n967), .A2(new_n854), .A3(KEYINPUT112), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT111), .B1(new_n967), .B2(new_n854), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n963), .A2(new_n956), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n921), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n934), .B1(new_n969), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n967), .A2(new_n854), .ZN(new_n976));
  INV_X1    g551(.A(new_n964), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n976), .A2(new_n977), .A3(new_n929), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n941), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n921), .A2(new_n971), .A3(new_n972), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n971), .B1(new_n921), .B2(new_n972), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n966), .B(new_n968), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n935), .ZN(new_n983));
  INV_X1    g558(.A(new_n978), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(new_n940), .A3(new_n984), .ZN(new_n985));
  XOR2_X1   g560(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n986));
  AND4_X1   g561(.A1(new_n908), .A2(new_n979), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n978), .B1(new_n982), .B2(new_n935), .ZN(new_n989));
  AOI21_X1  g564(.A(G37), .B1(new_n989), .B2(new_n940), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n976), .A2(new_n977), .ZN(new_n991));
  OAI22_X1  g566(.A1(new_n982), .A2(new_n929), .B1(new_n934), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n941), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n988), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT44), .B1(new_n987), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n979), .A2(new_n985), .A3(new_n908), .ZN(new_n997));
  INV_X1    g572(.A(new_n986), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n990), .A2(new_n986), .A3(new_n993), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n995), .A2(new_n996), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n996), .B1(new_n995), .B2(new_n1002), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(G397));
  NAND2_X1  g580(.A1(new_n871), .A2(new_n873), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n495), .ZN(new_n1007));
  XOR2_X1   g582(.A(KEYINPUT114), .B(G1384), .Z(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n473), .A2(G40), .A3(new_n482), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1013), .A2(G1996), .A3(new_n730), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n1014), .A2(KEYINPUT115), .ZN(new_n1015));
  XOR2_X1   g590(.A(new_n749), .B(G2067), .Z(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(G1996), .B2(new_n730), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n1013), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1014), .A2(KEYINPUT115), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1015), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1013), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n615), .A2(new_n825), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G290), .A2(G1986), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n819), .A2(new_n821), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n819), .A2(new_n821), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1021), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1020), .A2(new_n1024), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n1029));
  INV_X1    g604(.A(G1384), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1007), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1012), .B1(new_n1031), .B2(new_n1010), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1010), .A2(G1384), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n502), .A2(new_n505), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT119), .ZN(new_n1035));
  OR2_X1    g610(.A1(new_n1034), .A2(KEYINPUT119), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1032), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n1038));
  OR3_X1    g613(.A1(new_n1037), .A2(new_n1038), .A3(G2078), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n874), .A2(G1384), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1012), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n502), .A2(new_n505), .A3(new_n1030), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT50), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n789), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1044), .A2(new_n1010), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1007), .A2(KEYINPUT45), .A3(new_n1008), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1048), .A2(new_n1049), .A3(new_n760), .A4(new_n1043), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1050), .A2(KEYINPUT124), .A3(new_n1038), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT124), .B1(new_n1050), .B2(new_n1038), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1039), .B(new_n1047), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1029), .B1(new_n1054), .B2(G301), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1012), .A2(new_n1038), .A3(G2078), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1011), .A2(new_n1049), .A3(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1047), .B(new_n1057), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1058), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT125), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1058), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1060), .B1(new_n1061), .B2(G301), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1055), .A2(new_n1059), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1053), .A2(G171), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1064), .B1(G171), .B2(new_n1058), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n1029), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1068));
  INV_X1    g643(.A(G1976), .ZN(new_n1069));
  OAI211_X1 g644(.A(G8), .B(new_n1068), .C1(G288), .C2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n599), .B2(G1976), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1067), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1072), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1068), .A2(G8), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(G1976), .B2(new_n599), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1074), .A2(new_n1076), .A3(KEYINPUT117), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(G303), .A2(G8), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n1079), .B(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1043), .B1(new_n1044), .B2(KEYINPUT50), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1082), .A2(new_n1083), .A3(G2090), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1048), .A2(new_n1049), .A3(new_n1043), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n801), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G8), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1081), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n601), .A2(new_n602), .ZN(new_n1089));
  OAI21_X1  g664(.A(G1981), .B1(new_n1089), .B2(new_n605), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(G305), .B2(G1981), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT49), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1075), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1093), .A2(new_n1094), .B1(new_n1070), .B2(KEYINPUT52), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1085), .A2(new_n801), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(G2090), .B2(new_n1046), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1081), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(new_n1098), .A3(G8), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1078), .A2(new_n1088), .A3(new_n1095), .A4(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1037), .A2(new_n756), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1042), .A2(new_n1045), .A3(new_n775), .A4(new_n1043), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1101), .A2(G168), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(G8), .ZN(new_n1104));
  AOI21_X1  g679(.A(G168), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT51), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT51), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(new_n1107), .A3(G8), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1100), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1063), .A2(new_n1066), .A3(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1012), .A2(G1996), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1048), .A2(new_n1049), .A3(new_n1111), .ZN(new_n1112));
  XOR2_X1   g687(.A(KEYINPUT58), .B(G1341), .Z(new_n1113));
  NAND2_X1  g688(.A1(new_n1068), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1112), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1115), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n567), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT59), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1068), .A2(G2067), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1120), .B1(new_n767), .B2(new_n1046), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1121), .A2(new_n626), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1121), .A2(new_n626), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT60), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(G299), .B(KEYINPUT57), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G1956), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT56), .B(G2072), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1048), .A2(new_n1049), .A3(new_n1043), .A4(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1126), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n1125), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT61), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n626), .A2(KEYINPUT60), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1134), .A2(new_n1135), .B1(new_n1121), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT121), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1132), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1128), .A2(KEYINPUT121), .A3(new_n1130), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1139), .A2(new_n1125), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1141), .A2(KEYINPUT61), .A3(new_n1131), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1119), .A2(new_n1124), .A3(new_n1137), .A4(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1141), .B1(new_n626), .B2(new_n1121), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n1131), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1143), .A2(KEYINPUT123), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT123), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1110), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1078), .A2(new_n1095), .ZN(new_n1149));
  NOR2_X1   g724(.A1(G305), .A2(G1981), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT118), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1152));
  NOR2_X1   g727(.A1(G288), .A2(G1976), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI22_X1  g729(.A1(new_n1149), .A2(new_n1099), .B1(new_n1154), .B2(new_n1075), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1097), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1081), .B1(new_n1156), .B2(new_n1087), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1078), .A2(new_n1157), .A3(new_n1095), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(KEYINPUT120), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT120), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1078), .A2(new_n1157), .A3(new_n1160), .A4(new_n1095), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1162));
  AND4_X1   g737(.A1(G8), .A2(new_n1099), .A3(G168), .A4(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1159), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1155), .B1(new_n1164), .B2(KEYINPUT63), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1162), .A2(G8), .A3(G168), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1166), .A2(KEYINPUT63), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1064), .B1(new_n1168), .B2(KEYINPUT62), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1106), .A2(new_n1170), .A3(new_n1108), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1167), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1165), .B1(new_n1172), .B2(new_n1100), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1028), .B1(new_n1148), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT46), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1175), .B1(new_n1021), .B2(G1996), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1016), .B(new_n731), .C1(new_n1175), .C2(G1996), .ZN(new_n1177));
  AOI22_X1  g752(.A1(new_n1176), .A2(KEYINPUT126), .B1(new_n1013), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1178), .B1(KEYINPUT126), .B2(new_n1176), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT47), .ZN(new_n1180));
  OAI22_X1  g755(.A1(new_n1020), .A2(new_n1026), .B1(G2067), .B2(new_n749), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n1013), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT48), .ZN(new_n1184));
  OR3_X1    g759(.A1(new_n1184), .A2(new_n1020), .A3(new_n1027), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1180), .A2(new_n1182), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1174), .A2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g763(.A1(new_n915), .A2(new_n911), .ZN(new_n1190));
  NAND2_X1  g764(.A1(new_n999), .A2(new_n1001), .ZN(new_n1191));
  NOR4_X1   g765(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1192));
  AND3_X1   g766(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(G308));
  NAND3_X1  g767(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(G225));
endmodule


