//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n615, new_n616,
    new_n619, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195, new_n1196,
    new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT67), .Z(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n463), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n468), .A2(G137), .A3(new_n463), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n471), .A2(new_n475), .ZN(G160));
  AOI21_X1  g051(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(G136), .B2(new_n482), .ZN(G162));
  AND2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  OAI211_X1 g060(.A(G138), .B(new_n463), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT4), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n468), .A2(new_n488), .A3(G138), .A4(new_n463), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n463), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT68), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n494), .A2(new_n496), .A3(new_n497), .A4(G2104), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n493), .A2(new_n498), .B1(new_n477), .B2(G126), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n490), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(G62), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(G75), .A2(G543), .ZN(new_n508));
  OAI21_X1  g083(.A(G651), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n511));
  OAI21_X1  g086(.A(G651), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT6), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n512), .A2(G50), .A3(G543), .A4(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT5), .B(G543), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n512), .A2(G88), .A3(new_n514), .A4(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n509), .A2(new_n515), .A3(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n522));
  AND2_X1   g097(.A1(G63), .A2(G651), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n521), .A2(new_n522), .B1(new_n516), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n512), .A2(G543), .A3(new_n514), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  INV_X1    g101(.A(G89), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n512), .A2(new_n514), .A3(new_n516), .ZN(new_n528));
  OAI221_X1 g103(.A(new_n524), .B1(new_n525), .B2(new_n526), .C1(new_n527), .C2(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  AND2_X1   g106(.A1(KEYINPUT5), .A2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(KEYINPUT5), .A2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n531), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G651), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n512), .A2(G52), .A3(G543), .A4(new_n514), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n512), .A2(G90), .A3(new_n514), .A4(new_n516), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(KEYINPUT70), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT70), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n537), .A2(new_n542), .A3(new_n538), .A4(new_n539), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n541), .A2(new_n543), .ZN(G171));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n534), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n513), .B1(new_n547), .B2(KEYINPUT71), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n548), .B1(KEYINPUT71), .B2(new_n547), .ZN(new_n549));
  INV_X1    g124(.A(new_n525), .ZN(new_n550));
  XNOR2_X1  g125(.A(KEYINPUT72), .B(G43), .ZN(new_n551));
  AND3_X1   g126(.A1(new_n512), .A2(new_n514), .A3(new_n516), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n550), .A2(new_n551), .B1(new_n552), .B2(G81), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(G860), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT73), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(new_n516), .A2(G65), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n513), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n512), .A2(G91), .A3(new_n514), .A4(new_n516), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(KEYINPUT74), .ZN(new_n566));
  INV_X1    g141(.A(new_n514), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n534), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n568), .A2(new_n569), .A3(G91), .A4(new_n512), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n564), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT9), .B1(new_n525), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g148(.A(KEYINPUT69), .B(KEYINPUT6), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n567), .B1(new_n574), .B2(G651), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n575), .A2(new_n576), .A3(G53), .A4(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n571), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  INV_X1    g155(.A(G74), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n513), .B1(new_n534), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(new_n552), .B2(G87), .ZN(new_n583));
  INV_X1    g158(.A(G49), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n525), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT75), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR3_X1   g162(.A1(new_n525), .A2(KEYINPUT75), .A3(new_n584), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n583), .B1(new_n587), .B2(new_n588), .ZN(G288));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(new_n505), .B2(new_n506), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n512), .A2(G86), .A3(new_n514), .A4(new_n516), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n512), .A2(G48), .A3(G543), .A4(new_n514), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(new_n550), .A2(G47), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n552), .A2(G85), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  OAI211_X1 g175(.A(new_n598), .B(new_n599), .C1(new_n513), .C2(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(new_n552), .A2(G92), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n534), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n550), .A2(G54), .B1(G651), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  MUX2_X1   g185(.A(G301), .B(new_n609), .S(new_n610), .Z(G321));
  XOR2_X1   g186(.A(G321), .B(KEYINPUT76), .Z(G284));
  AOI21_X1  g187(.A(G868), .B1(G299), .B2(KEYINPUT78), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(KEYINPUT78), .B2(G299), .ZN(new_n614));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT77), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n616), .ZN(G297));
  NAND2_X1  g192(.A1(new_n614), .A2(new_n616), .ZN(G280));
  INV_X1    g193(.A(new_n609), .ZN(new_n619));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n554), .A2(new_n610), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n609), .A2(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(new_n610), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n468), .A2(new_n473), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n629), .A2(G2100), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT79), .Z(new_n631));
  NAND2_X1  g206(.A1(new_n482), .A2(G135), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n477), .A2(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n463), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2096), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n629), .B2(G2100), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n631), .A2(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT83), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2427), .B(G2430), .Z(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT82), .B(KEYINPUT14), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n642), .A2(new_n643), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G1341), .B(G1348), .Z(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT81), .ZN(new_n653));
  XOR2_X1   g228(.A(G2451), .B(G2454), .Z(new_n654));
  XOR2_X1   g229(.A(new_n653), .B(new_n654), .Z(new_n655));
  OR2_X1    g230(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n651), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G401));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT17), .Z(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  INV_X1    g240(.A(new_n662), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(new_n660), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n664), .B(new_n665), .C1(new_n663), .C2(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n660), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT18), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2100), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT84), .B(G2096), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  XOR2_X1   g249(.A(G1971), .B(G1976), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT20), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n677), .A2(new_n678), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n676), .A2(new_n679), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(new_n676), .B2(new_n682), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT85), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT86), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n688), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G229));
  INV_X1    g268(.A(G29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G33), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT25), .Z(new_n697));
  NAND2_X1  g272(.A1(new_n482), .A2(G139), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n468), .A2(G127), .ZN(new_n700));
  NAND2_X1  g275(.A1(G115), .A2(G2104), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n463), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n695), .B1(new_n703), .B2(new_n694), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n704), .A2(G2072), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT93), .Z(new_n706));
  NOR2_X1   g281(.A1(G4), .A2(G16), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n619), .B2(G16), .ZN(new_n708));
  NOR2_X1   g283(.A1(G29), .A2(G35), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G162), .B2(G29), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  OAI221_X1 g287(.A(new_n706), .B1(G1348), .B2(new_n708), .C1(G2090), .C2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n694), .A2(G32), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n477), .A2(G129), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT94), .Z(new_n716));
  AND2_X1   g291(.A1(new_n473), .A2(G105), .ZN(new_n717));
  NAND3_X1  g292(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT26), .ZN(new_n719));
  AOI211_X1 g294(.A(new_n717), .B(new_n719), .C1(G141), .C2(new_n482), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n714), .B1(new_n722), .B2(new_n694), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT27), .B(G1996), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  MUX2_X1   g300(.A(G21), .B(G286), .S(G16), .Z(new_n726));
  XOR2_X1   g301(.A(KEYINPUT95), .B(G1966), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n704), .A2(G2072), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT24), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n694), .B1(new_n730), .B2(G34), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n730), .B2(G34), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G160), .B2(G29), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(G2084), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n733), .A2(G2084), .ZN(new_n735));
  NOR3_X1   g310(.A1(new_n729), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n708), .A2(G1348), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n725), .A2(new_n728), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT89), .B(G16), .Z(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(G19), .ZN(new_n741));
  INV_X1    g316(.A(new_n554), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(new_n740), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(G1341), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n694), .A2(G26), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT28), .Z(new_n746));
  NAND2_X1  g321(.A1(new_n482), .A2(G140), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n477), .A2(G128), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n463), .A2(G116), .ZN(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n747), .B(new_n748), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT92), .Z(new_n752));
  AOI21_X1  g327(.A(new_n746), .B1(new_n752), .B2(G29), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G2067), .ZN(new_n754));
  NOR2_X1   g329(.A1(G27), .A2(G29), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G164), .B2(G29), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n756), .A2(G2078), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(G2078), .ZN(new_n758));
  OR3_X1    g333(.A1(new_n636), .A2(KEYINPUT96), .A3(new_n694), .ZN(new_n759));
  OAI21_X1  g334(.A(KEYINPUT96), .B1(new_n636), .B2(new_n694), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT31), .B(G11), .Z(new_n761));
  INV_X1    g336(.A(G28), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(KEYINPUT30), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT97), .ZN(new_n764));
  AOI21_X1  g339(.A(G29), .B1(new_n762), .B2(KEYINPUT30), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n761), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n759), .A2(new_n760), .A3(new_n766), .ZN(new_n767));
  NOR3_X1   g342(.A1(new_n757), .A2(new_n758), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n744), .A2(new_n754), .A3(new_n768), .ZN(new_n769));
  NOR3_X1   g344(.A1(new_n713), .A2(new_n738), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n712), .A2(G2090), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT99), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n739), .A2(G20), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT23), .Z(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G299), .B2(G16), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1956), .ZN(new_n776));
  NOR2_X1   g351(.A1(G5), .A2(G16), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G171), .B2(G16), .ZN(new_n778));
  INV_X1    g353(.A(G1961), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n770), .A2(new_n772), .A3(new_n776), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n482), .A2(G131), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n477), .A2(G119), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n463), .A2(G107), .ZN(new_n784));
  OAI21_X1  g359(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n782), .B(new_n783), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT87), .Z(new_n787));
  MUX2_X1   g362(.A(G25), .B(new_n787), .S(G29), .Z(new_n788));
  XOR2_X1   g363(.A(KEYINPUT35), .B(G1991), .Z(new_n789));
  OR2_X1    g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  AND3_X1   g366(.A1(new_n790), .A2(KEYINPUT88), .A3(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n740), .A2(G24), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G290), .B2(new_n739), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT90), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G1986), .Z(new_n796));
  AOI21_X1  g371(.A(KEYINPUT88), .B1(new_n790), .B2(new_n791), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n792), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  MUX2_X1   g373(.A(G6), .B(G305), .S(G16), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT91), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT32), .B(G1981), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(G23), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n803), .A2(G16), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G288), .B2(G16), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT33), .B(G1976), .Z(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n805), .A2(new_n807), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n740), .A2(G22), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G166), .B2(new_n740), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G1971), .Z(new_n812));
  NAND4_X1  g387(.A1(new_n802), .A2(new_n808), .A3(new_n809), .A4(new_n812), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(KEYINPUT34), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(KEYINPUT34), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n798), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(KEYINPUT36), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT36), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n798), .A2(new_n814), .A3(new_n818), .A4(new_n815), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n781), .B1(new_n817), .B2(new_n819), .ZN(G311));
  XNOR2_X1  g395(.A(G311), .B(KEYINPUT100), .ZN(G150));
  AOI22_X1  g396(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n822), .A2(new_n513), .ZN(new_n823));
  INV_X1    g398(.A(G55), .ZN(new_n824));
  INV_X1    g399(.A(G93), .ZN(new_n825));
  OAI22_X1  g400(.A1(new_n824), .A2(new_n525), .B1(new_n528), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT101), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n575), .A2(G55), .A3(G543), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n568), .A2(G93), .A3(new_n512), .ZN(new_n830));
  AOI21_X1  g405(.A(KEYINPUT101), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n823), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G860), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT37), .Z(new_n834));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n832), .A2(KEYINPUT102), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT102), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n837), .B(new_n823), .C1(new_n828), .C2(new_n831), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n836), .A2(new_n742), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n742), .B1(new_n836), .B2(new_n838), .ZN(new_n840));
  OR3_X1    g415(.A1(new_n839), .A2(new_n840), .A3(KEYINPUT38), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n609), .A2(new_n620), .ZN(new_n842));
  OAI21_X1  g417(.A(KEYINPUT38), .B1(new_n839), .B2(new_n840), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n842), .B1(new_n841), .B2(new_n843), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n835), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(new_n555), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n844), .A2(new_n845), .A3(new_n835), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n834), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT103), .ZN(G145));
  INV_X1    g425(.A(G37), .ZN(new_n851));
  XOR2_X1   g426(.A(G160), .B(new_n636), .Z(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(G162), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n752), .B(new_n721), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n854), .A2(G164), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(G164), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR3_X1   g432(.A1(new_n699), .A2(KEYINPUT104), .A3(new_n702), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n627), .B(new_n786), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n482), .A2(G142), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT105), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n477), .A2(G130), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n463), .A2(G118), .ZN(new_n864));
  OAI21_X1  g439(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n862), .B(new_n863), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n860), .B(new_n866), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n703), .B(KEYINPUT104), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(new_n855), .B2(new_n856), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n859), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n867), .B1(new_n859), .B2(new_n869), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n853), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n853), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT106), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n870), .A2(new_n875), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n851), .B(new_n873), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g455(.A(new_n623), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(new_n839), .B2(new_n840), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT41), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n609), .A2(G299), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n571), .A2(new_n578), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(new_n604), .B2(new_n608), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n883), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n609), .A2(G299), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(new_n604), .A3(new_n608), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(KEYINPUT41), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n826), .B(new_n827), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n837), .B1(new_n892), .B2(new_n823), .ZN(new_n893));
  INV_X1    g468(.A(new_n838), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n554), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n836), .A2(new_n742), .A3(new_n838), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(new_n623), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n882), .A2(new_n891), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n884), .A2(new_n886), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n900), .B1(new_n882), .B2(new_n897), .ZN(new_n901));
  OAI21_X1  g476(.A(KEYINPUT42), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n901), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n904), .A3(new_n898), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  XOR2_X1   g481(.A(G288), .B(G305), .Z(new_n907));
  XNOR2_X1  g482(.A(G290), .B(G166), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n907), .B(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n909), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n902), .A2(new_n905), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n610), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(G868), .B1(new_n892), .B2(new_n823), .ZN(new_n914));
  OR3_X1    g489(.A1(new_n913), .A2(KEYINPUT107), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT107), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(G295));
  OR2_X1    g492(.A1(new_n913), .A2(new_n914), .ZN(G331));
  AND2_X1   g493(.A1(new_n887), .A2(new_n890), .ZN(new_n919));
  XNOR2_X1  g494(.A(G171), .B(G168), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n839), .A2(new_n840), .A3(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(G171), .B(G286), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n922), .B1(new_n895), .B2(new_n896), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n919), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n920), .B1(new_n839), .B2(new_n840), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n895), .A2(new_n896), .A3(new_n922), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(new_n926), .A3(new_n900), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(new_n909), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n851), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n909), .B1(new_n924), .B2(new_n927), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT43), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n928), .A2(new_n851), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n924), .A2(new_n927), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT108), .B1(new_n933), .B2(new_n911), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n935));
  AOI211_X1 g510(.A(new_n935), .B(new_n909), .C1(new_n924), .C2(new_n927), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n932), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n931), .B1(new_n937), .B2(KEYINPUT43), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n929), .A2(new_n930), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n939), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n941), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n942), .B1(new_n941), .B2(new_n945), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n940), .B1(new_n946), .B2(new_n947), .ZN(G397));
  INV_X1    g523(.A(KEYINPUT57), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n571), .A2(new_n949), .A3(new_n578), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n949), .B1(new_n571), .B2(new_n578), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G1956), .ZN(new_n953));
  XNOR2_X1  g528(.A(KEYINPUT110), .B(G40), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n471), .A2(new_n475), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(G1384), .B1(new_n490), .B2(new_n499), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT50), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI211_X1 g533(.A(KEYINPUT50), .B(G1384), .C1(new_n490), .C2(new_n499), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n953), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G1384), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n487), .A2(new_n489), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n493), .A2(new_n498), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n477), .A2(G126), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n961), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n956), .A2(KEYINPUT45), .ZN(new_n969));
  XNOR2_X1  g544(.A(KEYINPUT56), .B(G2072), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n968), .A2(new_n955), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n952), .B1(new_n960), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n952), .A2(new_n960), .A3(new_n971), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n973), .A2(new_n619), .ZN(new_n974));
  INV_X1    g549(.A(G1348), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n975), .B1(new_n958), .B2(new_n959), .ZN(new_n976));
  INV_X1    g551(.A(G2067), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n955), .A2(new_n956), .A3(new_n977), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n976), .A2(new_n978), .A3(KEYINPUT121), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT121), .B1(new_n976), .B2(new_n978), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n972), .B1(new_n974), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT122), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n973), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(new_n972), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n960), .A2(new_n971), .ZN(new_n987));
  INV_X1    g562(.A(new_n952), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(new_n988), .A3(KEYINPUT122), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT61), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n986), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n987), .A2(new_n988), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n993), .A2(KEYINPUT61), .A3(new_n973), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT59), .ZN(new_n995));
  INV_X1    g570(.A(G1996), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n968), .A2(new_n996), .A3(new_n955), .A4(new_n969), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n955), .A2(new_n956), .ZN(new_n998));
  XOR2_X1   g573(.A(KEYINPUT58), .B(G1341), .Z(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n995), .B1(new_n1001), .B2(new_n742), .ZN(new_n1002));
  AOI211_X1 g577(.A(KEYINPUT59), .B(new_n554), .C1(new_n997), .C2(new_n1000), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n994), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n992), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT60), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n981), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT121), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n469), .A2(new_n470), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(G2105), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n472), .A2(new_n474), .ZN(new_n1011));
  INV_X1    g586(.A(new_n954), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1013), .B1(new_n966), .B2(KEYINPUT50), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n956), .A2(new_n957), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1348), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n978), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1008), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n976), .A2(KEYINPUT121), .A3(new_n978), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n609), .B1(new_n1020), .B2(KEYINPUT60), .ZN(new_n1021));
  AOI211_X1 g596(.A(new_n1006), .B(new_n619), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1007), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n983), .B1(new_n1005), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1976), .ZN(new_n1025));
  OAI211_X1 g600(.A(G8), .B(new_n998), .C1(G288), .C2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT52), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n1028));
  INV_X1    g603(.A(G288), .ZN(new_n1029));
  XNOR2_X1  g604(.A(KEYINPUT115), .B(G1976), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1028), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1027), .B1(new_n1031), .B2(new_n1026), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT49), .ZN(new_n1034));
  XNOR2_X1  g609(.A(KEYINPUT116), .B(G1981), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n594), .A2(new_n595), .A3(new_n596), .A4(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT117), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n592), .B1(new_n534), .B2(new_n590), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1035), .B1(new_n1039), .B2(G651), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1040), .A2(new_n1041), .A3(new_n595), .A4(new_n596), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n1038), .A2(new_n1042), .B1(G1981), .B2(G305), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1034), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI221_X4 g620(.A(KEYINPUT118), .B1(G305), .B2(G1981), .C1(new_n1038), .C2(new_n1042), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1033), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G305), .A2(G1981), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1037), .A2(KEYINPUT117), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1037), .A2(KEYINPUT117), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT118), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1052), .A2(new_n1053), .A3(KEYINPUT119), .A4(new_n1034), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1047), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n998), .A2(G8), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1056), .B1(KEYINPUT49), .B2(new_n1043), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1032), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n966), .A2(KEYINPUT50), .ZN(new_n1059));
  INV_X1    g634(.A(G2090), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n955), .A4(new_n1015), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT45), .B1(new_n500), .B2(new_n961), .ZN(new_n1062));
  AOI211_X1 g637(.A(new_n967), .B(G1384), .C1(new_n490), .C2(new_n499), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1062), .A2(new_n1063), .A3(new_n1013), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT112), .B(G1971), .Z(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1061), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n1068));
  AND3_X1   g643(.A1(G303), .A2(G8), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1068), .B1(G303), .B2(G8), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT114), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(G303), .A2(G8), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1068), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n1075));
  NAND3_X1  g650(.A1(G303), .A2(G8), .A3(new_n1068), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1071), .A2(new_n1077), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1067), .A2(G8), .A3(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1080), .B1(new_n1067), .B2(G8), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(G2078), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1064), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G2078), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n968), .A2(new_n1086), .A3(new_n955), .A4(new_n969), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n1083), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n958), .A2(new_n959), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1085), .B(new_n1088), .C1(G1961), .C2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n1091));
  XNOR2_X1  g666(.A(G171), .B(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(G160), .A2(G40), .A3(new_n1084), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1062), .A2(new_n1063), .A3(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1089), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1096), .A2(new_n779), .B1(new_n1087), .B2(new_n1083), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1090), .A2(new_n1092), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1058), .A2(new_n1082), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G2084), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1059), .A2(new_n1100), .A3(new_n955), .A4(new_n1015), .ZN(new_n1101));
  INV_X1    g676(.A(new_n727), .ZN(new_n1102));
  OAI211_X1 g677(.A(G168), .B(new_n1101), .C1(new_n1064), .C2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1103), .A2(new_n1104), .A3(G8), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n1106), .A3(KEYINPUT51), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n968), .A2(new_n955), .A3(new_n969), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1100), .A2(new_n1089), .B1(new_n1108), .B2(new_n727), .ZN(new_n1109));
  INV_X1    g684(.A(G8), .ZN(new_n1110));
  OR3_X1    g685(.A1(new_n1109), .A2(new_n1110), .A3(G168), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1103), .A2(KEYINPUT124), .A3(G8), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1107), .B(new_n1111), .C1(new_n1112), .C2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1099), .A2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1024), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1057), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n1047), .B2(new_n1054), .ZN(new_n1120));
  NOR2_X1   g695(.A1(G288), .A2(G1976), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  OAI22_X1  g697(.A1(new_n1120), .A2(new_n1122), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1123));
  XOR2_X1   g698(.A(new_n1056), .B(KEYINPUT120), .Z(new_n1124));
  AOI22_X1  g699(.A1(new_n1123), .A2(new_n1124), .B1(new_n1058), .B2(new_n1079), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1066), .B1(new_n1126), .B2(new_n955), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n958), .A2(new_n959), .A3(G2090), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1078), .B(G8), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1108), .A2(new_n1065), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1110), .B1(new_n1130), .B2(new_n1061), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1129), .B1(new_n1131), .B2(new_n1080), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1132), .A2(new_n1120), .A3(new_n1032), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1109), .A2(new_n1110), .A3(G286), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT63), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  AND4_X1   g710(.A1(KEYINPUT63), .A2(new_n1058), .A3(new_n1082), .A4(new_n1134), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1125), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT125), .B1(new_n1118), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1058), .A2(new_n1079), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1058), .A2(new_n1082), .A3(new_n1134), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT63), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1133), .A2(KEYINPUT63), .A3(new_n1134), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1141), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1058), .A2(new_n1082), .A3(new_n1098), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n619), .B1(new_n981), .B2(new_n1006), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1020), .A2(KEYINPUT60), .A3(new_n609), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n1151), .A2(new_n1152), .B1(new_n981), .B2(new_n1006), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1154), .B(new_n994), .C1(new_n986), .C2(new_n991), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n982), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1150), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1146), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n1116), .A2(KEYINPUT62), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1116), .A2(KEYINPUT62), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1133), .A2(G171), .A3(new_n1090), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1138), .A2(new_n1159), .A3(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n752), .B(new_n977), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(new_n996), .B2(new_n722), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1062), .A2(new_n955), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT111), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1167), .A2(G1996), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1166), .A2(new_n1168), .B1(new_n722), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1168), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n786), .B(new_n789), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1167), .ZN(new_n1174));
  XNOR2_X1  g749(.A(G290), .B(G1986), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1173), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1164), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1171), .B1(new_n1165), .B2(new_n722), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1178), .B(new_n1179), .ZN(new_n1180));
  XOR2_X1   g755(.A(new_n1169), .B(KEYINPUT46), .Z(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT47), .Z(new_n1183));
  NOR2_X1   g758(.A1(new_n752), .A2(G2067), .ZN(new_n1184));
  INV_X1    g759(.A(new_n789), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n787), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1184), .B1(new_n1170), .B2(new_n1186), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1167), .A2(G1986), .A3(G290), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n1188), .B(KEYINPUT48), .ZN(new_n1189));
  OAI22_X1  g764(.A1(new_n1187), .A2(new_n1171), .B1(new_n1173), .B2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1183), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1177), .A2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g767(.A1(G227), .A2(new_n461), .A3(G401), .ZN(new_n1194));
  AND2_X1   g768(.A1(new_n1194), .A2(KEYINPUT127), .ZN(new_n1195));
  NOR2_X1   g769(.A1(new_n1194), .A2(KEYINPUT127), .ZN(new_n1196));
  NOR3_X1   g770(.A1(new_n1195), .A2(new_n1196), .A3(G229), .ZN(new_n1197));
  NAND3_X1  g771(.A1(new_n1197), .A2(new_n879), .A3(new_n938), .ZN(G225));
  INV_X1    g772(.A(G225), .ZN(G308));
endmodule


