//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1270, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  XOR2_X1   g0007(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT65), .ZN(new_n209));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n209), .B(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n211), .ZN(new_n218));
  INV_X1    g0018(.A(new_n201), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT66), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n216), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT67), .B(G68), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G58), .A2(G232), .ZN(new_n230));
  NAND4_X1  g0030(.A1(new_n227), .A2(new_n228), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n213), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n222), .B1(KEYINPUT1), .B2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G68), .Z(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G41), .ZN(new_n251));
  OAI211_X1 g0051(.A(G1), .B(G13), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n253));
  AND2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G226), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n256));
  INV_X1    g0056(.A(G274), .ZN(new_n257));
  NOR3_X1   g0057(.A1(new_n256), .A2(new_n257), .A3(new_n253), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(G222), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G77), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(G1698), .ZN(new_n265));
  INV_X1    g0065(.A(G223), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n263), .B1(new_n264), .B2(new_n261), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n260), .B1(new_n256), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G190), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n267), .A2(new_n256), .ZN(new_n270));
  OAI21_X1  g0070(.A(G200), .B1(new_n270), .B2(new_n260), .ZN(new_n271));
  NAND3_X1  g0071(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n217), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n211), .A2(G33), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n274), .B(KEYINPUT70), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT69), .ZN(new_n276));
  INV_X1    g0076(.A(G58), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT8), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT8), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G58), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT68), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n279), .A2(KEYINPUT68), .A3(G58), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n276), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n282), .A2(new_n276), .A3(new_n283), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n275), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n273), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT9), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n202), .ZN(new_n295));
  INV_X1    g0095(.A(new_n273), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n210), .A2(G20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n295), .B1(new_n298), .B2(new_n202), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  AND3_X1   g0100(.A1(new_n291), .A2(new_n292), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n292), .B1(new_n291), .B2(new_n300), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n269), .B(new_n271), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(KEYINPUT73), .A2(KEYINPUT10), .ZN(new_n304));
  OR2_X1    g0104(.A1(KEYINPUT73), .A2(KEYINPUT10), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n302), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n291), .A2(new_n292), .A3(new_n300), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n271), .A2(new_n269), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n309), .A2(KEYINPUT73), .A3(new_n310), .A4(KEYINPUT10), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n291), .A2(new_n300), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT71), .B(G179), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n268), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n312), .B(new_n314), .C1(G169), .C2(new_n268), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n306), .A2(new_n311), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT72), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n293), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n293), .A2(new_n317), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(new_n273), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(G68), .A3(new_n297), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(KEYINPUT12), .A3(new_n224), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n293), .A2(G68), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n323), .B(new_n324), .C1(KEYINPUT12), .C2(new_n325), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n224), .A2(G20), .B1(G50), .B2(new_n288), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n275), .B2(new_n264), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n328), .A2(KEYINPUT11), .A3(new_n273), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT11), .B1(new_n328), .B2(new_n273), .ZN(new_n330));
  NOR3_X1   g0130(.A1(new_n326), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT14), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n261), .A2(G232), .A3(G1698), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n261), .A2(G226), .A3(new_n262), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G33), .A2(G97), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n256), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n258), .B1(G238), .B2(new_n254), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT13), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n340), .B1(new_n338), .B2(new_n339), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n333), .B(G169), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n343), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n345), .A2(G179), .A3(new_n341), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n341), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n333), .B1(new_n348), .B2(G169), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n332), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(G200), .ZN(new_n351));
  INV_X1    g0151(.A(G190), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n331), .B(new_n351), .C1(new_n352), .C2(new_n348), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n322), .A2(G77), .A3(new_n297), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n278), .A2(new_n280), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n356), .A2(new_n288), .B1(G20), .B2(G77), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT15), .B(G87), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n357), .B1(new_n274), .B2(new_n358), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n359), .A2(new_n273), .B1(new_n264), .B2(new_n321), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n261), .A2(G232), .A3(new_n262), .ZN(new_n362));
  INV_X1    g0162(.A(G107), .ZN(new_n363));
  OAI221_X1 g0163(.A(new_n362), .B1(new_n363), .B2(new_n261), .C1(new_n265), .C2(new_n225), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n256), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n258), .B1(G244), .B2(new_n254), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n361), .B1(new_n368), .B2(G190), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(G200), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n313), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G169), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n367), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n361), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n371), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  OR3_X1    g0177(.A1(new_n316), .A2(new_n354), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT75), .ZN(new_n379));
  AND2_X1   g0179(.A1(KEYINPUT67), .A2(G68), .ZN(new_n380));
  NOR2_X1   g0180(.A1(KEYINPUT67), .A2(G68), .ZN(new_n381));
  OAI21_X1  g0181(.A(G58), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n211), .B1(new_n382), .B2(new_n219), .ZN(new_n383));
  INV_X1    g0183(.A(new_n288), .ZN(new_n384));
  INV_X1    g0184(.A(G159), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n379), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n386), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n201), .B1(new_n223), .B2(G58), .ZN(new_n389));
  OAI211_X1 g0189(.A(KEYINPUT75), .B(new_n388), .C1(new_n389), .C2(new_n211), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G68), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT3), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G33), .ZN(new_n396));
  AOI211_X1 g0196(.A(new_n393), .B(G20), .C1(new_n394), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n394), .A2(new_n396), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT74), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT74), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n261), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n401), .A3(new_n211), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n397), .B1(new_n402), .B2(new_n393), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n391), .B(KEYINPUT16), .C1(new_n392), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT76), .ZN(new_n405));
  INV_X1    g0205(.A(new_n397), .ZN(new_n406));
  AND3_X1   g0206(.A1(new_n394), .A2(new_n396), .A3(new_n400), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n400), .B1(new_n394), .B2(new_n396), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n407), .A2(new_n408), .A3(G20), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n406), .B1(new_n409), .B2(KEYINPUT7), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G68), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT76), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n411), .A2(new_n412), .A3(KEYINPUT16), .A4(new_n391), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n405), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT16), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT7), .B1(new_n398), .B2(new_n211), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n224), .B1(new_n417), .B2(new_n406), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n388), .B1(new_n389), .B2(new_n211), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n415), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n273), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n414), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n285), .A2(new_n286), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(new_n294), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n424), .B2(new_n298), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n261), .A2(G226), .A3(G1698), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n261), .A2(G223), .A3(new_n262), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G87), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n256), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n258), .B1(G232), .B2(new_n254), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n352), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(G200), .B2(new_n434), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n423), .A2(new_n427), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT17), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT77), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n432), .A2(new_n433), .A3(new_n372), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n440), .B(new_n441), .C1(new_n434), .C2(new_n374), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n432), .A2(new_n433), .A3(new_n372), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n374), .B1(new_n432), .B2(new_n433), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT77), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n421), .B1(new_n405), .B2(new_n413), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n446), .B1(new_n447), .B2(new_n426), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT18), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT18), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n446), .B(new_n450), .C1(new_n447), .C2(new_n426), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n423), .A2(KEYINPUT17), .A3(new_n427), .A4(new_n436), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n439), .A2(new_n449), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n378), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G45), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n455), .A2(G1), .ZN(new_n456));
  XNOR2_X1  g0256(.A(KEYINPUT5), .B(G41), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n256), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT84), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(new_n459), .A3(G264), .ZN(new_n460));
  AND2_X1   g0260(.A1(KEYINPUT5), .A2(G41), .ZN(new_n461));
  NOR2_X1   g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n456), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(G264), .A3(new_n252), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT84), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n463), .A2(new_n256), .A3(new_n257), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n261), .A2(G257), .A3(G1698), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G294), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n394), .A2(new_n396), .A3(G250), .A4(new_n262), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n467), .B1(new_n471), .B2(new_n256), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n464), .ZN(new_n474));
  OAI22_X1  g0274(.A1(new_n473), .A2(G200), .B1(G190), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n294), .A2(KEYINPUT25), .A3(new_n363), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT83), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT25), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(new_n293), .B2(G107), .ZN(new_n479));
  OR2_X1    g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n477), .A2(new_n479), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n210), .A2(G33), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n296), .A2(new_n482), .A3(new_n293), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n480), .A2(new_n481), .B1(G107), .B2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n394), .A2(new_n396), .A3(new_n211), .A4(G87), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT22), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT22), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n261), .A2(new_n488), .A3(new_n211), .A4(G87), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n363), .A2(KEYINPUT23), .A3(G20), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT23), .B1(new_n363), .B2(G20), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G116), .ZN(new_n493));
  OAI22_X1  g0293(.A1(new_n491), .A2(new_n492), .B1(G20), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT24), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT24), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n490), .A2(new_n498), .A3(new_n495), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT82), .B1(new_n500), .B2(new_n273), .ZN(new_n501));
  AOI211_X1 g0301(.A(KEYINPUT24), .B(new_n494), .C1(new_n487), .C2(new_n489), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n498), .B1(new_n490), .B2(new_n495), .ZN(new_n503));
  OAI211_X1 g0303(.A(KEYINPUT82), .B(new_n273), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n475), .B(new_n485), .C1(new_n501), .C2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT85), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n473), .A2(G179), .B1(G169), .B2(new_n474), .ZN(new_n508));
  INV_X1    g0308(.A(new_n485), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n273), .B1(new_n502), .B2(new_n503), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT82), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n509), .B1(new_n512), .B2(new_n504), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n506), .B(new_n507), .C1(new_n508), .C2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n485), .B1(new_n501), .B2(new_n505), .ZN(new_n516));
  INV_X1    g0316(.A(new_n508), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n507), .B1(new_n518), .B2(new_n506), .ZN(new_n519));
  OR2_X1    g0319(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT6), .ZN(new_n521));
  AND2_X1   g0321(.A1(G97), .A2(G107), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n521), .B1(new_n522), .B2(new_n205), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n363), .A2(KEYINPUT6), .A3(G97), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n211), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n384), .A2(new_n264), .ZN(new_n526));
  OAI21_X1  g0326(.A(KEYINPUT78), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(G107), .B1(new_n416), .B2(new_n397), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT78), .ZN(new_n529));
  INV_X1    g0329(.A(new_n526), .ZN(new_n530));
  NAND2_X1  g0330(.A1(KEYINPUT6), .A2(G97), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(G107), .ZN(new_n532));
  XNOR2_X1  g0332(.A(G97), .B(G107), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n532), .B1(new_n533), .B2(new_n521), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n529), .B(new_n530), .C1(new_n534), .C2(new_n211), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n527), .A2(new_n528), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n273), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n293), .A2(G97), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n484), .B2(G97), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n394), .A2(new_n396), .A3(G244), .A4(new_n262), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT4), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n261), .A2(KEYINPUT4), .A3(G244), .A4(new_n262), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G283), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n261), .A2(G250), .A3(G1698), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n543), .A2(new_n544), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n256), .ZN(new_n548));
  INV_X1    g0348(.A(new_n467), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n463), .A2(G257), .A3(new_n252), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n374), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n550), .B1(new_n547), .B2(new_n256), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n554), .A2(new_n549), .A3(new_n313), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n540), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT79), .ZN(new_n557));
  AOI211_X1 g0357(.A(new_n467), .B(new_n550), .C1(new_n547), .C2(new_n256), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n537), .A2(new_n539), .B1(new_n558), .B2(new_n313), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT79), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n560), .A3(new_n553), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(G190), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n552), .A2(G200), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n562), .A2(new_n563), .A3(new_n537), .A4(new_n539), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n557), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n394), .A2(new_n396), .A3(G257), .A4(new_n262), .ZN(new_n566));
  INV_X1    g0366(.A(G303), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(new_n261), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n261), .A2(G264), .A3(G1698), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n256), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n256), .A2(new_n257), .ZN(new_n571));
  INV_X1    g0371(.A(new_n463), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n458), .A2(G270), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n374), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(G97), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n545), .B(new_n211), .C1(G33), .C2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(G116), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G20), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n273), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT20), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n576), .A2(KEYINPUT20), .A3(new_n273), .A4(new_n578), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(KEYINPUT80), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT80), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n579), .A2(new_n584), .A3(new_n580), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n321), .A2(new_n577), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n577), .B1(new_n210), .B2(G33), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n296), .B(new_n587), .C1(new_n319), .C2(new_n320), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n583), .A2(new_n585), .A3(new_n586), .A4(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n574), .A2(new_n589), .A3(KEYINPUT21), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT81), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT81), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n574), .A2(new_n589), .A3(new_n592), .A4(KEYINPUT21), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n261), .A2(new_n211), .A3(G68), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT19), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n211), .B1(new_n336), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(G87), .B2(new_n206), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n596), .B1(new_n274), .B2(new_n575), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n595), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n600), .A2(new_n273), .B1(new_n321), .B2(new_n358), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n484), .A2(G87), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n394), .A2(new_n396), .A3(G244), .A4(G1698), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n394), .A2(new_n396), .A3(G238), .A4(new_n262), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n604), .A3(new_n493), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n256), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n252), .A2(G274), .A3(new_n456), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n210), .A2(G45), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n252), .A2(G250), .A3(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n601), .B(new_n602), .C1(new_n611), .C2(new_n352), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n607), .A2(new_n609), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n256), .B2(new_n605), .ZN(new_n615));
  INV_X1    g0415(.A(G200), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n601), .B1(new_n483), .B2(new_n358), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n611), .A2(G169), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n606), .A2(new_n610), .A3(new_n372), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n613), .A2(new_n618), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n570), .A2(new_n573), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n589), .B1(G200), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n352), .B2(new_n624), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n574), .A2(new_n589), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT21), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n573), .A2(G179), .A3(new_n570), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n627), .A2(new_n628), .B1(new_n629), .B2(new_n589), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n594), .A2(new_n623), .A3(new_n626), .A4(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n565), .A2(new_n631), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n454), .A2(new_n520), .A3(new_n632), .ZN(G372));
  AND2_X1   g0433(.A1(new_n449), .A2(new_n451), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n439), .A2(new_n452), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n376), .A2(new_n373), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n353), .A2(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n637), .A2(new_n350), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n634), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n639), .A2(new_n306), .A3(new_n311), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n315), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n454), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n560), .B1(new_n559), .B2(new_n553), .ZN(new_n644));
  AND4_X1   g0444(.A1(new_n560), .A2(new_n540), .A3(new_n553), .A4(new_n555), .ZN(new_n645));
  OAI211_X1 g0445(.A(KEYINPUT26), .B(new_n623), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n540), .A2(new_n553), .A3(new_n555), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n606), .A2(new_n372), .A3(new_n610), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n374), .B1(new_n606), .B2(new_n610), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT86), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT86), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n620), .A2(new_n651), .A3(new_n621), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n619), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT87), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n615), .B2(new_n616), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n611), .A2(KEYINPUT87), .A3(G200), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n612), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n647), .A2(new_n654), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n646), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n644), .A2(new_n645), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n594), .B(new_n630), .C1(new_n513), .C2(new_n508), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n658), .B1(new_n513), .B2(new_n475), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n664), .A2(new_n665), .A3(new_n564), .A4(new_n666), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n663), .A2(new_n667), .A3(new_n654), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n642), .B1(new_n643), .B2(new_n668), .ZN(G369));
  NAND3_X1  g0469(.A1(new_n210), .A2(new_n211), .A3(G13), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n520), .B1(new_n513), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n518), .B2(new_n676), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n594), .A2(new_n630), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n589), .A2(new_n675), .ZN(new_n680));
  XOR2_X1   g0480(.A(new_n680), .B(KEYINPUT88), .Z(new_n681));
  NAND3_X1  g0481(.A1(new_n679), .A2(new_n626), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n679), .B2(new_n681), .ZN(new_n683));
  XOR2_X1   g0483(.A(KEYINPUT89), .B(G330), .Z(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n678), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n679), .A2(new_n675), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n520), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n516), .A2(new_n517), .A3(new_n676), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT90), .ZN(G399));
  INV_X1    g0495(.A(new_n214), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G1), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n220), .B2(new_n698), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT28), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n663), .A2(new_n667), .A3(new_n654), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT29), .B1(new_n703), .B2(new_n676), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n622), .A2(new_n619), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n617), .B2(new_n612), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n557), .B2(new_n561), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT92), .B1(new_n707), .B2(KEYINPUT26), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n623), .B1(new_n644), .B2(new_n645), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT92), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(new_n710), .A3(new_n661), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n660), .A2(new_n661), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n708), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n654), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n665), .A2(new_n666), .ZN(new_n715));
  INV_X1    g0515(.A(new_n565), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n675), .B1(new_n713), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n704), .B1(KEYINPUT29), .B2(new_n718), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n632), .B(new_n676), .C1(new_n515), .C2(new_n519), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n473), .A2(new_n558), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n615), .A2(new_n372), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n722), .A2(KEYINPUT91), .A3(new_n624), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT91), .B1(new_n722), .B2(new_n624), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n721), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n615), .A2(new_n466), .A3(new_n472), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(new_n554), .A3(new_n629), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n726), .A2(KEYINPUT30), .A3(new_n554), .A4(new_n629), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n725), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n731), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT31), .B1(new_n731), .B2(new_n675), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n720), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n685), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n719), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n702), .B1(new_n738), .B2(G1), .ZN(G364));
  NOR2_X1   g0539(.A1(G13), .A2(G33), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G20), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n683), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(G13), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n210), .B1(new_n746), .B2(G45), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n697), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n696), .A2(new_n398), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n750), .A2(G355), .B1(new_n577), .B2(new_n696), .ZN(new_n751));
  XOR2_X1   g0551(.A(new_n751), .B(KEYINPUT94), .Z(new_n752));
  NOR2_X1   g0552(.A1(new_n248), .A2(new_n455), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n407), .A2(new_n408), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n696), .ZN(new_n756));
  INV_X1    g0556(.A(new_n221), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n756), .B1(new_n757), .B2(G45), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n752), .B1(new_n753), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n217), .B1(G20), .B2(new_n374), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n742), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT95), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n749), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n313), .A2(G200), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT97), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n211), .A2(G190), .ZN(new_n767));
  AND3_X1   g0567(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n766), .B1(new_n765), .B2(new_n767), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n211), .A2(new_n616), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n372), .A2(G190), .A3(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n771), .A2(G77), .B1(G50), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n211), .A2(new_n352), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n765), .A2(new_n776), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT96), .Z(new_n778));
  OAI21_X1  g0578(.A(new_n775), .B1(new_n277), .B2(new_n778), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT98), .Z(new_n780));
  NOR2_X1   g0580(.A1(new_n616), .A2(G179), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n398), .B1(new_n783), .B2(G87), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n767), .A2(new_n781), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n784), .B1(new_n363), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G179), .A2(G200), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n767), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G159), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n787), .A2(G190), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n790), .A2(KEYINPUT32), .B1(G97), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(KEYINPUT32), .B2(new_n790), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n372), .A2(new_n352), .A3(new_n772), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n786), .B(new_n794), .C1(G68), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n780), .A2(new_n797), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n798), .A2(KEYINPUT99), .ZN(new_n799));
  INV_X1    g0599(.A(new_n777), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n800), .A2(G322), .B1(new_n774), .B2(G326), .ZN(new_n801));
  XOR2_X1   g0601(.A(KEYINPUT33), .B(G317), .Z(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n795), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G311), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n770), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n792), .ZN(new_n806));
  INV_X1    g0606(.A(G294), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n785), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n809), .A2(G283), .B1(new_n789), .B2(G329), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n810), .B(new_n398), .C1(new_n567), .C2(new_n782), .ZN(new_n811));
  NOR4_X1   g0611(.A1(new_n803), .A2(new_n805), .A3(new_n808), .A4(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(new_n798), .B2(KEYINPUT99), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n799), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n764), .B1(new_n814), .B2(new_n761), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n744), .B1(new_n815), .B2(KEYINPUT100), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(KEYINPUT100), .B2(new_n815), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n687), .A2(new_n749), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n685), .B2(new_n683), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT93), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n817), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT101), .ZN(G396));
  NAND2_X1  g0624(.A1(new_n636), .A2(KEYINPUT102), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT102), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n376), .B2(new_n373), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(new_n370), .B2(new_n369), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n703), .A2(new_n676), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n668), .A2(new_n675), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n361), .A2(new_n675), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n825), .A2(new_n371), .A3(new_n832), .A4(new_n827), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n636), .A2(new_n675), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n830), .B1(new_n831), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n836), .A2(new_n736), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT103), .Z(new_n838));
  AOI21_X1  g0638(.A(new_n749), .B1(new_n836), .B2(new_n736), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G137), .A2(new_n774), .B1(new_n796), .B2(G150), .ZN(new_n841));
  INV_X1    g0641(.A(G143), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n841), .B1(new_n385), .B2(new_n770), .C1(new_n778), .C2(new_n842), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT34), .Z(new_n844));
  NAND2_X1  g0644(.A1(new_n809), .A2(G68), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n202), .B2(new_n782), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G132), .B2(new_n789), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n847), .B(new_n755), .C1(new_n277), .C2(new_n806), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n261), .B1(new_n783), .B2(G107), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n792), .A2(G97), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n809), .A2(G87), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n789), .A2(G311), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n850), .A2(new_n851), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n800), .A2(G294), .B1(new_n796), .B2(G283), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n567), .B2(new_n773), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n854), .B(new_n856), .C1(G116), .C2(new_n771), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n761), .B1(new_n849), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n749), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n761), .A2(new_n740), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n859), .B1(new_n264), .B2(new_n860), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n858), .B(new_n861), .C1(new_n741), .C2(new_n835), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n840), .A2(new_n862), .ZN(G384));
  NAND2_X1  g0663(.A1(new_n218), .A2(G116), .ZN(new_n864));
  INV_X1    g0664(.A(new_n534), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n864), .B1(new_n865), .B2(KEYINPUT35), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(KEYINPUT35), .B2(new_n865), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT36), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n264), .B(new_n220), .C1(new_n223), .C2(G58), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n392), .A2(G50), .ZN(new_n870));
  OAI211_X1 g0670(.A(G1), .B(new_n745), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT104), .ZN(new_n873));
  INV_X1    g0673(.A(new_n673), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n410), .A2(G68), .B1(new_n387), .B2(new_n390), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n273), .B1(new_n875), .B2(KEYINPUT16), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n413), .B2(new_n405), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n874), .B1(new_n877), .B2(new_n426), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n446), .B1(new_n877), .B2(new_n426), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n878), .A2(new_n879), .A3(new_n437), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT37), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n874), .B1(new_n447), .B2(new_n426), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n437), .A2(new_n448), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n878), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n453), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n885), .A2(new_n887), .A3(KEYINPUT38), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT106), .ZN(new_n889));
  INV_X1    g0689(.A(new_n882), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n437), .A2(new_n448), .A3(new_n882), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT37), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n453), .A2(new_n890), .B1(new_n892), .B2(new_n884), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n888), .B(new_n889), .C1(KEYINPUT38), .C2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n720), .A2(new_n734), .A3(KEYINPUT108), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT108), .B1(new_n720), .B2(new_n734), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n331), .A2(new_n676), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n354), .A2(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n350), .B(new_n353), .C1(new_n331), .C2(new_n676), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n835), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n896), .A2(new_n897), .A3(new_n902), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n884), .A2(new_n881), .B1(new_n453), .B2(new_n886), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n904), .A2(KEYINPUT106), .A3(KEYINPUT38), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n894), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n885), .A2(new_n887), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT40), .B1(new_n909), .B2(new_n888), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n906), .A2(KEYINPUT40), .B1(new_n903), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n896), .A2(new_n897), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n454), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n911), .B(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n914), .A2(new_n684), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n634), .A2(new_n874), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n909), .A2(new_n888), .ZN(new_n917));
  INV_X1    g0717(.A(new_n901), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n828), .A2(new_n676), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n919), .B(KEYINPUT105), .Z(new_n920));
  AOI21_X1  g0720(.A(new_n918), .B1(new_n920), .B2(new_n830), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n916), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n888), .A2(new_n889), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n893), .A2(KEYINPUT38), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n923), .B(new_n905), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n909), .A2(KEYINPUT39), .A3(new_n888), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n350), .A2(new_n675), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n922), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n713), .A2(new_n717), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(KEYINPUT29), .A3(new_n676), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT29), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n668), .B2(new_n675), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n932), .A2(new_n454), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT107), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT107), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n719), .A2(new_n937), .A3(new_n454), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n641), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n930), .B(new_n939), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n915), .A2(new_n940), .B1(new_n210), .B2(new_n746), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n915), .A2(new_n940), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n873), .B1(new_n941), .B2(new_n942), .ZN(G367));
  AOI21_X1  g0743(.A(new_n565), .B1(new_n540), .B2(new_n675), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT109), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n944), .B(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n647), .A2(new_n675), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(new_n520), .A3(new_n689), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT42), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT43), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n676), .B1(new_n601), .B2(new_n602), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n714), .A2(new_n658), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n714), .B2(new_n953), .ZN(new_n955));
  INV_X1    g0755(.A(new_n948), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(new_n518), .ZN(new_n957));
  INV_X1    g0757(.A(new_n664), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n676), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n951), .A2(new_n952), .A3(new_n955), .A4(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n955), .A2(new_n952), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n955), .A2(new_n952), .ZN(new_n962));
  INV_X1    g0762(.A(new_n959), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n961), .B(new_n962), .C1(new_n963), .C2(new_n950), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n688), .A2(new_n956), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n960), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n960), .A2(new_n964), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n688), .B2(new_n956), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n697), .B(KEYINPUT41), .Z(new_n969));
  NAND3_X1  g0769(.A1(new_n956), .A2(KEYINPUT44), .A3(new_n692), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT44), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n693), .B2(new_n948), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n693), .A2(new_n948), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT45), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT45), .B1(new_n693), .B2(new_n948), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n973), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(new_n687), .A3(new_n678), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n976), .A2(new_n977), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n980), .A2(new_n688), .A3(new_n973), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n690), .B1(new_n678), .B2(new_n689), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n687), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n686), .B(new_n690), .C1(new_n678), .C2(new_n689), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n738), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n979), .A2(new_n981), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n969), .B1(new_n988), .B2(new_n738), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n966), .B(new_n968), .C1(new_n989), .C2(new_n748), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n955), .A2(new_n742), .ZN(new_n991));
  INV_X1    g0791(.A(new_n763), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n214), .B2(new_n358), .ZN(new_n993));
  INV_X1    g0793(.A(new_n756), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n994), .A2(new_n241), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n749), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT110), .Z(new_n997));
  INV_X1    g0797(.A(G150), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n777), .A2(new_n998), .B1(new_n795), .B2(new_n385), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(G143), .B2(new_n774), .ZN(new_n1000));
  INV_X1    g0800(.A(G137), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n261), .B1(new_n788), .B2(new_n1001), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n782), .A2(new_n277), .B1(new_n785), .B2(new_n264), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n1002), .B(new_n1003), .C1(G68), .C2(new_n792), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1000), .B(new_n1004), .C1(new_n202), .C2(new_n770), .ZN(new_n1005));
  INV_X1    g0805(.A(G283), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n778), .A2(new_n567), .B1(new_n770), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n783), .A2(G116), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT46), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n1008), .A2(new_n1009), .B1(new_n363), .B2(new_n806), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n1009), .B2(new_n1008), .ZN(new_n1011));
  INV_X1    g0811(.A(G317), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n785), .A2(new_n575), .B1(new_n788), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n755), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n796), .A2(G294), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n774), .A2(G311), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1011), .A2(new_n1014), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1005), .B1(new_n1007), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT47), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n761), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n997), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n991), .A2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT111), .Z(new_n1025));
  NAND2_X1  g0825(.A1(new_n990), .A2(new_n1025), .ZN(G387));
  NAND2_X1  g0826(.A1(new_n985), .A2(new_n748), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n699), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n750), .A2(new_n1028), .B1(new_n363), .B2(new_n696), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n238), .A2(new_n455), .ZN(new_n1030));
  AOI21_X1  g0830(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1031));
  AND3_X1   g0831(.A1(new_n356), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1032));
  AOI21_X1  g0832(.A(KEYINPUT50), .B1(new_n356), .B2(new_n202), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n699), .B(new_n1031), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n756), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1029), .B1(new_n1030), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n859), .B1(new_n1036), .B2(new_n992), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n783), .A2(G77), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n575), .B2(new_n785), .C1(new_n998), .C2(new_n788), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n777), .A2(new_n202), .B1(new_n773), .B2(new_n385), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n806), .A2(new_n358), .ZN(new_n1041));
  NOR4_X1   g0841(.A1(new_n1039), .A2(new_n1040), .A3(new_n754), .A4(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n424), .A2(new_n796), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(new_n392), .C2(new_n770), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT112), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G311), .A2(new_n796), .B1(new_n774), .B2(G322), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n567), .B2(new_n770), .C1(new_n778), .C2(new_n1012), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT48), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n783), .A2(G294), .B1(new_n792), .B2(G283), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT49), .Z(new_n1053));
  OR2_X1    g0853(.A1(new_n1053), .A2(KEYINPUT113), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n789), .A2(G326), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n754), .B(new_n1055), .C1(new_n577), .C2(new_n785), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n1053), .B2(KEYINPUT113), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1045), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1037), .B1(new_n678), .B2(new_n743), .C1(new_n1058), .C2(new_n1021), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n986), .A2(new_n697), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n985), .A2(new_n738), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1027), .B(new_n1059), .C1(new_n1060), .C2(new_n1061), .ZN(G393));
  INV_X1    g0862(.A(new_n981), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n688), .B1(new_n980), .B2(new_n973), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n986), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1065), .A2(new_n697), .A3(new_n988), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n994), .A2(new_n245), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n992), .B1(new_n575), .B2(new_n214), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n795), .A2(new_n567), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G283), .A2(new_n783), .B1(new_n789), .B2(G322), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1070), .B(new_n398), .C1(new_n363), .C2(new_n785), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1069), .B(new_n1071), .C1(G116), .C2(new_n792), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n777), .A2(new_n804), .B1(new_n773), .B2(new_n1012), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT52), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1072), .B(new_n1074), .C1(new_n807), .C2(new_n770), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n792), .A2(G77), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n755), .A2(new_n1076), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n852), .B1(new_n842), .B2(new_n788), .C1(new_n224), .C2(new_n782), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(G50), .C2(new_n796), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n777), .A2(new_n385), .B1(new_n773), .B2(new_n998), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT51), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n771), .A2(new_n356), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1075), .A2(new_n1083), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n749), .B1(new_n1067), .B2(new_n1068), .C1(new_n1084), .C2(new_n1021), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n956), .B2(new_n742), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1086), .B1(new_n1087), .B2(new_n748), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1066), .A2(new_n1088), .ZN(G390));
  NAND4_X1  g0889(.A1(new_n735), .A2(new_n685), .A3(new_n835), .A4(new_n901), .ZN(new_n1090));
  AND4_X1   g0890(.A1(KEYINPUT106), .A2(new_n885), .A3(KEYINPUT38), .A4(new_n887), .ZN(new_n1091));
  AOI21_X1  g0891(.A(KEYINPUT106), .B1(new_n904), .B2(KEYINPUT38), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n453), .A2(new_n890), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n892), .A2(new_n884), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n908), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1091), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n718), .A2(new_n829), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n919), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n901), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1096), .A2(new_n1099), .A3(new_n929), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n888), .ZN(new_n1101));
  AOI21_X1  g0901(.A(KEYINPUT38), .B1(new_n885), .B2(new_n887), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n1101), .A2(new_n1102), .A3(new_n923), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n1096), .B2(new_n923), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n929), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n921), .A2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1090), .B(new_n1100), .C1(new_n1104), .C2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT108), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n735), .A2(new_n1108), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n901), .A2(new_n835), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1109), .A2(G330), .A3(new_n895), .A4(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1106), .B1(new_n926), .B2(new_n927), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n929), .B(new_n905), .C1(new_n924), .C2(new_n925), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n918), .B1(new_n1097), .B2(new_n919), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1112), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1107), .A2(new_n748), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n860), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n749), .B1(new_n424), .B2(new_n1119), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n770), .A2(new_n575), .B1(new_n363), .B2(new_n795), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1121), .A2(KEYINPUT116), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(KEYINPUT116), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n261), .B1(new_n783), .B2(G87), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n789), .A2(G294), .ZN(new_n1125));
  AND4_X1   g0925(.A1(new_n845), .A2(new_n1124), .A3(new_n1076), .A4(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n800), .A2(G116), .B1(new_n774), .B2(G283), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1122), .A2(new_n1123), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT117), .ZN(new_n1129));
  OR2_X1    g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(G125), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n261), .B1(new_n788), .B2(new_n1131), .C1(new_n202), .C2(new_n785), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n782), .A2(new_n998), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT115), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1134), .A2(KEYINPUT53), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1132), .B(new_n1135), .C1(G159), .C2(new_n792), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1134), .A2(KEYINPUT53), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT54), .B(G143), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n771), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(G128), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n1141), .A2(new_n773), .B1(new_n795), .B2(new_n1001), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G132), .B2(new_n800), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1136), .A2(new_n1137), .A3(new_n1140), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1130), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1120), .B1(new_n1146), .B2(new_n761), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT118), .Z(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n1104), .B2(new_n741), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1118), .A2(KEYINPUT119), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT119), .B1(new_n1118), .B2(new_n1149), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n912), .A2(G330), .A3(new_n454), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n937), .B1(new_n719), .B2(new_n454), .ZN(new_n1154));
  AND4_X1   g0954(.A1(new_n937), .A2(new_n932), .A3(new_n454), .A4(new_n934), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n642), .B(new_n1153), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1109), .A2(G330), .A3(new_n835), .A4(new_n895), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n918), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1097), .A2(new_n919), .A3(new_n1090), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n735), .A2(new_n685), .A3(new_n835), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n918), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1111), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n920), .A2(new_n830), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1158), .A2(new_n1159), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1156), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1107), .A2(new_n1165), .A3(new_n1117), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n1166), .A2(new_n697), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT114), .ZN(new_n1168));
  AND4_X1   g0968(.A1(G330), .A2(new_n454), .A3(new_n1109), .A4(new_n895), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n641), .B(new_n1169), .C1(new_n936), .C2(new_n938), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1159), .A2(new_n1158), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AOI221_X4 g0973(.A(new_n1168), .B1(new_n1170), .B2(new_n1173), .C1(new_n1107), .C2(new_n1117), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1107), .A2(new_n1117), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1165), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT114), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1167), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1152), .A2(new_n1178), .ZN(G378));
  NOR2_X1   g0979(.A1(new_n785), .A2(new_n277), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT120), .Z(new_n1181));
  OAI221_X1 g0981(.A(new_n1181), .B1(new_n575), .B2(new_n795), .C1(new_n577), .C2(new_n773), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n754), .A2(new_n251), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1038), .B1(new_n1006), .B2(new_n788), .C1(new_n392), .C2(new_n806), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n800), .A2(G107), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT121), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1185), .B(new_n1187), .C1(new_n358), .C2(new_n770), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT58), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1183), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n806), .A2(new_n998), .B1(new_n1138), .B2(new_n782), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n796), .B2(G132), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n1131), .B2(new_n773), .C1(new_n1141), .C2(new_n777), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G137), .B2(new_n771), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT122), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n250), .B(new_n251), .C1(new_n785), .C2(new_n385), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(G124), .C2(new_n789), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1190), .B(new_n1193), .C1(new_n1199), .C2(new_n1202), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n749), .B1(G50), .B2(new_n1119), .C1(new_n1203), .C2(new_n1021), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n673), .B1(new_n291), .B2(new_n300), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n316), .B(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT123), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1209), .A2(KEYINPUT123), .A3(new_n1210), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n741), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1204), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1209), .A2(KEYINPUT124), .A3(new_n1210), .ZN(new_n1217));
  INV_X1    g1017(.A(G330), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1217), .B1(new_n911), .B2(new_n1218), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1209), .A2(KEYINPUT123), .A3(KEYINPUT124), .A4(new_n1210), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1213), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT40), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n1096), .B2(new_n903), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n910), .A2(new_n903), .ZN(new_n1224));
  OAI211_X1 g1024(.A(G330), .B(new_n1221), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1219), .A2(new_n1225), .A3(new_n930), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n930), .B1(new_n1219), .B2(new_n1225), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1216), .B1(new_n1228), .B2(new_n748), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT125), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1156), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT125), .B1(new_n939), .B2(new_n1153), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1166), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT57), .B1(new_n1228), .B2(new_n1234), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1234), .B(KEYINPUT57), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n697), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1229), .B1(new_n1235), .B2(new_n1237), .ZN(G375));
  NAND2_X1  g1038(.A1(new_n918), .A2(new_n740), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n749), .B1(G68), .B2(new_n1119), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n777), .A2(new_n1006), .B1(new_n795), .B2(new_n577), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(G294), .B2(new_n774), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n398), .B1(new_n785), .B2(new_n264), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n782), .A2(new_n575), .B1(new_n788), .B2(new_n567), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1041), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1242), .B(new_n1245), .C1(new_n363), .C2(new_n770), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1181), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G132), .B2(new_n774), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n792), .A2(G50), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n782), .A2(new_n385), .B1(new_n788), .B2(new_n1141), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n754), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n796), .A2(new_n1139), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1248), .A2(new_n1249), .A3(new_n1251), .A4(new_n1252), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n778), .A2(new_n1001), .B1(new_n770), .B2(new_n998), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1246), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1240), .B1(new_n1255), .B2(new_n761), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1173), .A2(new_n748), .B1(new_n1239), .B2(new_n1256), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1165), .A2(new_n969), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1156), .A2(new_n1164), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1257), .B1(new_n1259), .B2(new_n1260), .ZN(G381));
  OR4_X1    g1061(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1262), .A2(G387), .A3(G381), .ZN(new_n1263));
  INV_X1    g1063(.A(G375), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1118), .A2(new_n1149), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1178), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1263), .A2(new_n1264), .A3(new_n1266), .ZN(G407));
  NAND2_X1  g1067(.A1(new_n674), .A2(G213), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1264), .A2(new_n1266), .A3(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(G407), .A2(new_n1270), .A3(G213), .ZN(G409));
  INV_X1    g1071(.A(KEYINPUT61), .ZN(new_n1272));
  OAI211_X1 g1072(.A(G378), .B(new_n1229), .C1(new_n1235), .C2(new_n1237), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n969), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1234), .B(new_n1274), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1216), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1275), .B(new_n1276), .C1(new_n747), .C2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1266), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1269), .B1(new_n1273), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1260), .A2(KEYINPUT60), .ZN(new_n1281));
  XOR2_X1   g1081(.A(KEYINPUT126), .B(KEYINPUT60), .Z(new_n1282));
  NOR2_X1   g1082(.A1(new_n1165), .A2(new_n1282), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1281), .B(new_n697), .C1(new_n1283), .C2(new_n1260), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1257), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT127), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G384), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(G384), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(KEYINPUT127), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1285), .A2(new_n1287), .A3(new_n1289), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1284), .A2(new_n1288), .A3(KEYINPUT127), .A4(new_n1257), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1269), .A2(G2897), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1290), .A2(G2897), .A3(new_n1269), .A4(new_n1291), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1272), .B1(new_n1280), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1280), .A2(new_n1292), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT63), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  XOR2_X1   g1101(.A(G396), .B(G393), .Z(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n990), .A2(G390), .A3(new_n1025), .ZN(new_n1304));
  AOI21_X1  g1104(.A(G390), .B1(new_n990), .B2(new_n1025), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1303), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(G390), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(G387), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n990), .A2(G390), .A3(new_n1025), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1308), .A2(new_n1302), .A3(new_n1309), .ZN(new_n1310));
  AND2_X1   g1110(.A1(new_n1306), .A2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1280), .A2(KEYINPUT63), .A3(new_n1292), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1298), .A2(new_n1301), .A3(new_n1311), .A4(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT62), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1280), .A2(new_n1314), .A3(new_n1292), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1314), .B1(new_n1280), .B2(new_n1292), .ZN(new_n1316));
  NOR3_X1   g1116(.A1(new_n1315), .A2(new_n1297), .A3(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1313), .B1(new_n1317), .B2(new_n1311), .ZN(G405));
  NAND2_X1  g1118(.A1(G375), .A2(new_n1266), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1273), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1311), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1292), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1306), .A2(new_n1310), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1323), .A2(new_n1273), .A3(new_n1319), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1321), .A2(new_n1322), .A3(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1322), .B1(new_n1321), .B2(new_n1324), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(G402));
endmodule


