

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U552 ( .A1(n601), .A2(n600), .ZN(n988) );
  NOR2_X2 U553 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X2 U554 ( .A1(n758), .A2(n757), .ZN(n780) );
  XNOR2_X2 U555 ( .A(n525), .B(KEYINPUT66), .ZN(n531) );
  BUF_X1 U556 ( .A(n701), .Z(n742) );
  INV_X2 U557 ( .A(n701), .ZN(n715) );
  XNOR2_X1 U558 ( .A(n710), .B(n709), .ZN(n712) );
  XNOR2_X1 U559 ( .A(n706), .B(KEYINPUT31), .ZN(n707) );
  NOR2_X2 U560 ( .A1(n531), .A2(n530), .ZN(n694) );
  XOR2_X1 U561 ( .A(n789), .B(KEYINPUT106), .Z(n518) );
  XNOR2_X1 U562 ( .A(KEYINPUT98), .B(KEYINPUT27), .ZN(n709) );
  NOR2_X1 U563 ( .A1(n718), .A2(n717), .ZN(n719) );
  OR2_X1 U564 ( .A1(n971), .A2(n719), .ZN(n725) );
  NAND2_X1 U565 ( .A1(n732), .A2(n731), .ZN(n734) );
  AND2_X1 U566 ( .A1(n700), .A2(n699), .ZN(n705) );
  NOR2_X1 U567 ( .A1(n783), .A2(G1966), .ZN(n756) );
  INV_X1 U568 ( .A(n830), .ZN(n818) );
  XNOR2_X1 U569 ( .A(KEYINPUT23), .B(KEYINPUT65), .ZN(n519) );
  INV_X1 U570 ( .A(G651), .ZN(n539) );
  NAND2_X1 U571 ( .A1(n654), .A2(G56), .ZN(n598) );
  INV_X1 U572 ( .A(G2105), .ZN(n522) );
  NOR2_X1 U573 ( .A1(G651), .A2(n641), .ZN(n659) );
  NOR2_X2 U574 ( .A1(G2104), .A2(n522), .ZN(n892) );
  BUF_X1 U575 ( .A(n694), .Z(G160) );
  XNOR2_X1 U576 ( .A(n519), .B(KEYINPUT64), .ZN(n521) );
  AND2_X1 U577 ( .A1(n522), .A2(G2104), .ZN(n549) );
  NAND2_X1 U578 ( .A1(G101), .A2(n549), .ZN(n520) );
  XNOR2_X1 U579 ( .A(n521), .B(n520), .ZN(n524) );
  NAND2_X1 U580 ( .A1(n892), .A2(G125), .ZN(n523) );
  NAND2_X1 U581 ( .A1(n524), .A2(n523), .ZN(n525) );
  AND2_X1 U582 ( .A1(G2105), .A2(G2104), .ZN(n891) );
  NAND2_X1 U583 ( .A1(G113), .A2(n891), .ZN(n529) );
  XNOR2_X1 U584 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n527) );
  NOR2_X1 U585 ( .A1(G2105), .A2(G2104), .ZN(n526) );
  XNOR2_X2 U586 ( .A(n527), .B(n526), .ZN(n888) );
  NAND2_X1 U587 ( .A1(G137), .A2(n888), .ZN(n528) );
  NAND2_X1 U588 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U589 ( .A(G543), .B(KEYINPUT0), .Z(n641) );
  NAND2_X1 U590 ( .A1(G51), .A2(n659), .ZN(n535) );
  NOR2_X1 U591 ( .A1(G543), .A2(n539), .ZN(n532) );
  XOR2_X1 U592 ( .A(KEYINPUT1), .B(n532), .Z(n533) );
  XNOR2_X2 U593 ( .A(KEYINPUT68), .B(n533), .ZN(n654) );
  NAND2_X1 U594 ( .A1(G63), .A2(n654), .ZN(n534) );
  NAND2_X1 U595 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U596 ( .A(KEYINPUT6), .B(n536), .ZN(n544) );
  NOR2_X1 U597 ( .A1(G543), .A2(G651), .ZN(n658) );
  NAND2_X1 U598 ( .A1(G89), .A2(n658), .ZN(n537) );
  XNOR2_X1 U599 ( .A(n537), .B(KEYINPUT74), .ZN(n538) );
  XNOR2_X1 U600 ( .A(n538), .B(KEYINPUT4), .ZN(n541) );
  NOR2_X1 U601 ( .A1(n641), .A2(n539), .ZN(n652) );
  NAND2_X1 U602 ( .A1(G76), .A2(n652), .ZN(n540) );
  NAND2_X1 U603 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U604 ( .A(n542), .B(KEYINPUT5), .Z(n543) );
  NOR2_X1 U605 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U606 ( .A(KEYINPUT7), .B(n545), .Z(n547) );
  XOR2_X1 U607 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n546) );
  XNOR2_X1 U608 ( .A(n547), .B(n546), .ZN(G168) );
  NAND2_X1 U609 ( .A1(n891), .A2(G114), .ZN(n548) );
  XNOR2_X1 U610 ( .A(n548), .B(KEYINPUT92), .ZN(n552) );
  INV_X1 U611 ( .A(n549), .ZN(n550) );
  INV_X1 U612 ( .A(n550), .ZN(n887) );
  NAND2_X1 U613 ( .A1(G102), .A2(n887), .ZN(n551) );
  NAND2_X1 U614 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U615 ( .A1(G138), .A2(n888), .ZN(n554) );
  NAND2_X1 U616 ( .A1(G126), .A2(n892), .ZN(n553) );
  NAND2_X1 U617 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U618 ( .A1(n556), .A2(n555), .ZN(G164) );
  NAND2_X1 U619 ( .A1(G85), .A2(n658), .ZN(n558) );
  NAND2_X1 U620 ( .A1(G72), .A2(n652), .ZN(n557) );
  NAND2_X1 U621 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U622 ( .A1(G47), .A2(n659), .ZN(n560) );
  NAND2_X1 U623 ( .A1(G60), .A2(n654), .ZN(n559) );
  NAND2_X1 U624 ( .A1(n560), .A2(n559), .ZN(n561) );
  OR2_X1 U625 ( .A1(n562), .A2(n561), .ZN(G290) );
  XOR2_X1 U626 ( .A(G2430), .B(G2451), .Z(n564) );
  XNOR2_X1 U627 ( .A(KEYINPUT111), .B(G2443), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n564), .B(n563), .ZN(n571) );
  XOR2_X1 U629 ( .A(G2435), .B(G2446), .Z(n566) );
  XNOR2_X1 U630 ( .A(G2427), .B(G2454), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(n567) );
  XOR2_X1 U632 ( .A(n567), .B(G2438), .Z(n569) );
  XNOR2_X1 U633 ( .A(G1348), .B(G1341), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n571), .B(n570), .ZN(n572) );
  AND2_X1 U636 ( .A1(n572), .A2(G14), .ZN(G401) );
  NAND2_X1 U637 ( .A1(G52), .A2(n659), .ZN(n574) );
  NAND2_X1 U638 ( .A1(G64), .A2(n654), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n579) );
  NAND2_X1 U640 ( .A1(G90), .A2(n658), .ZN(n576) );
  NAND2_X1 U641 ( .A1(G77), .A2(n652), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U643 ( .A(KEYINPUT9), .B(n577), .Z(n578) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(G171) );
  AND2_X1 U645 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U646 ( .A1(G123), .A2(n892), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n580), .B(KEYINPUT18), .ZN(n587) );
  NAND2_X1 U648 ( .A1(G111), .A2(n891), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G99), .A2(n887), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U651 ( .A1(G135), .A2(n888), .ZN(n583) );
  XNOR2_X1 U652 ( .A(KEYINPUT77), .B(n583), .ZN(n584) );
  NOR2_X1 U653 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n587), .A2(n586), .ZN(n923) );
  XNOR2_X1 U655 ( .A(G2096), .B(n923), .ZN(n588) );
  OR2_X1 U656 ( .A1(G2100), .A2(n588), .ZN(G156) );
  INV_X1 U657 ( .A(G132), .ZN(G219) );
  INV_X1 U658 ( .A(G82), .ZN(G220) );
  INV_X1 U659 ( .A(G57), .ZN(G237) );
  INV_X1 U660 ( .A(G69), .ZN(G235) );
  INV_X1 U661 ( .A(G108), .ZN(G238) );
  INV_X1 U662 ( .A(G120), .ZN(G236) );
  XOR2_X1 U663 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U664 ( .A1(G7), .A2(G661), .ZN(n589) );
  XNOR2_X1 U665 ( .A(n589), .B(KEYINPUT10), .ZN(n590) );
  XNOR2_X1 U666 ( .A(KEYINPUT70), .B(n590), .ZN(G223) );
  INV_X1 U667 ( .A(G223), .ZN(n840) );
  NAND2_X1 U668 ( .A1(n840), .A2(G567), .ZN(n591) );
  XOR2_X1 U669 ( .A(KEYINPUT11), .B(n591), .Z(G234) );
  NAND2_X1 U670 ( .A1(n658), .A2(G81), .ZN(n592) );
  XNOR2_X1 U671 ( .A(n592), .B(KEYINPUT12), .ZN(n594) );
  NAND2_X1 U672 ( .A1(G68), .A2(n652), .ZN(n593) );
  NAND2_X1 U673 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U674 ( .A(n595), .B(KEYINPUT13), .ZN(n597) );
  NAND2_X1 U675 ( .A1(G43), .A2(n659), .ZN(n596) );
  NAND2_X1 U676 ( .A1(n597), .A2(n596), .ZN(n601) );
  XNOR2_X1 U677 ( .A(n598), .B(KEYINPUT14), .ZN(n599) );
  XNOR2_X1 U678 ( .A(n599), .B(KEYINPUT71), .ZN(n600) );
  NAND2_X1 U679 ( .A1(n988), .A2(G860), .ZN(G153) );
  XOR2_X1 U680 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  INV_X1 U681 ( .A(G868), .ZN(n674) );
  NOR2_X1 U682 ( .A1(G301), .A2(n674), .ZN(n610) );
  NAND2_X1 U683 ( .A1(G92), .A2(n658), .ZN(n603) );
  NAND2_X1 U684 ( .A1(G79), .A2(n652), .ZN(n602) );
  NAND2_X1 U685 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U686 ( .A1(G54), .A2(n659), .ZN(n605) );
  NAND2_X1 U687 ( .A1(G66), .A2(n654), .ZN(n604) );
  NAND2_X1 U688 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U689 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U690 ( .A(KEYINPUT15), .B(n608), .Z(n971) );
  AND2_X1 U691 ( .A1(n674), .A2(n971), .ZN(n609) );
  NOR2_X1 U692 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U693 ( .A(KEYINPUT73), .B(n611), .Z(G284) );
  NAND2_X1 U694 ( .A1(G53), .A2(n659), .ZN(n613) );
  NAND2_X1 U695 ( .A1(G65), .A2(n654), .ZN(n612) );
  NAND2_X1 U696 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U697 ( .A1(G91), .A2(n658), .ZN(n615) );
  NAND2_X1 U698 ( .A1(G78), .A2(n652), .ZN(n614) );
  NAND2_X1 U699 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U700 ( .A1(n617), .A2(n616), .ZN(n972) );
  XNOR2_X1 U701 ( .A(n972), .B(KEYINPUT69), .ZN(G299) );
  NAND2_X1 U702 ( .A1(G868), .A2(G286), .ZN(n619) );
  NAND2_X1 U703 ( .A1(G299), .A2(n674), .ZN(n618) );
  NAND2_X1 U704 ( .A1(n619), .A2(n618), .ZN(G297) );
  INV_X1 U705 ( .A(G860), .ZN(n620) );
  NAND2_X1 U706 ( .A1(n620), .A2(G559), .ZN(n621) );
  NAND2_X1 U707 ( .A1(n621), .A2(n971), .ZN(n622) );
  XNOR2_X1 U708 ( .A(n622), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U709 ( .A1(n971), .A2(G868), .ZN(n623) );
  NOR2_X1 U710 ( .A1(G559), .A2(n623), .ZN(n625) );
  AND2_X1 U711 ( .A1(n674), .A2(n988), .ZN(n624) );
  NOR2_X1 U712 ( .A1(n625), .A2(n624), .ZN(G282) );
  NAND2_X1 U713 ( .A1(G559), .A2(n971), .ZN(n626) );
  XNOR2_X1 U714 ( .A(n626), .B(n988), .ZN(n671) );
  XOR2_X1 U715 ( .A(n671), .B(KEYINPUT78), .Z(n627) );
  NOR2_X1 U716 ( .A1(G860), .A2(n627), .ZN(n628) );
  XOR2_X1 U717 ( .A(KEYINPUT80), .B(n628), .Z(n636) );
  NAND2_X1 U718 ( .A1(G55), .A2(n659), .ZN(n630) );
  NAND2_X1 U719 ( .A1(G67), .A2(n654), .ZN(n629) );
  NAND2_X1 U720 ( .A1(n630), .A2(n629), .ZN(n635) );
  NAND2_X1 U721 ( .A1(G93), .A2(n658), .ZN(n632) );
  NAND2_X1 U722 ( .A1(G80), .A2(n652), .ZN(n631) );
  NAND2_X1 U723 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U724 ( .A(KEYINPUT79), .B(n633), .Z(n634) );
  NOR2_X1 U725 ( .A1(n635), .A2(n634), .ZN(n673) );
  XOR2_X1 U726 ( .A(n636), .B(n673), .Z(G145) );
  NAND2_X1 U727 ( .A1(G49), .A2(n659), .ZN(n638) );
  NAND2_X1 U728 ( .A1(G74), .A2(G651), .ZN(n637) );
  NAND2_X1 U729 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U730 ( .A(KEYINPUT81), .B(n639), .Z(n640) );
  NOR2_X1 U731 ( .A1(n654), .A2(n640), .ZN(n643) );
  NAND2_X1 U732 ( .A1(n641), .A2(G87), .ZN(n642) );
  NAND2_X1 U733 ( .A1(n643), .A2(n642), .ZN(G288) );
  XOR2_X1 U734 ( .A(KEYINPUT82), .B(KEYINPUT2), .Z(n645) );
  NAND2_X1 U735 ( .A1(G73), .A2(n652), .ZN(n644) );
  XNOR2_X1 U736 ( .A(n645), .B(n644), .ZN(n649) );
  NAND2_X1 U737 ( .A1(G86), .A2(n658), .ZN(n647) );
  NAND2_X1 U738 ( .A1(G48), .A2(n659), .ZN(n646) );
  NAND2_X1 U739 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U740 ( .A1(n649), .A2(n648), .ZN(n651) );
  NAND2_X1 U741 ( .A1(G61), .A2(n654), .ZN(n650) );
  NAND2_X1 U742 ( .A1(n651), .A2(n650), .ZN(G305) );
  NAND2_X1 U743 ( .A1(G75), .A2(n652), .ZN(n653) );
  XNOR2_X1 U744 ( .A(n653), .B(KEYINPUT84), .ZN(n657) );
  NAND2_X1 U745 ( .A1(n654), .A2(G62), .ZN(n655) );
  XOR2_X1 U746 ( .A(KEYINPUT83), .B(n655), .Z(n656) );
  NAND2_X1 U747 ( .A1(n657), .A2(n656), .ZN(n663) );
  NAND2_X1 U748 ( .A1(G88), .A2(n658), .ZN(n661) );
  NAND2_X1 U749 ( .A1(G50), .A2(n659), .ZN(n660) );
  NAND2_X1 U750 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U751 ( .A1(n663), .A2(n662), .ZN(G166) );
  XNOR2_X1 U752 ( .A(KEYINPUT86), .B(KEYINPUT19), .ZN(n665) );
  XNOR2_X1 U753 ( .A(G290), .B(KEYINPUT85), .ZN(n664) );
  XNOR2_X1 U754 ( .A(n665), .B(n664), .ZN(n668) );
  XNOR2_X1 U755 ( .A(n673), .B(G288), .ZN(n666) );
  XNOR2_X1 U756 ( .A(n666), .B(G299), .ZN(n667) );
  XNOR2_X1 U757 ( .A(n668), .B(n667), .ZN(n670) );
  XNOR2_X1 U758 ( .A(G305), .B(G166), .ZN(n669) );
  XNOR2_X1 U759 ( .A(n670), .B(n669), .ZN(n908) );
  XOR2_X1 U760 ( .A(n908), .B(n671), .Z(n672) );
  NOR2_X1 U761 ( .A1(n674), .A2(n672), .ZN(n676) );
  AND2_X1 U762 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U763 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U764 ( .A1(G2084), .A2(G2078), .ZN(n677) );
  XOR2_X1 U765 ( .A(KEYINPUT20), .B(n677), .Z(n678) );
  NAND2_X1 U766 ( .A1(G2090), .A2(n678), .ZN(n680) );
  XOR2_X1 U767 ( .A(KEYINPUT87), .B(KEYINPUT21), .Z(n679) );
  XNOR2_X1 U768 ( .A(n680), .B(n679), .ZN(n681) );
  NAND2_X1 U769 ( .A1(G2072), .A2(n681), .ZN(G158) );
  XNOR2_X1 U770 ( .A(KEYINPUT88), .B(G44), .ZN(n682) );
  XNOR2_X1 U771 ( .A(n682), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U772 ( .A1(G236), .A2(G238), .ZN(n684) );
  NOR2_X1 U773 ( .A1(G235), .A2(G237), .ZN(n683) );
  NAND2_X1 U774 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U775 ( .A(KEYINPUT90), .B(n685), .ZN(n845) );
  NAND2_X1 U776 ( .A1(G567), .A2(n845), .ZN(n691) );
  NOR2_X1 U777 ( .A1(G220), .A2(G219), .ZN(n686) );
  XOR2_X1 U778 ( .A(KEYINPUT22), .B(n686), .Z(n687) );
  NOR2_X1 U779 ( .A1(G218), .A2(n687), .ZN(n688) );
  NAND2_X1 U780 ( .A1(G96), .A2(n688), .ZN(n844) );
  NAND2_X1 U781 ( .A1(G2106), .A2(n844), .ZN(n689) );
  XOR2_X1 U782 ( .A(KEYINPUT89), .B(n689), .Z(n690) );
  NAND2_X1 U783 ( .A1(n691), .A2(n690), .ZN(n920) );
  NAND2_X1 U784 ( .A1(G483), .A2(G661), .ZN(n692) );
  NOR2_X1 U785 ( .A1(n920), .A2(n692), .ZN(n693) );
  XOR2_X1 U786 ( .A(KEYINPUT91), .B(n693), .Z(n843) );
  NAND2_X1 U787 ( .A1(n843), .A2(G36), .ZN(G176) );
  XNOR2_X1 U788 ( .A(KEYINPUT93), .B(G166), .ZN(G303) );
  NAND2_X1 U789 ( .A1(n694), .A2(G40), .ZN(n806) );
  INV_X1 U790 ( .A(n806), .ZN(n695) );
  NOR2_X1 U791 ( .A1(G164), .A2(G1384), .ZN(n807) );
  NAND2_X1 U792 ( .A1(n695), .A2(n807), .ZN(n701) );
  NAND2_X1 U793 ( .A1(n701), .A2(G8), .ZN(n696) );
  XOR2_X1 U794 ( .A(KEYINPUT96), .B(n696), .Z(n776) );
  INV_X1 U795 ( .A(n776), .ZN(n783) );
  NOR2_X1 U796 ( .A1(G2084), .A2(n742), .ZN(n752) );
  NOR2_X1 U797 ( .A1(n756), .A2(n752), .ZN(n697) );
  AND2_X1 U798 ( .A1(n697), .A2(G8), .ZN(n698) );
  XNOR2_X1 U799 ( .A(n698), .B(KEYINPUT30), .ZN(n700) );
  INV_X1 U800 ( .A(G168), .ZN(n699) );
  XNOR2_X1 U801 ( .A(G1961), .B(KEYINPUT97), .ZN(n1006) );
  NAND2_X1 U802 ( .A1(n742), .A2(n1006), .ZN(n703) );
  XNOR2_X1 U803 ( .A(G2078), .B(KEYINPUT25), .ZN(n957) );
  NAND2_X1 U804 ( .A1(n715), .A2(n957), .ZN(n702) );
  NAND2_X1 U805 ( .A1(n703), .A2(n702), .ZN(n735) );
  NOR2_X1 U806 ( .A1(G171), .A2(n735), .ZN(n704) );
  NOR2_X2 U807 ( .A1(n705), .A2(n704), .ZN(n708) );
  INV_X1 U808 ( .A(KEYINPUT102), .ZN(n706) );
  XNOR2_X1 U809 ( .A(n708), .B(n707), .ZN(n740) );
  NAND2_X1 U810 ( .A1(G2072), .A2(n715), .ZN(n710) );
  INV_X1 U811 ( .A(G1956), .ZN(n997) );
  NOR2_X1 U812 ( .A1(n715), .A2(n997), .ZN(n711) );
  NOR2_X1 U813 ( .A1(n712), .A2(n711), .ZN(n728) );
  NAND2_X1 U814 ( .A1(n728), .A2(n972), .ZN(n727) );
  NAND2_X1 U815 ( .A1(n742), .A2(G1341), .ZN(n713) );
  XNOR2_X1 U816 ( .A(n713), .B(KEYINPUT100), .ZN(n714) );
  NAND2_X1 U817 ( .A1(n714), .A2(n988), .ZN(n718) );
  NAND2_X1 U818 ( .A1(G1996), .A2(n715), .ZN(n716) );
  XOR2_X1 U819 ( .A(KEYINPUT26), .B(n716), .Z(n717) );
  NAND2_X1 U820 ( .A1(n719), .A2(n971), .ZN(n723) );
  NAND2_X1 U821 ( .A1(G1348), .A2(n742), .ZN(n721) );
  NAND2_X1 U822 ( .A1(G2067), .A2(n715), .ZN(n720) );
  NAND2_X1 U823 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U824 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U825 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U826 ( .A1(n727), .A2(n726), .ZN(n732) );
  NOR2_X1 U827 ( .A1(n728), .A2(n972), .ZN(n730) );
  XNOR2_X1 U828 ( .A(KEYINPUT99), .B(KEYINPUT28), .ZN(n729) );
  XNOR2_X1 U829 ( .A(n730), .B(n729), .ZN(n731) );
  INV_X1 U830 ( .A(KEYINPUT29), .ZN(n733) );
  XNOR2_X1 U831 ( .A(n734), .B(n733), .ZN(n737) );
  NAND2_X1 U832 ( .A1(G171), .A2(n735), .ZN(n736) );
  AND2_X1 U833 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U834 ( .A(n738), .B(KEYINPUT101), .ZN(n739) );
  NAND2_X1 U835 ( .A1(n740), .A2(n739), .ZN(n754) );
  AND2_X1 U836 ( .A1(G286), .A2(G8), .ZN(n741) );
  NAND2_X1 U837 ( .A1(n754), .A2(n741), .ZN(n750) );
  INV_X1 U838 ( .A(G8), .ZN(n748) );
  NOR2_X1 U839 ( .A1(n783), .A2(G1971), .ZN(n744) );
  NOR2_X1 U840 ( .A1(G2090), .A2(n742), .ZN(n743) );
  NOR2_X1 U841 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U842 ( .A(KEYINPUT103), .B(n745), .Z(n746) );
  NAND2_X1 U843 ( .A1(n746), .A2(G303), .ZN(n747) );
  OR2_X1 U844 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U845 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U846 ( .A(n751), .B(KEYINPUT32), .ZN(n758) );
  NAND2_X1 U847 ( .A1(G8), .A2(n752), .ZN(n753) );
  NAND2_X1 U848 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U849 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n761) );
  NOR2_X1 U851 ( .A1(G1971), .A2(G303), .ZN(n759) );
  OR2_X1 U852 ( .A1(n761), .A2(n759), .ZN(n992) );
  NOR2_X1 U853 ( .A1(n780), .A2(n992), .ZN(n760) );
  NOR2_X1 U854 ( .A1(n783), .A2(n760), .ZN(n768) );
  NAND2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n980) );
  INV_X1 U856 ( .A(KEYINPUT33), .ZN(n770) );
  NAND2_X1 U857 ( .A1(n761), .A2(n776), .ZN(n762) );
  NOR2_X1 U858 ( .A1(n770), .A2(n762), .ZN(n763) );
  XOR2_X1 U859 ( .A(n763), .B(KEYINPUT104), .Z(n769) );
  AND2_X1 U860 ( .A1(n980), .A2(n769), .ZN(n766) );
  OR2_X1 U861 ( .A1(G1981), .A2(G305), .ZN(n775) );
  NAND2_X1 U862 ( .A1(G1981), .A2(G305), .ZN(n764) );
  NAND2_X1 U863 ( .A1(n775), .A2(n764), .ZN(n983) );
  INV_X1 U864 ( .A(n983), .ZN(n765) );
  AND2_X1 U865 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U866 ( .A1(n768), .A2(n767), .ZN(n774) );
  INV_X1 U867 ( .A(n769), .ZN(n771) );
  OR2_X1 U868 ( .A1(n771), .A2(n770), .ZN(n772) );
  OR2_X1 U869 ( .A1(n983), .A2(n772), .ZN(n773) );
  NAND2_X1 U870 ( .A1(n774), .A2(n773), .ZN(n788) );
  XOR2_X1 U871 ( .A(KEYINPUT24), .B(n775), .Z(n777) );
  NAND2_X1 U872 ( .A1(n777), .A2(n776), .ZN(n786) );
  NOR2_X1 U873 ( .A1(G2090), .A2(G303), .ZN(n778) );
  XOR2_X1 U874 ( .A(KEYINPUT105), .B(n778), .Z(n779) );
  NAND2_X1 U875 ( .A1(n779), .A2(G8), .ZN(n782) );
  INV_X1 U876 ( .A(n780), .ZN(n781) );
  NAND2_X1 U877 ( .A1(n782), .A2(n781), .ZN(n784) );
  NAND2_X1 U878 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U879 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U880 ( .A1(G95), .A2(n887), .ZN(n791) );
  NAND2_X1 U881 ( .A1(G131), .A2(n888), .ZN(n790) );
  NAND2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U883 ( .A(KEYINPUT94), .B(n792), .Z(n796) );
  NAND2_X1 U884 ( .A1(n891), .A2(G107), .ZN(n794) );
  NAND2_X1 U885 ( .A1(G119), .A2(n892), .ZN(n793) );
  AND2_X1 U886 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n874) );
  NAND2_X1 U888 ( .A1(G1991), .A2(n874), .ZN(n805) );
  NAND2_X1 U889 ( .A1(G117), .A2(n891), .ZN(n798) );
  NAND2_X1 U890 ( .A1(G129), .A2(n892), .ZN(n797) );
  NAND2_X1 U891 ( .A1(n798), .A2(n797), .ZN(n801) );
  NAND2_X1 U892 ( .A1(n887), .A2(G105), .ZN(n799) );
  XOR2_X1 U893 ( .A(KEYINPUT38), .B(n799), .Z(n800) );
  NOR2_X1 U894 ( .A1(n801), .A2(n800), .ZN(n803) );
  NAND2_X1 U895 ( .A1(n888), .A2(G141), .ZN(n802) );
  NAND2_X1 U896 ( .A1(n803), .A2(n802), .ZN(n898) );
  NAND2_X1 U897 ( .A1(G1996), .A2(n898), .ZN(n804) );
  NAND2_X1 U898 ( .A1(n805), .A2(n804), .ZN(n921) );
  NOR2_X1 U899 ( .A1(n807), .A2(n806), .ZN(n835) );
  NAND2_X1 U900 ( .A1(n921), .A2(n835), .ZN(n808) );
  XNOR2_X1 U901 ( .A(n808), .B(KEYINPUT95), .ZN(n827) );
  NAND2_X1 U902 ( .A1(G104), .A2(n887), .ZN(n810) );
  NAND2_X1 U903 ( .A1(G140), .A2(n888), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U905 ( .A(KEYINPUT34), .B(n811), .ZN(n816) );
  NAND2_X1 U906 ( .A1(G116), .A2(n891), .ZN(n813) );
  NAND2_X1 U907 ( .A1(G128), .A2(n892), .ZN(n812) );
  NAND2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U909 ( .A(KEYINPUT35), .B(n814), .Z(n815) );
  NOR2_X1 U910 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U911 ( .A(KEYINPUT36), .B(n817), .ZN(n905) );
  XNOR2_X1 U912 ( .A(G2067), .B(KEYINPUT37), .ZN(n832) );
  NOR2_X1 U913 ( .A1(n905), .A2(n832), .ZN(n937) );
  NAND2_X1 U914 ( .A1(n835), .A2(n937), .ZN(n830) );
  NOR2_X1 U915 ( .A1(n827), .A2(n818), .ZN(n819) );
  NAND2_X1 U916 ( .A1(n518), .A2(n819), .ZN(n820) );
  XNOR2_X1 U917 ( .A(n820), .B(KEYINPUT107), .ZN(n822) );
  XNOR2_X1 U918 ( .A(G1986), .B(G290), .ZN(n974) );
  NAND2_X1 U919 ( .A1(n835), .A2(n974), .ZN(n821) );
  NAND2_X1 U920 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U921 ( .A(n823), .B(KEYINPUT108), .ZN(n838) );
  NOR2_X1 U922 ( .A1(G1996), .A2(n898), .ZN(n926) );
  NOR2_X1 U923 ( .A1(G1991), .A2(n874), .ZN(n922) );
  NOR2_X1 U924 ( .A1(G1986), .A2(G290), .ZN(n824) );
  XOR2_X1 U925 ( .A(n824), .B(KEYINPUT109), .Z(n825) );
  NOR2_X1 U926 ( .A1(n922), .A2(n825), .ZN(n826) );
  NOR2_X1 U927 ( .A1(n827), .A2(n826), .ZN(n828) );
  NOR2_X1 U928 ( .A1(n926), .A2(n828), .ZN(n829) );
  XNOR2_X1 U929 ( .A(n829), .B(KEYINPUT39), .ZN(n831) );
  NAND2_X1 U930 ( .A1(n831), .A2(n830), .ZN(n833) );
  NAND2_X1 U931 ( .A1(n905), .A2(n832), .ZN(n938) );
  NAND2_X1 U932 ( .A1(n833), .A2(n938), .ZN(n834) );
  NAND2_X1 U933 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U934 ( .A(KEYINPUT110), .B(n836), .ZN(n837) );
  NAND2_X1 U935 ( .A1(n838), .A2(n837), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n839), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U937 ( .A1(G2106), .A2(n840), .ZN(G217) );
  AND2_X1 U938 ( .A1(G15), .A2(G2), .ZN(n841) );
  NAND2_X1 U939 ( .A1(G661), .A2(n841), .ZN(G259) );
  NAND2_X1 U940 ( .A1(G3), .A2(G1), .ZN(n842) );
  NAND2_X1 U941 ( .A1(n843), .A2(n842), .ZN(G188) );
  INV_X1 U943 ( .A(G96), .ZN(G221) );
  NOR2_X1 U944 ( .A1(n845), .A2(n844), .ZN(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U946 ( .A(G1956), .B(G2474), .ZN(n855) );
  XOR2_X1 U947 ( .A(G1976), .B(G1971), .Z(n847) );
  XNOR2_X1 U948 ( .A(G1966), .B(G1961), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U950 ( .A(G1981), .B(G1996), .Z(n849) );
  XNOR2_X1 U951 ( .A(G1986), .B(G1991), .ZN(n848) );
  XNOR2_X1 U952 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U953 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U954 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(G229) );
  XOR2_X1 U957 ( .A(G2100), .B(G2096), .Z(n857) );
  XNOR2_X1 U958 ( .A(KEYINPUT42), .B(G2678), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U960 ( .A(KEYINPUT43), .B(G2090), .Z(n859) );
  XNOR2_X1 U961 ( .A(G2067), .B(G2072), .ZN(n858) );
  XNOR2_X1 U962 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U963 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U964 ( .A(G2084), .B(G2078), .ZN(n862) );
  XNOR2_X1 U965 ( .A(n863), .B(n862), .ZN(G227) );
  NAND2_X1 U966 ( .A1(n892), .A2(G124), .ZN(n864) );
  XNOR2_X1 U967 ( .A(n864), .B(KEYINPUT44), .ZN(n866) );
  NAND2_X1 U968 ( .A1(G136), .A2(n888), .ZN(n865) );
  NAND2_X1 U969 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U970 ( .A(n867), .B(KEYINPUT113), .ZN(n869) );
  NAND2_X1 U971 ( .A1(G100), .A2(n887), .ZN(n868) );
  NAND2_X1 U972 ( .A1(n869), .A2(n868), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n891), .A2(G112), .ZN(n870) );
  XOR2_X1 U974 ( .A(KEYINPUT114), .B(n870), .Z(n871) );
  NOR2_X1 U975 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U976 ( .A(KEYINPUT115), .B(n873), .Z(G162) );
  XNOR2_X1 U977 ( .A(G160), .B(n874), .ZN(n904) );
  NAND2_X1 U978 ( .A1(G118), .A2(n891), .ZN(n876) );
  NAND2_X1 U979 ( .A1(G130), .A2(n892), .ZN(n875) );
  NAND2_X1 U980 ( .A1(n876), .A2(n875), .ZN(n882) );
  NAND2_X1 U981 ( .A1(G106), .A2(n887), .ZN(n878) );
  NAND2_X1 U982 ( .A1(G142), .A2(n888), .ZN(n877) );
  NAND2_X1 U983 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U984 ( .A(KEYINPUT45), .B(n879), .Z(n880) );
  XNOR2_X1 U985 ( .A(KEYINPUT116), .B(n880), .ZN(n881) );
  NOR2_X1 U986 ( .A1(n882), .A2(n881), .ZN(n886) );
  XOR2_X1 U987 ( .A(KEYINPUT48), .B(KEYINPUT117), .Z(n884) );
  XNOR2_X1 U988 ( .A(G164), .B(KEYINPUT46), .ZN(n883) );
  XNOR2_X1 U989 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U990 ( .A(n886), .B(n885), .ZN(n900) );
  NAND2_X1 U991 ( .A1(G103), .A2(n887), .ZN(n890) );
  NAND2_X1 U992 ( .A1(G139), .A2(n888), .ZN(n889) );
  NAND2_X1 U993 ( .A1(n890), .A2(n889), .ZN(n897) );
  NAND2_X1 U994 ( .A1(G115), .A2(n891), .ZN(n894) );
  NAND2_X1 U995 ( .A1(G127), .A2(n892), .ZN(n893) );
  NAND2_X1 U996 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U997 ( .A(KEYINPUT47), .B(n895), .Z(n896) );
  NOR2_X1 U998 ( .A1(n897), .A2(n896), .ZN(n931) );
  XNOR2_X1 U999 ( .A(n898), .B(n931), .ZN(n899) );
  XNOR2_X1 U1000 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(G162), .B(n901), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n902), .B(n923), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n906) );
  XOR2_X1 U1004 ( .A(n906), .B(n905), .Z(n907) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n907), .ZN(G395) );
  XNOR2_X1 U1006 ( .A(G286), .B(n908), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(G171), .B(n971), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n911), .B(n988), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n912), .ZN(G397) );
  NOR2_X1 U1011 ( .A1(G229), .A2(G227), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(n913), .B(KEYINPUT49), .ZN(n916) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(n914), .B(KEYINPUT119), .ZN(n915) );
  NOR2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(n919) );
  NOR2_X1 U1016 ( .A1(G401), .A2(n920), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(n917), .B(KEYINPUT118), .ZN(n918) );
  NAND2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(n920), .ZN(G319) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n924) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n930) );
  XOR2_X1 U1023 ( .A(G2090), .B(G162), .Z(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1025 ( .A(KEYINPUT120), .B(n927), .Z(n928) );
  XOR2_X1 U1026 ( .A(KEYINPUT51), .B(n928), .Z(n929) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n943) );
  XOR2_X1 U1028 ( .A(G2072), .B(n931), .Z(n933) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1031 ( .A(KEYINPUT50), .B(n934), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(G160), .B(G2084), .ZN(n935) );
  NAND2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n941) );
  INV_X1 U1034 ( .A(n937), .ZN(n939) );
  NAND2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(KEYINPUT52), .B(n944), .ZN(n945) );
  XNOR2_X1 U1039 ( .A(KEYINPUT121), .B(n945), .ZN(n946) );
  INV_X1 U1040 ( .A(KEYINPUT55), .ZN(n966) );
  NAND2_X1 U1041 ( .A1(n946), .A2(n966), .ZN(n947) );
  NAND2_X1 U1042 ( .A1(n947), .A2(G29), .ZN(n1027) );
  XOR2_X1 U1043 ( .A(KEYINPUT122), .B(G34), .Z(n949) );
  XNOR2_X1 U1044 ( .A(G2084), .B(KEYINPUT54), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(n949), .B(n948), .ZN(n964) );
  XNOR2_X1 U1046 ( .A(G2090), .B(G35), .ZN(n962) );
  XNOR2_X1 U1047 ( .A(G2067), .B(G26), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(G33), .B(G2072), .ZN(n950) );
  NOR2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n956) );
  XOR2_X1 U1050 ( .A(G1991), .B(G25), .Z(n952) );
  NAND2_X1 U1051 ( .A1(n952), .A2(G28), .ZN(n954) );
  XNOR2_X1 U1052 ( .A(G32), .B(G1996), .ZN(n953) );
  NOR2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n959) );
  XOR2_X1 U1055 ( .A(G27), .B(n957), .Z(n958) );
  NOR2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1057 ( .A(KEYINPUT53), .B(n960), .ZN(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(n966), .B(n965), .ZN(n968) );
  INV_X1 U1061 ( .A(G29), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(G11), .A2(n969), .ZN(n1025) );
  INV_X1 U1064 ( .A(G16), .ZN(n1021) );
  XNOR2_X1 U1065 ( .A(KEYINPUT56), .B(KEYINPUT123), .ZN(n970) );
  XNOR2_X1 U1066 ( .A(n1021), .B(n970), .ZN(n996) );
  XNOR2_X1 U1067 ( .A(G1348), .B(n971), .ZN(n977) );
  XNOR2_X1 U1068 ( .A(n972), .B(G1956), .ZN(n973) );
  XNOR2_X1 U1069 ( .A(n973), .B(KEYINPUT125), .ZN(n975) );
  NOR2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n979) );
  XOR2_X1 U1072 ( .A(G171), .B(G1961), .Z(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n987) );
  XOR2_X1 U1075 ( .A(G1966), .B(KEYINPUT124), .Z(n982) );
  XNOR2_X1 U1076 ( .A(G168), .B(n982), .ZN(n984) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(KEYINPUT57), .B(n985), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n994) );
  XNOR2_X1 U1080 ( .A(n988), .B(G1341), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(G1971), .A2(G303), .ZN(n989) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n1023) );
  XNOR2_X1 U1086 ( .A(G20), .B(n997), .ZN(n1001) );
  XNOR2_X1 U1087 ( .A(G1981), .B(G6), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(G19), .B(G1341), .ZN(n998) );
  NOR2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1004) );
  XOR2_X1 U1091 ( .A(KEYINPUT59), .B(G1348), .Z(n1002) );
  XNOR2_X1 U1092 ( .A(G4), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(KEYINPUT60), .B(n1005), .ZN(n1017) );
  XOR2_X1 U1095 ( .A(G1966), .B(G21), .Z(n1008) );
  XNOR2_X1 U1096 ( .A(n1006), .B(G5), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1015) );
  XNOR2_X1 U1098 ( .A(G1986), .B(G24), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(G1971), .B(G22), .ZN(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XOR2_X1 U1101 ( .A(G1976), .B(G23), .Z(n1011) );
  NAND2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(KEYINPUT58), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(n1018), .B(KEYINPUT126), .ZN(n1019) );
  XOR2_X1 U1107 ( .A(KEYINPUT61), .B(n1019), .Z(n1020) );
  NAND2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(n1028), .B(KEYINPUT62), .ZN(n1029) );
  XNOR2_X1 U1113 ( .A(KEYINPUT127), .B(n1029), .ZN(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

