

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738;

  INV_X1 U369 ( .A(n673), .ZN(n348) );
  XNOR2_X1 U370 ( .A(n547), .B(n503), .ZN(n673) );
  INV_X2 U371 ( .A(G953), .ZN(n724) );
  NOR2_X4 U372 ( .A1(n513), .A2(n524), .ZN(n642) );
  NOR2_X2 U373 ( .A1(n400), .A2(n398), .ZN(n399) );
  NOR2_X2 U374 ( .A1(n409), .A2(n408), .ZN(n407) );
  INV_X1 U375 ( .A(n642), .ZN(n639) );
  NOR2_X1 U376 ( .A1(n529), .A2(n583), .ZN(n376) );
  XNOR2_X1 U377 ( .A(n401), .B(n350), .ZN(n657) );
  XNOR2_X1 U378 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n428) );
  AND2_X1 U379 ( .A1(n370), .A2(n369), .ZN(n368) );
  XNOR2_X1 U380 ( .A(n507), .B(n506), .ZN(n735) );
  OR2_X1 U381 ( .A1(n519), .A2(n688), .ZN(n507) );
  NOR2_X1 U382 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U383 ( .A(n505), .B(n356), .ZN(n688) );
  XNOR2_X1 U384 ( .A(n376), .B(KEYINPUT28), .ZN(n458) );
  AND2_X1 U385 ( .A1(n657), .A2(n658), .ZN(n508) );
  AND2_X1 U386 ( .A1(n372), .A2(G221), .ZN(n433) );
  XNOR2_X1 U387 ( .A(n429), .B(n428), .ZN(n372) );
  XNOR2_X1 U388 ( .A(n464), .B(KEYINPUT4), .ZN(n489) );
  XOR2_X1 U389 ( .A(G116), .B(G107), .Z(n486) );
  AND2_X2 U390 ( .A1(n368), .A2(n365), .ZN(n353) );
  NOR2_X1 U391 ( .A1(n568), .A2(n357), .ZN(n380) );
  XNOR2_X1 U392 ( .A(n589), .B(KEYINPUT45), .ZN(n594) );
  NAND2_X1 U393 ( .A1(n379), .A2(n405), .ZN(n388) );
  AND2_X1 U394 ( .A1(n383), .A2(n382), .ZN(n386) );
  NOR2_X1 U395 ( .A1(G953), .A2(G237), .ZN(n475) );
  XNOR2_X1 U396 ( .A(G902), .B(KEYINPUT15), .ZN(n590) );
  XOR2_X1 U397 ( .A(G122), .B(G104), .Z(n485) );
  AND2_X1 U398 ( .A1(G224), .A2(n724), .ZN(n495) );
  NAND2_X1 U399 ( .A1(n712), .A2(n598), .ZN(n655) );
  NOR2_X1 U400 ( .A1(n738), .A2(n731), .ZN(n568) );
  NOR2_X1 U401 ( .A1(n736), .A2(KEYINPUT44), .ZN(n406) );
  NOR2_X1 U402 ( .A1(G902), .A2(G237), .ZN(n459) );
  XNOR2_X1 U403 ( .A(n404), .B(G146), .ZN(n490) );
  INV_X1 U404 ( .A(G125), .ZN(n404) );
  XOR2_X1 U405 ( .A(KEYINPUT11), .B(KEYINPUT98), .Z(n477) );
  XNOR2_X1 U406 ( .A(G143), .B(G113), .ZN(n473) );
  XOR2_X1 U407 ( .A(G140), .B(G131), .Z(n474) );
  INV_X1 U408 ( .A(KEYINPUT73), .ZN(n371) );
  NAND2_X1 U409 ( .A1(n650), .A2(n371), .ZN(n369) );
  XNOR2_X1 U410 ( .A(n481), .B(G475), .ZN(n482) );
  OR2_X2 U411 ( .A1(n704), .A2(G902), .ZN(n401) );
  XNOR2_X1 U412 ( .A(KEYINPUT1), .B(n528), .ZN(n663) );
  XNOR2_X1 U413 ( .A(n361), .B(n421), .ZN(n620) );
  XNOR2_X1 U414 ( .A(n454), .B(n351), .ZN(n361) );
  XNOR2_X1 U415 ( .A(G128), .B(KEYINPUT82), .ZN(n430) );
  XNOR2_X1 U416 ( .A(G119), .B(G110), .ZN(n436) );
  XNOR2_X1 U417 ( .A(n490), .B(n403), .ZN(n721) );
  INV_X1 U418 ( .A(KEYINPUT10), .ZN(n403) );
  XNOR2_X1 U419 ( .A(n467), .B(n466), .ZN(n468) );
  BUF_X1 U420 ( .A(n547), .Z(n360) );
  BUF_X1 U421 ( .A(n512), .Z(n524) );
  OR2_X1 U422 ( .A1(n565), .A2(n570), .ZN(n409) );
  XNOR2_X1 U423 ( .A(n390), .B(n487), .ZN(n710) );
  XNOR2_X1 U424 ( .A(n484), .B(n391), .ZN(n390) );
  XNOR2_X1 U425 ( .A(n488), .B(KEYINPUT71), .ZN(n391) );
  AND2_X2 U426 ( .A1(n599), .A2(n655), .ZN(n705) );
  OR2_X1 U427 ( .A1(n638), .A2(n354), .ZN(n374) );
  NAND2_X1 U428 ( .A1(KEYINPUT85), .A2(KEYINPUT44), .ZN(n387) );
  XNOR2_X1 U429 ( .A(n588), .B(KEYINPUT104), .ZN(n379) );
  XNOR2_X1 U430 ( .A(G116), .B(G146), .ZN(n418) );
  XNOR2_X1 U431 ( .A(n489), .B(n417), .ZN(n454) );
  XNOR2_X1 U432 ( .A(G134), .B(G131), .ZN(n417) );
  XNOR2_X1 U433 ( .A(n491), .B(n494), .ZN(n413) );
  XNOR2_X1 U434 ( .A(n492), .B(n494), .ZN(n414) );
  NAND2_X1 U435 ( .A1(G237), .A2(G234), .ZN(n441) );
  NOR2_X1 U436 ( .A1(n663), .A2(n664), .ZN(n580) );
  XNOR2_X1 U437 ( .A(n502), .B(n501), .ZN(n516) );
  NAND2_X1 U438 ( .A1(n378), .A2(n355), .ZN(n529) );
  INV_X1 U439 ( .A(n658), .ZN(n377) );
  XNOR2_X1 U440 ( .A(n396), .B(n395), .ZN(n528) );
  XNOR2_X1 U441 ( .A(n456), .B(G469), .ZN(n395) );
  OR2_X1 U442 ( .A1(n700), .A2(G902), .ZN(n396) );
  XOR2_X1 U443 ( .A(G110), .B(KEYINPUT16), .Z(n488) );
  XNOR2_X1 U444 ( .A(n349), .B(n420), .ZN(n484) );
  XNOR2_X1 U445 ( .A(n364), .B(n480), .ZN(n613) );
  XNOR2_X1 U446 ( .A(n479), .B(n352), .ZN(n364) );
  NOR2_X1 U447 ( .A1(n650), .A2(n371), .ZN(n366) );
  NOR2_X1 U448 ( .A1(n594), .A2(n590), .ZN(n358) );
  XNOR2_X1 U449 ( .A(G107), .B(G104), .ZN(n448) );
  NOR2_X1 U450 ( .A1(n504), .A2(n673), .ZN(n505) );
  NAND2_X1 U451 ( .A1(n676), .A2(n558), .ZN(n504) );
  XNOR2_X1 U452 ( .A(n517), .B(KEYINPUT19), .ZN(n556) );
  NAND2_X1 U453 ( .A1(n516), .A2(n676), .ZN(n517) );
  XNOR2_X1 U454 ( .A(n402), .B(n435), .ZN(n704) );
  XNOR2_X1 U455 ( .A(n721), .B(n427), .ZN(n435) );
  XNOR2_X1 U456 ( .A(KEYINPUT23), .B(KEYINPUT94), .ZN(n427) );
  XNOR2_X1 U457 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U458 ( .A(n606), .B(n607), .ZN(n608) );
  XNOR2_X1 U459 ( .A(n534), .B(KEYINPUT36), .ZN(n535) );
  XNOR2_X1 U460 ( .A(n394), .B(n392), .ZN(n736) );
  XNOR2_X1 U461 ( .A(n393), .B(KEYINPUT35), .ZN(n392) );
  INV_X1 U462 ( .A(KEYINPUT77), .ZN(n393) );
  XNOR2_X1 U463 ( .A(n407), .B(KEYINPUT32), .ZN(n738) );
  XNOR2_X1 U464 ( .A(n702), .B(n701), .ZN(n703) );
  XOR2_X1 U465 ( .A(G101), .B(KEYINPUT3), .Z(n349) );
  XNOR2_X1 U466 ( .A(n440), .B(n439), .ZN(n350) );
  XOR2_X1 U467 ( .A(n419), .B(n418), .Z(n351) );
  XOR2_X1 U468 ( .A(n474), .B(n473), .Z(n352) );
  BUF_X1 U469 ( .A(n657), .Z(n363) );
  OR2_X1 U470 ( .A1(n678), .A2(n375), .ZN(n354) );
  NOR2_X1 U471 ( .A1(n510), .A2(n377), .ZN(n355) );
  XNOR2_X1 U472 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n356) );
  INV_X1 U473 ( .A(KEYINPUT85), .ZN(n389) );
  AND2_X1 U474 ( .A1(n389), .A2(KEYINPUT44), .ZN(n357) );
  NAND2_X1 U475 ( .A1(n353), .A2(n358), .ZN(n593) );
  INV_X1 U476 ( .A(n516), .ZN(n547) );
  XNOR2_X2 U477 ( .A(n359), .B(KEYINPUT0), .ZN(n569) );
  NAND2_X1 U478 ( .A1(n556), .A2(n557), .ZN(n359) );
  NOR2_X2 U479 ( .A1(n386), .A2(n388), .ZN(n589) );
  XNOR2_X1 U480 ( .A(n455), .B(n720), .ZN(n700) );
  NAND2_X1 U481 ( .A1(n576), .A2(n575), .ZN(n394) );
  XNOR2_X1 U482 ( .A(n497), .B(n710), .ZN(n606) );
  XNOR2_X1 U483 ( .A(n362), .B(KEYINPUT30), .ZN(n509) );
  NAND2_X1 U484 ( .A1(n661), .A2(n676), .ZN(n362) );
  NAND2_X1 U485 ( .A1(n733), .A2(n735), .ZN(n515) );
  XNOR2_X2 U486 ( .A(n514), .B(KEYINPUT40), .ZN(n733) );
  NOR2_X2 U487 ( .A1(n509), .A2(n510), .ZN(n511) );
  XNOR2_X1 U488 ( .A(n536), .B(n535), .ZN(n537) );
  NOR2_X1 U489 ( .A1(n597), .A2(n650), .ZN(n722) );
  NAND2_X1 U490 ( .A1(n367), .A2(n366), .ZN(n365) );
  INV_X1 U491 ( .A(n597), .ZN(n367) );
  NAND2_X1 U492 ( .A1(n597), .A2(n371), .ZN(n370) );
  NAND2_X1 U493 ( .A1(n372), .A2(G217), .ZN(n462) );
  XNOR2_X1 U494 ( .A(n374), .B(n373), .ZN(n527) );
  INV_X1 U495 ( .A(KEYINPUT47), .ZN(n373) );
  INV_X1 U496 ( .A(KEYINPUT66), .ZN(n375) );
  INV_X1 U497 ( .A(n657), .ZN(n378) );
  NAND2_X1 U498 ( .A1(n381), .A2(n380), .ZN(n382) );
  NAND2_X1 U499 ( .A1(n406), .A2(KEYINPUT85), .ZN(n381) );
  NAND2_X1 U500 ( .A1(n384), .A2(n385), .ZN(n383) );
  AND2_X1 U501 ( .A1(n568), .A2(n387), .ZN(n384) );
  NAND2_X1 U502 ( .A1(n406), .A2(n389), .ZN(n385) );
  XNOR2_X1 U503 ( .A(n483), .B(n482), .ZN(n512) );
  XNOR2_X1 U504 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U505 ( .A(n434), .B(n437), .ZN(n402) );
  INV_X1 U506 ( .A(n400), .ZN(n584) );
  OR2_X1 U507 ( .A1(n400), .A2(n397), .ZN(n522) );
  INV_X1 U508 ( .A(n511), .ZN(n397) );
  NAND2_X1 U509 ( .A1(n348), .A2(n511), .ZN(n398) );
  XNOR2_X1 U510 ( .A(n399), .B(KEYINPUT39), .ZN(n550) );
  OR2_X2 U511 ( .A1(n664), .A2(n528), .ZN(n400) );
  NAND2_X1 U512 ( .A1(n736), .A2(KEYINPUT44), .ZN(n405) );
  INV_X1 U513 ( .A(n409), .ZN(n577) );
  NAND2_X1 U514 ( .A1(n567), .A2(n378), .ZN(n408) );
  NAND2_X1 U515 ( .A1(n411), .A2(n410), .ZN(n496) );
  NAND2_X1 U516 ( .A1(n493), .A2(n414), .ZN(n410) );
  NAND2_X1 U517 ( .A1(n412), .A2(n413), .ZN(n411) );
  INV_X1 U518 ( .A(n493), .ZN(n412) );
  AND2_X1 U519 ( .A1(G210), .A2(n475), .ZN(n415) );
  XNOR2_X1 U520 ( .A(KEYINPUT103), .B(n559), .ZN(n416) );
  INV_X1 U521 ( .A(n648), .ZN(n538) );
  NAND2_X1 U522 ( .A1(n539), .A2(n538), .ZN(n540) );
  INV_X1 U523 ( .A(n464), .ZN(n465) );
  INV_X1 U524 ( .A(KEYINPUT102), .ZN(n466) );
  INV_X1 U525 ( .A(KEYINPUT90), .ZN(n499) );
  INV_X1 U526 ( .A(KEYINPUT86), .ZN(n534) );
  XNOR2_X1 U527 ( .A(n500), .B(n499), .ZN(n501) );
  INV_X1 U528 ( .A(n600), .ZN(n601) );
  XNOR2_X1 U529 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U530 ( .A(n617), .B(KEYINPUT64), .ZN(n618) );
  XNOR2_X2 U531 ( .A(G143), .B(G128), .ZN(n464) );
  XOR2_X1 U532 ( .A(G137), .B(KEYINPUT5), .Z(n419) );
  XNOR2_X1 U533 ( .A(G113), .B(G119), .ZN(n420) );
  XNOR2_X1 U534 ( .A(n484), .B(n415), .ZN(n421) );
  NOR2_X1 U535 ( .A1(n620), .A2(G902), .ZN(n422) );
  XNOR2_X2 U536 ( .A(n422), .B(G472), .ZN(n583) );
  XOR2_X1 U537 ( .A(KEYINPUT96), .B(KEYINPUT21), .Z(n426) );
  XOR2_X1 U538 ( .A(KEYINPUT95), .B(KEYINPUT20), .Z(n424) );
  NAND2_X1 U539 ( .A1(G234), .A2(n590), .ZN(n423) );
  XNOR2_X1 U540 ( .A(n424), .B(n423), .ZN(n438) );
  NAND2_X1 U541 ( .A1(G221), .A2(n438), .ZN(n425) );
  XNOR2_X1 U542 ( .A(n426), .B(n425), .ZN(n658) );
  NAND2_X1 U543 ( .A1(n724), .A2(G234), .ZN(n429) );
  XOR2_X1 U544 ( .A(KEYINPUT75), .B(KEYINPUT24), .Z(n431) );
  XNOR2_X1 U545 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U546 ( .A(G140), .B(G137), .Z(n453) );
  XNOR2_X1 U547 ( .A(n436), .B(n453), .ZN(n437) );
  XOR2_X1 U548 ( .A(KEYINPUT25), .B(KEYINPUT74), .Z(n440) );
  NAND2_X1 U549 ( .A1(n438), .A2(G217), .ZN(n439) );
  XNOR2_X1 U550 ( .A(n441), .B(KEYINPUT14), .ZN(n443) );
  NAND2_X1 U551 ( .A1(G952), .A2(n443), .ZN(n442) );
  XOR2_X1 U552 ( .A(KEYINPUT91), .B(n442), .Z(n687) );
  NOR2_X1 U553 ( .A1(G953), .A2(n687), .ZN(n554) );
  INV_X1 U554 ( .A(n554), .ZN(n446) );
  NAND2_X1 U555 ( .A1(G902), .A2(n443), .ZN(n552) );
  NOR2_X1 U556 ( .A1(G900), .A2(n552), .ZN(n444) );
  NAND2_X1 U557 ( .A1(G953), .A2(n444), .ZN(n445) );
  NAND2_X1 U558 ( .A1(n446), .A2(n445), .ZN(n447) );
  XOR2_X1 U559 ( .A(KEYINPUT80), .B(n447), .Z(n510) );
  XOR2_X1 U560 ( .A(G110), .B(G101), .Z(n449) );
  XNOR2_X1 U561 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U562 ( .A(G146), .B(n450), .Z(n452) );
  NAND2_X1 U563 ( .A1(G227), .A2(n724), .ZN(n451) );
  XNOR2_X1 U564 ( .A(n452), .B(n451), .ZN(n455) );
  XNOR2_X1 U565 ( .A(n454), .B(n453), .ZN(n720) );
  XNOR2_X1 U566 ( .A(KEYINPUT68), .B(KEYINPUT69), .ZN(n456) );
  XNOR2_X1 U567 ( .A(n528), .B(KEYINPUT109), .ZN(n457) );
  NAND2_X1 U568 ( .A1(n458), .A2(n457), .ZN(n519) );
  XOR2_X1 U569 ( .A(KEYINPUT72), .B(n459), .Z(n498) );
  NAND2_X1 U570 ( .A1(G214), .A2(n498), .ZN(n676) );
  XOR2_X1 U571 ( .A(KEYINPUT100), .B(KEYINPUT9), .Z(n461) );
  XNOR2_X1 U572 ( .A(KEYINPUT101), .B(KEYINPUT7), .ZN(n460) );
  XNOR2_X1 U573 ( .A(n461), .B(n460), .ZN(n471) );
  XOR2_X1 U574 ( .A(n486), .B(G134), .Z(n463) );
  XNOR2_X1 U575 ( .A(n463), .B(n462), .ZN(n469) );
  XNOR2_X1 U576 ( .A(n465), .B(G122), .ZN(n467) );
  XNOR2_X1 U577 ( .A(n471), .B(n470), .ZN(n600) );
  NOR2_X1 U578 ( .A1(n600), .A2(G902), .ZN(n472) );
  XNOR2_X1 U579 ( .A(n472), .B(G478), .ZN(n525) );
  INV_X1 U580 ( .A(n525), .ZN(n513) );
  NAND2_X1 U581 ( .A1(n475), .A2(G214), .ZN(n476) );
  XNOR2_X1 U582 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U583 ( .A(n478), .B(KEYINPUT12), .Z(n480) );
  XNOR2_X1 U584 ( .A(n721), .B(n485), .ZN(n479) );
  NOR2_X1 U585 ( .A1(G902), .A2(n613), .ZN(n483) );
  XNOR2_X1 U586 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n481) );
  INV_X1 U587 ( .A(n512), .ZN(n521) );
  NOR2_X2 U588 ( .A1(n513), .A2(n521), .ZN(n558) );
  INV_X1 U589 ( .A(n558), .ZN(n675) );
  XNOR2_X1 U590 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U591 ( .A(n489), .B(n490), .ZN(n493) );
  XOR2_X1 U592 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n492) );
  INV_X1 U593 ( .A(n492), .ZN(n491) );
  INV_X1 U594 ( .A(KEYINPUT76), .ZN(n494) );
  XNOR2_X1 U595 ( .A(n496), .B(n495), .ZN(n497) );
  NAND2_X1 U596 ( .A1(n606), .A2(n590), .ZN(n502) );
  NAND2_X1 U597 ( .A1(G210), .A2(n498), .ZN(n500) );
  INV_X1 U598 ( .A(KEYINPUT38), .ZN(n503) );
  XOR2_X1 U599 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n506) );
  XNOR2_X1 U600 ( .A(n508), .B(KEYINPUT65), .ZN(n664) );
  INV_X2 U601 ( .A(n583), .ZN(n661) );
  OR2_X2 U602 ( .A1(n550), .A2(n639), .ZN(n514) );
  XNOR2_X1 U603 ( .A(n515), .B(KEYINPUT46), .ZN(n541) );
  INV_X1 U604 ( .A(n556), .ZN(n518) );
  XNOR2_X1 U605 ( .A(n520), .B(KEYINPUT79), .ZN(n638) );
  NOR2_X1 U606 ( .A1(n521), .A2(n525), .ZN(n645) );
  NOR2_X1 U607 ( .A1(n642), .A2(n645), .ZN(n678) );
  NOR2_X1 U608 ( .A1(n360), .A2(n522), .ZN(n523) );
  XNOR2_X1 U609 ( .A(KEYINPUT108), .B(n523), .ZN(n526) );
  NOR2_X1 U610 ( .A1(n525), .A2(n524), .ZN(n575) );
  NAND2_X1 U611 ( .A1(n526), .A2(n575), .ZN(n637) );
  AND2_X1 U612 ( .A1(n527), .A2(n637), .ZN(n539) );
  XOR2_X1 U613 ( .A(KEYINPUT87), .B(n663), .Z(n566) );
  XNOR2_X1 U614 ( .A(KEYINPUT6), .B(n583), .ZN(n570) );
  INV_X1 U615 ( .A(n529), .ZN(n530) );
  NAND2_X1 U616 ( .A1(n570), .A2(n530), .ZN(n531) );
  NOR2_X1 U617 ( .A1(n639), .A2(n531), .ZN(n532) );
  XNOR2_X1 U618 ( .A(n532), .B(KEYINPUT106), .ZN(n533) );
  NAND2_X1 U619 ( .A1(n533), .A2(n676), .ZN(n543) );
  NOR2_X1 U620 ( .A1(n543), .A2(n360), .ZN(n536) );
  NOR2_X1 U621 ( .A1(n566), .A2(n537), .ZN(n648) );
  NOR2_X2 U622 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U623 ( .A(n542), .B(KEYINPUT48), .ZN(n548) );
  INV_X1 U624 ( .A(n663), .ZN(n579) );
  NOR2_X1 U625 ( .A1(n579), .A2(n543), .ZN(n545) );
  XNOR2_X1 U626 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n544) );
  XNOR2_X1 U627 ( .A(n545), .B(n544), .ZN(n546) );
  NAND2_X1 U628 ( .A1(n360), .A2(n546), .ZN(n652) );
  NAND2_X1 U629 ( .A1(n548), .A2(n652), .ZN(n549) );
  XNOR2_X2 U630 ( .A(n549), .B(KEYINPUT84), .ZN(n597) );
  INV_X1 U631 ( .A(n645), .ZN(n633) );
  NOR2_X1 U632 ( .A1(n633), .A2(n550), .ZN(n650) );
  NOR2_X1 U633 ( .A1(G898), .A2(n724), .ZN(n551) );
  XOR2_X1 U634 ( .A(KEYINPUT92), .B(n551), .Z(n711) );
  NOR2_X1 U635 ( .A1(n711), .A2(n552), .ZN(n553) );
  NOR2_X1 U636 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U637 ( .A(KEYINPUT93), .B(n555), .ZN(n557) );
  INV_X1 U638 ( .A(n569), .ZN(n560) );
  NAND2_X1 U639 ( .A1(n658), .A2(n558), .ZN(n559) );
  NAND2_X1 U640 ( .A1(n560), .A2(n416), .ZN(n561) );
  XNOR2_X1 U641 ( .A(n561), .B(KEYINPUT22), .ZN(n565) );
  NOR2_X1 U642 ( .A1(n363), .A2(n565), .ZN(n563) );
  NOR2_X1 U643 ( .A1(n661), .A2(n579), .ZN(n562) );
  NAND2_X1 U644 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U645 ( .A(KEYINPUT105), .B(n564), .ZN(n731) );
  INV_X1 U646 ( .A(n566), .ZN(n567) );
  XNOR2_X1 U647 ( .A(KEYINPUT34), .B(KEYINPUT78), .ZN(n574) );
  XOR2_X1 U648 ( .A(KEYINPUT33), .B(KEYINPUT70), .Z(n572) );
  NAND2_X1 U649 ( .A1(n570), .A2(n580), .ZN(n571) );
  XNOR2_X1 U650 ( .A(n572), .B(n571), .ZN(n689) );
  NOR2_X1 U651 ( .A1(n569), .A2(n689), .ZN(n573) );
  XNOR2_X1 U652 ( .A(n574), .B(n573), .ZN(n576) );
  NAND2_X1 U653 ( .A1(n363), .A2(n577), .ZN(n578) );
  NOR2_X1 U654 ( .A1(n579), .A2(n578), .ZN(n627) );
  NAND2_X1 U655 ( .A1(n661), .A2(n580), .ZN(n669) );
  NOR2_X1 U656 ( .A1(n569), .A2(n669), .ZN(n581) );
  XNOR2_X1 U657 ( .A(n581), .B(KEYINPUT97), .ZN(n582) );
  XNOR2_X1 U658 ( .A(n582), .B(KEYINPUT31), .ZN(n646) );
  NAND2_X1 U659 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U660 ( .A1(n569), .A2(n585), .ZN(n629) );
  NOR2_X1 U661 ( .A1(n646), .A2(n629), .ZN(n586) );
  NOR2_X1 U662 ( .A1(n678), .A2(n586), .ZN(n587) );
  NOR2_X1 U663 ( .A1(n627), .A2(n587), .ZN(n588) );
  XNOR2_X1 U664 ( .A(n590), .B(KEYINPUT83), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n591), .A2(KEYINPUT2), .ZN(n592) );
  NAND2_X1 U666 ( .A1(n593), .A2(n592), .ZN(n599) );
  INV_X1 U667 ( .A(n594), .ZN(n712) );
  INV_X1 U668 ( .A(KEYINPUT2), .ZN(n653) );
  OR2_X1 U669 ( .A1(n653), .A2(n650), .ZN(n595) );
  XOR2_X1 U670 ( .A(KEYINPUT81), .B(n595), .Z(n596) );
  NOR2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U672 ( .A1(n705), .A2(G478), .ZN(n602) );
  XNOR2_X1 U673 ( .A(n602), .B(n601), .ZN(n604) );
  NOR2_X1 U674 ( .A1(G952), .A2(n724), .ZN(n603) );
  XNOR2_X1 U675 ( .A(KEYINPUT89), .B(n603), .ZN(n698) );
  NAND2_X1 U676 ( .A1(n604), .A2(n698), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n605), .B(KEYINPUT123), .ZN(G63) );
  NAND2_X1 U678 ( .A1(n705), .A2(G210), .ZN(n609) );
  XOR2_X1 U679 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n607) );
  XNOR2_X1 U680 ( .A(n609), .B(n608), .ZN(n610) );
  NAND2_X1 U681 ( .A1(n610), .A2(n698), .ZN(n612) );
  INV_X1 U682 ( .A(KEYINPUT56), .ZN(n611) );
  XNOR2_X1 U683 ( .A(n612), .B(n611), .ZN(G51) );
  NAND2_X1 U684 ( .A1(n705), .A2(G475), .ZN(n615) );
  XNOR2_X1 U685 ( .A(n613), .B(KEYINPUT59), .ZN(n614) );
  XNOR2_X1 U686 ( .A(n615), .B(n614), .ZN(n616) );
  NAND2_X1 U687 ( .A1(n616), .A2(n698), .ZN(n619) );
  INV_X1 U688 ( .A(KEYINPUT60), .ZN(n617) );
  XNOR2_X1 U689 ( .A(n619), .B(n618), .ZN(G60) );
  NAND2_X1 U690 ( .A1(n705), .A2(G472), .ZN(n622) );
  XOR2_X1 U691 ( .A(n620), .B(KEYINPUT62), .Z(n621) );
  XNOR2_X1 U692 ( .A(n622), .B(n621), .ZN(n623) );
  NAND2_X1 U693 ( .A1(n623), .A2(n698), .ZN(n626) );
  XNOR2_X1 U694 ( .A(KEYINPUT88), .B(KEYINPUT112), .ZN(n624) );
  XNOR2_X1 U695 ( .A(n624), .B(KEYINPUT63), .ZN(n625) );
  XNOR2_X1 U696 ( .A(n626), .B(n625), .ZN(G57) );
  XOR2_X1 U697 ( .A(G101), .B(n627), .Z(G3) );
  NAND2_X1 U698 ( .A1(n629), .A2(n642), .ZN(n628) );
  XNOR2_X1 U699 ( .A(n628), .B(G104), .ZN(G6) );
  XOR2_X1 U700 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n631) );
  NAND2_X1 U701 ( .A1(n629), .A2(n645), .ZN(n630) );
  XNOR2_X1 U702 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U703 ( .A(G107), .B(n632), .ZN(G9) );
  NOR2_X1 U704 ( .A1(n633), .A2(n638), .ZN(n635) );
  XNOR2_X1 U705 ( .A(KEYINPUT114), .B(KEYINPUT29), .ZN(n634) );
  XNOR2_X1 U706 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U707 ( .A(G128), .B(n636), .ZN(G30) );
  XNOR2_X1 U708 ( .A(G143), .B(n637), .ZN(G45) );
  NOR2_X1 U709 ( .A1(n639), .A2(n638), .ZN(n641) );
  XNOR2_X1 U710 ( .A(G146), .B(KEYINPUT115), .ZN(n640) );
  XNOR2_X1 U711 ( .A(n641), .B(n640), .ZN(G48) );
  NAND2_X1 U712 ( .A1(n646), .A2(n642), .ZN(n643) );
  XNOR2_X1 U713 ( .A(n643), .B(KEYINPUT116), .ZN(n644) );
  XNOR2_X1 U714 ( .A(G113), .B(n644), .ZN(G15) );
  NAND2_X1 U715 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U716 ( .A(n647), .B(G116), .ZN(G18) );
  XNOR2_X1 U717 ( .A(G125), .B(n648), .ZN(n649) );
  XNOR2_X1 U718 ( .A(n649), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U719 ( .A(G134), .B(n650), .Z(G36) );
  XOR2_X1 U720 ( .A(G140), .B(KEYINPUT117), .Z(n651) );
  XNOR2_X1 U721 ( .A(n652), .B(n651), .ZN(G42) );
  NAND2_X1 U722 ( .A1(n722), .A2(n712), .ZN(n654) );
  NAND2_X1 U723 ( .A1(n654), .A2(n653), .ZN(n656) );
  NAND2_X1 U724 ( .A1(n656), .A2(n655), .ZN(n695) );
  NOR2_X1 U725 ( .A1(n658), .A2(n363), .ZN(n659) );
  XOR2_X1 U726 ( .A(KEYINPUT49), .B(n659), .Z(n660) );
  NOR2_X1 U727 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U728 ( .A(n662), .B(KEYINPUT118), .ZN(n668) );
  XOR2_X1 U729 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n666) );
  NAND2_X1 U730 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U731 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U732 ( .A1(n668), .A2(n667), .ZN(n670) );
  NAND2_X1 U733 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U734 ( .A(KEYINPUT51), .B(n671), .ZN(n672) );
  NOR2_X1 U735 ( .A1(n688), .A2(n672), .ZN(n684) );
  NOR2_X1 U736 ( .A1(n676), .A2(n348), .ZN(n674) );
  NOR2_X1 U737 ( .A1(n675), .A2(n674), .ZN(n681) );
  NAND2_X1 U738 ( .A1(n676), .A2(n348), .ZN(n677) );
  NOR2_X1 U739 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U740 ( .A(n679), .B(KEYINPUT120), .ZN(n680) );
  NOR2_X1 U741 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U742 ( .A1(n689), .A2(n682), .ZN(n683) );
  NOR2_X1 U743 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U744 ( .A(n685), .B(KEYINPUT52), .ZN(n686) );
  NOR2_X1 U745 ( .A1(n687), .A2(n686), .ZN(n691) );
  NOR2_X1 U746 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U747 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U748 ( .A(n692), .B(KEYINPUT121), .ZN(n693) );
  NOR2_X1 U749 ( .A1(G953), .A2(n693), .ZN(n694) );
  NAND2_X1 U750 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U751 ( .A(KEYINPUT122), .B(n696), .Z(n697) );
  XNOR2_X1 U752 ( .A(KEYINPUT53), .B(n697), .ZN(G75) );
  INV_X1 U753 ( .A(n698), .ZN(n709) );
  NAND2_X1 U754 ( .A1(n705), .A2(G469), .ZN(n702) );
  XOR2_X1 U755 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n699) );
  NOR2_X1 U756 ( .A1(n709), .A2(n703), .ZN(G54) );
  XNOR2_X1 U757 ( .A(n704), .B(KEYINPUT124), .ZN(n707) );
  NAND2_X1 U758 ( .A1(G217), .A2(n705), .ZN(n706) );
  XNOR2_X1 U759 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U760 ( .A1(n709), .A2(n708), .ZN(G66) );
  NAND2_X1 U761 ( .A1(n711), .A2(n710), .ZN(n719) );
  NAND2_X1 U762 ( .A1(n724), .A2(n712), .ZN(n716) );
  NAND2_X1 U763 ( .A1(G953), .A2(G224), .ZN(n713) );
  XNOR2_X1 U764 ( .A(KEYINPUT61), .B(n713), .ZN(n714) );
  NAND2_X1 U765 ( .A1(n714), .A2(G898), .ZN(n715) );
  NAND2_X1 U766 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U767 ( .A(n717), .B(KEYINPUT125), .ZN(n718) );
  XNOR2_X1 U768 ( .A(n719), .B(n718), .ZN(G69) );
  XNOR2_X1 U769 ( .A(n721), .B(n720), .ZN(n726) );
  INV_X1 U770 ( .A(n726), .ZN(n723) );
  XNOR2_X1 U771 ( .A(n723), .B(n722), .ZN(n725) );
  NAND2_X1 U772 ( .A1(n725), .A2(n724), .ZN(n730) );
  XNOR2_X1 U773 ( .A(G227), .B(n726), .ZN(n727) );
  NAND2_X1 U774 ( .A1(n727), .A2(G900), .ZN(n728) );
  NAND2_X1 U775 ( .A1(n728), .A2(G953), .ZN(n729) );
  NAND2_X1 U776 ( .A1(n730), .A2(n729), .ZN(G72) );
  XNOR2_X1 U777 ( .A(G110), .B(n731), .ZN(n732) );
  XNOR2_X1 U778 ( .A(n732), .B(KEYINPUT113), .ZN(G12) );
  XOR2_X1 U779 ( .A(n733), .B(G131), .Z(n734) );
  XNOR2_X1 U780 ( .A(KEYINPUT127), .B(n734), .ZN(G33) );
  XNOR2_X1 U781 ( .A(G137), .B(n735), .ZN(G39) );
  XOR2_X1 U782 ( .A(G122), .B(n736), .Z(n737) );
  XNOR2_X1 U783 ( .A(KEYINPUT126), .B(n737), .ZN(G24) );
  XOR2_X1 U784 ( .A(G119), .B(n738), .Z(G21) );
endmodule

