//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 0 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1254, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1341,
    new_n1342;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR3_X1   g0001(.A1(new_n201), .A2(G58), .A3(G68), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  AND2_X1   g0003(.A1(new_n202), .A2(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(KEYINPUT65), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT65), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G20), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  AND2_X1   g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n214), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n206), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n209), .B(new_n218), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT66), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NOR2_X1   g0046(.A1(G20), .A2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G150), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT65), .B(G20), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G33), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT8), .B(G58), .ZN(new_n251));
  OAI221_X1 g0051(.A(new_n248), .B1(new_n250), .B2(new_n251), .C1(new_n202), .C2(new_n210), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G1), .A2(G13), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G13), .ZN(new_n257));
  NOR3_X1   g0057(.A1(new_n257), .A2(new_n210), .A3(G1), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n255), .ZN(new_n259));
  INV_X1    g0059(.A(G50), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n260), .B1(new_n261), .B2(G20), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n259), .A2(new_n262), .B1(new_n260), .B2(new_n258), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n256), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  OR2_X1    g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1698), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G222), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G223), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(G1698), .ZN(new_n272));
  OAI221_X1 g0072(.A(new_n269), .B1(new_n203), .B2(new_n270), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G1), .A3(G13), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G45), .ZN(new_n279));
  AOI21_X1  g0079(.A(G1), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(new_n275), .A3(G274), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n278), .A2(new_n279), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n261), .A2(new_n283), .B1(new_n215), .B2(new_n274), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n282), .B1(G226), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n277), .A2(new_n285), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n265), .A2(KEYINPUT9), .B1(G200), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n286), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT9), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n288), .A2(G190), .B1(new_n264), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n291), .B(KEYINPUT10), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n286), .A2(G179), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n294), .B(new_n264), .C1(G169), .C2(new_n288), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n251), .B1(new_n261), .B2(G20), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n297), .A2(new_n259), .B1(new_n258), .B2(new_n251), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT7), .B1(new_n214), .B2(new_n270), .ZN(new_n300));
  AND2_X1   g0100(.A1(KEYINPUT3), .A2(G33), .ZN(new_n301));
  NOR2_X1   g0101(.A1(KEYINPUT3), .A2(G33), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT7), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n303), .A2(new_n304), .A3(new_n210), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n300), .A2(G68), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(KEYINPUT72), .B1(new_n247), .B2(G159), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n247), .A2(KEYINPUT72), .A3(G159), .ZN(new_n309));
  XNOR2_X1  g0109(.A(G58), .B(G68), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n308), .A2(new_n309), .B1(G20), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT16), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n255), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n310), .A2(G20), .ZN(new_n316));
  INV_X1    g0116(.A(new_n309), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n316), .B(KEYINPUT16), .C1(new_n317), .C2(new_n307), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT7), .B1(new_n270), .B2(G20), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n303), .A2(new_n249), .A3(new_n304), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(new_n321), .A3(G68), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n315), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n299), .B1(new_n314), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G1698), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n271), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G226), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G1698), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n326), .B(new_n328), .C1(new_n301), .C2(new_n302), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G33), .A2(G87), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n275), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n275), .A2(G232), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n281), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(G169), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n329), .A2(new_n330), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n276), .ZN(new_n337));
  INV_X1    g0137(.A(G274), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n338), .B1(new_n215), .B2(new_n274), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n284), .A2(G232), .B1(new_n339), .B2(new_n280), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G179), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n335), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n324), .A2(new_n344), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n345), .A2(KEYINPUT73), .A3(KEYINPUT18), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n314), .A2(new_n323), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n298), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT18), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n349), .A3(new_n343), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT18), .B1(new_n324), .B2(new_n344), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n346), .B1(KEYINPUT73), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G190), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n337), .A2(new_n354), .A3(new_n340), .ZN(new_n355));
  INV_X1    g0155(.A(G200), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n331), .B2(new_n334), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT17), .B1(new_n324), .B2(new_n358), .ZN(new_n359));
  AND3_X1   g0159(.A1(new_n320), .A2(new_n321), .A3(G68), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n255), .B1(new_n360), .B2(new_n318), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT16), .B1(new_n306), .B2(new_n311), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n358), .B(new_n298), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT74), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n347), .A2(KEYINPUT74), .A3(new_n298), .A4(new_n358), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n359), .B1(new_n367), .B2(KEYINPUT17), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n353), .A2(new_n368), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n247), .A2(G50), .B1(G20), .B2(new_n220), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n250), .B2(new_n203), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n255), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT11), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n371), .A2(KEYINPUT11), .A3(new_n255), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n257), .A2(G1), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G20), .ZN(new_n377));
  OR3_X1    g0177(.A1(new_n377), .A2(KEYINPUT12), .A3(G68), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT12), .B1(new_n377), .B2(G68), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n220), .B1(new_n261), .B2(G20), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n378), .A2(new_n379), .B1(new_n259), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n374), .A2(new_n375), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n327), .A2(new_n325), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n270), .B(new_n383), .C1(G232), .C2(new_n325), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G33), .A2(G97), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n275), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  XOR2_X1   g0186(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n284), .A2(G238), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n281), .ZN(new_n390));
  OR3_X1    g0190(.A1(new_n386), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n388), .B1(new_n386), .B2(new_n390), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n382), .B1(new_n393), .B2(G200), .ZN(new_n394));
  OR3_X1    g0194(.A1(new_n386), .A2(new_n390), .A3(KEYINPUT70), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT70), .B1(new_n386), .B2(new_n390), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(KEYINPUT13), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(G190), .A3(new_n391), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT71), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n394), .A2(new_n398), .A3(KEYINPUT71), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n393), .A2(G169), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT14), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n397), .A2(G179), .A3(new_n391), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT14), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n393), .A2(new_n407), .A3(G169), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n382), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n403), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n268), .A2(G232), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n412), .B(KEYINPUT67), .ZN(new_n413));
  INV_X1    g0213(.A(G107), .ZN(new_n414));
  OAI22_X1  g0214(.A1(new_n272), .A2(new_n221), .B1(new_n414), .B2(new_n270), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n416), .A2(new_n275), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n282), .B1(G244), .B2(new_n284), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n342), .ZN(new_n421));
  XNOR2_X1  g0221(.A(KEYINPUT15), .B(G87), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT68), .B1(new_n250), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n251), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n424), .A2(new_n247), .B1(new_n214), .B2(G77), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NOR3_X1   g0226(.A1(new_n250), .A2(KEYINPUT68), .A3(new_n422), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n255), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n203), .B1(new_n261), .B2(G20), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n259), .A2(new_n429), .B1(new_n203), .B2(new_n258), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n421), .B(new_n431), .C1(G169), .C2(new_n420), .ZN(new_n432));
  INV_X1    g0232(.A(new_n431), .ZN(new_n433));
  OAI211_X1 g0233(.A(G190), .B(new_n418), .C1(new_n416), .C2(new_n275), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n433), .B(new_n434), .C1(new_n420), .C2(new_n356), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  NOR4_X1   g0236(.A1(new_n296), .A2(new_n369), .A3(new_n411), .A4(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G116), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n258), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n261), .A2(G33), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n315), .A2(new_n377), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G116), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n253), .A2(new_n254), .B1(G20), .B2(new_n439), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G33), .A2(G283), .ZN(new_n445));
  INV_X1    g0245(.A(G97), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n445), .B1(new_n446), .B2(G33), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n444), .B1(new_n214), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT20), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n448), .A2(new_n449), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n440), .B(new_n443), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n325), .B1(new_n266), .B2(new_n267), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G264), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n270), .A2(G257), .A3(new_n325), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n303), .A2(G303), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n276), .ZN(new_n459));
  XNOR2_X1  g0259(.A(KEYINPUT5), .B(G41), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n279), .A2(G1), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n462), .A2(G270), .A3(new_n275), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n339), .A2(new_n461), .A3(new_n460), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n459), .A2(new_n465), .A3(G190), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n463), .A2(new_n464), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n467), .B1(new_n276), .B2(new_n458), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n453), .B(new_n466), .C1(new_n356), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n459), .A2(new_n465), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n452), .A2(new_n470), .A3(G169), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT21), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n468), .A2(new_n452), .A3(G179), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n452), .A2(new_n470), .A3(KEYINPUT21), .A4(G169), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n469), .A2(new_n473), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT81), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n475), .A2(new_n474), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT81), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n478), .A2(new_n479), .A3(new_n473), .A4(new_n469), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT19), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n249), .B1(new_n482), .B2(new_n385), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n222), .A2(new_n446), .A3(new_n414), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n249), .A2(G33), .A3(G97), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n483), .A2(new_n484), .B1(new_n485), .B2(new_n482), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n211), .B(new_n213), .C1(new_n301), .C2(new_n302), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT79), .B1(new_n487), .B2(new_n220), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT79), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n249), .A2(new_n270), .A3(new_n489), .A4(G68), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n255), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n422), .A2(new_n258), .ZN(new_n494));
  INV_X1    g0294(.A(new_n422), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n442), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n493), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT80), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n492), .A2(new_n255), .B1(new_n258), .B2(new_n422), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT80), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(new_n500), .A3(new_n496), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n339), .A2(new_n461), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n275), .B(G250), .C1(G1), .C2(new_n279), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(G238), .B(new_n325), .C1(new_n301), .C2(new_n302), .ZN(new_n506));
  INV_X1    g0306(.A(G33), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n506), .B1(new_n507), .B2(new_n439), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT78), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n454), .A2(new_n509), .A3(G244), .ZN(new_n510));
  OAI211_X1 g0310(.A(G244), .B(G1698), .C1(new_n301), .C2(new_n302), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT78), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n508), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(G179), .B(new_n505), .C1(new_n513), .C2(new_n275), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n510), .A2(new_n512), .ZN(new_n515));
  INV_X1    g0315(.A(new_n508), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n504), .B1(new_n517), .B2(new_n276), .ZN(new_n518));
  INV_X1    g0318(.A(G169), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n514), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n498), .A2(new_n501), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n442), .A2(G97), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n258), .A2(new_n446), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT76), .ZN(new_n525));
  OR2_X1    g0325(.A1(new_n524), .A2(KEYINPUT76), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n300), .A2(G107), .A3(new_n305), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n247), .A2(G77), .ZN(new_n529));
  XNOR2_X1  g0329(.A(G97), .B(G107), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT75), .ZN(new_n531));
  OR2_X1    g0331(.A1(new_n531), .A2(KEYINPUT6), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  MUX2_X1   g0333(.A(new_n531), .B(G97), .S(KEYINPUT6), .Z(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(new_n530), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n528), .B(new_n529), .C1(new_n249), .C2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n527), .B1(new_n536), .B2(new_n255), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n462), .A2(G257), .A3(new_n275), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n464), .ZN(new_n539));
  OAI211_X1 g0339(.A(G250), .B(G1698), .C1(new_n301), .C2(new_n302), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT77), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT77), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n270), .A2(new_n542), .A3(G250), .A4(G1698), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n270), .A2(KEYINPUT4), .A3(G244), .A4(new_n325), .ZN(new_n545));
  OAI211_X1 g0345(.A(G244), .B(new_n325), .C1(new_n301), .C2(new_n302), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT4), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n546), .A2(new_n547), .B1(G33), .B2(G283), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  AOI211_X1 g0349(.A(G190), .B(new_n539), .C1(new_n549), .C2(new_n276), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n541), .A2(new_n543), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n546), .A2(new_n547), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n552), .A2(new_n545), .A3(new_n445), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n276), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n539), .ZN(new_n555));
  AOI21_X1  g0355(.A(G200), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n537), .B1(new_n550), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n529), .B1(new_n535), .B2(new_n249), .ZN(new_n558));
  INV_X1    g0358(.A(new_n528), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n255), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n527), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI211_X1 g0362(.A(new_n342), .B(new_n539), .C1(new_n549), .C2(new_n276), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n519), .B1(new_n554), .B2(new_n555), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n275), .B1(new_n515), .B2(new_n516), .ZN(new_n566));
  OAI21_X1  g0366(.A(G200), .B1(new_n566), .B2(new_n504), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n442), .A2(G87), .ZN(new_n568));
  OAI211_X1 g0368(.A(G190), .B(new_n505), .C1(new_n513), .C2(new_n275), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n499), .A2(new_n567), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n557), .A2(new_n565), .A3(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n522), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(KEYINPUT22), .B1(new_n487), .B2(new_n222), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT22), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n249), .A2(new_n270), .A3(new_n574), .A4(G87), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(KEYINPUT23), .B1(new_n210), .B2(G107), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n210), .A2(G33), .A3(G116), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(KEYINPUT23), .A2(G107), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(KEYINPUT82), .B1(new_n249), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT82), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n214), .A2(new_n583), .A3(new_n580), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n579), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT24), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n576), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n586), .B1(new_n576), .B2(new_n585), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n255), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT83), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(KEYINPUT83), .B(new_n255), .C1(new_n587), .C2(new_n588), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n376), .A2(G20), .A3(new_n414), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT25), .ZN(new_n595));
  OAI21_X1  g0395(.A(KEYINPUT84), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n595), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n594), .A2(KEYINPUT84), .A3(new_n595), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n598), .A2(new_n599), .B1(G107), .B2(new_n442), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n593), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n270), .A2(G257), .A3(G1698), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n270), .A2(G250), .A3(new_n325), .ZN(new_n603));
  INV_X1    g0403(.A(G294), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n602), .B(new_n603), .C1(new_n507), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n276), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT85), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT85), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n605), .A2(new_n608), .A3(new_n276), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n462), .A2(G264), .A3(new_n275), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n607), .A2(new_n464), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n606), .A2(new_n464), .A3(new_n610), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n611), .A2(G169), .B1(new_n613), .B2(G179), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n601), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n600), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n591), .B2(new_n592), .ZN(new_n618));
  OAI22_X1  g0418(.A1(new_n611), .A2(G190), .B1(new_n613), .B2(G200), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n481), .A2(new_n572), .A3(new_n616), .A4(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n438), .A2(new_n621), .ZN(G372));
  INV_X1    g0422(.A(new_n403), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n410), .B1(new_n623), .B2(new_n432), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n352), .B1(new_n624), .B2(new_n368), .ZN(new_n625));
  INV_X1    g0425(.A(new_n292), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n295), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n571), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n614), .B1(new_n593), .B2(new_n600), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n478), .A2(new_n473), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n629), .B(new_n620), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT86), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n563), .B2(new_n564), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n554), .A2(G179), .A3(new_n555), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n539), .B1(new_n549), .B2(new_n276), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n636), .B(KEYINPUT86), .C1(new_n519), .C2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n635), .A2(new_n562), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n520), .A2(new_n497), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n570), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n633), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n565), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n521), .A2(new_n643), .A3(KEYINPUT26), .A4(new_n570), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n632), .A2(new_n645), .A3(new_n640), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n628), .B1(new_n438), .B2(new_n646), .ZN(G369));
  INV_X1    g0447(.A(G330), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n249), .A2(new_n376), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(G213), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G343), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n481), .B1(new_n453), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n453), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n631), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n648), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n601), .A2(new_n654), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n616), .A2(new_n660), .A3(new_n620), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT87), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n662), .B1(new_n630), .B2(new_n654), .ZN(new_n663));
  NOR4_X1   g0463(.A1(new_n618), .A2(new_n614), .A3(KEYINPUT87), .A4(new_n655), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n616), .A2(new_n654), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n478), .A2(new_n473), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(new_n654), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n667), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n666), .A2(new_n670), .ZN(G399));
  INV_X1    g0471(.A(new_n207), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(G41), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n484), .A2(G116), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G1), .A3(new_n675), .ZN(new_n676));
  OAI22_X1  g0476(.A1(new_n676), .A2(KEYINPUT88), .B1(new_n216), .B2(new_n674), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(KEYINPUT88), .B2(new_n676), .ZN(new_n678));
  XOR2_X1   g0478(.A(new_n678), .B(KEYINPUT28), .Z(new_n679));
  OAI21_X1  g0479(.A(new_n505), .B1(new_n513), .B2(new_n275), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n680), .A2(new_n342), .A3(new_n470), .ZN(new_n681));
  OR3_X1    g0481(.A1(new_n681), .A2(new_n613), .A3(new_n637), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n637), .A2(G179), .A3(new_n468), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT89), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n518), .A2(new_n684), .A3(new_n606), .A4(new_n610), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n606), .A2(new_n610), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT89), .B1(new_n680), .B2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n683), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n682), .B1(new_n688), .B2(KEYINPUT30), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT30), .ZN(new_n690));
  AOI211_X1 g0490(.A(new_n690), .B(new_n683), .C1(new_n685), .C2(new_n687), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n654), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT31), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI211_X1 g0494(.A(KEYINPUT31), .B(new_n654), .C1(new_n689), .C2(new_n691), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n694), .B(new_n695), .C1(new_n621), .C2(new_n654), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n632), .A2(new_n645), .A3(new_n640), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT29), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(new_n699), .A3(new_n655), .ZN(new_n700));
  INV_X1    g0500(.A(new_n640), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n571), .B1(new_n618), .B2(new_n619), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n668), .B1(new_n614), .B2(new_n618), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(KEYINPUT26), .B1(new_n639), .B2(new_n641), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n521), .A2(new_n643), .A3(new_n633), .A4(new_n570), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n654), .B1(new_n704), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n700), .B1(new_n709), .B2(new_n699), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n697), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n679), .B1(new_n711), .B2(G1), .ZN(G364));
  NOR2_X1   g0512(.A1(G13), .A2(G33), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G20), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n656), .A2(new_n658), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n254), .B1(G20), .B2(new_n519), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n214), .A2(new_n354), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n719), .A2(G179), .A3(new_n356), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n720), .A2(KEYINPUT91), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(KEYINPUT91), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n342), .A2(new_n354), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n214), .A2(G200), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT92), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n723), .A2(G283), .B1(G326), .B2(new_n727), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n719), .A2(new_n342), .A3(G200), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G311), .ZN(new_n730));
  NOR4_X1   g0530(.A1(new_n210), .A2(new_n354), .A3(new_n356), .A4(G179), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT93), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n731), .B(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n214), .A2(new_n356), .A3(new_n724), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n734), .A2(G303), .B1(G322), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G179), .A2(G200), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n249), .B1(G190), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n303), .B1(new_n739), .B2(new_n604), .ZN(new_n740));
  INV_X1    g0540(.A(new_n719), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(G179), .A3(G200), .ZN(new_n742));
  XOR2_X1   g0542(.A(KEYINPUT33), .B(G317), .Z(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n741), .A2(new_n738), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n740), .B(new_n744), .C1(G329), .C2(new_n746), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n728), .A2(new_n730), .A3(new_n737), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n723), .A2(G107), .ZN(new_n749));
  INV_X1    g0549(.A(new_n729), .ZN(new_n750));
  OAI22_X1  g0550(.A1(new_n750), .A2(new_n203), .B1(new_n742), .B2(new_n220), .ZN(new_n751));
  INV_X1    g0551(.A(new_n731), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n270), .B1(new_n752), .B2(new_n222), .C1(new_n446), .C2(new_n739), .ZN(new_n753));
  INV_X1    g0553(.A(G58), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n260), .A2(new_n725), .B1(new_n735), .B2(new_n754), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n751), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G159), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n745), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT32), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n749), .A2(new_n756), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n718), .B1(new_n748), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n715), .A2(new_n717), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n672), .A2(new_n303), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT90), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n765), .A2(G355), .B1(new_n439), .B2(new_n672), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n672), .A2(new_n270), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n768), .B1(new_n279), .B2(new_n217), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(new_n245), .B2(new_n279), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n763), .B1(new_n766), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n214), .A2(new_n257), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n261), .B1(new_n772), .B2(G45), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n673), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n761), .A2(new_n771), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n716), .A2(new_n777), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT94), .Z(new_n779));
  INV_X1    g0579(.A(new_n659), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n656), .A2(new_n648), .A3(new_n658), .ZN(new_n781));
  AND3_X1   g0581(.A1(new_n780), .A2(new_n776), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(G396));
  NOR2_X1   g0584(.A1(new_n432), .A2(new_n654), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n435), .B1(new_n433), .B2(new_n655), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n785), .B1(new_n432), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(new_n646), .B2(new_n654), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n432), .A2(new_n435), .A3(new_n655), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n698), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n696), .A2(G330), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n775), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n794), .B2(new_n793), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n717), .A2(new_n713), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT95), .Z(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n776), .B1(new_n203), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT97), .B(G143), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n729), .A2(G159), .B1(new_n736), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G137), .ZN(new_n803));
  INV_X1    g0603(.A(G150), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n802), .B1(new_n803), .B2(new_n725), .C1(new_n804), .C2(new_n742), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT34), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G132), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n733), .A2(new_n260), .B1(new_n808), .B2(new_n745), .ZN(new_n809));
  INV_X1    g0609(.A(new_n739), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n303), .B(new_n809), .C1(G58), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n805), .A2(new_n806), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n723), .A2(G68), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n807), .A2(new_n811), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G311), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n750), .A2(new_n439), .B1(new_n745), .B2(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n270), .B(new_n816), .C1(G97), .C2(new_n810), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n723), .A2(G87), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n719), .A2(new_n342), .A3(new_n356), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n819), .A2(KEYINPUT96), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(KEYINPUT96), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(G283), .ZN(new_n824));
  INV_X1    g0624(.A(G303), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n604), .A2(new_n735), .B1(new_n725), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n734), .B2(G107), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n817), .A2(new_n818), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n814), .A2(new_n828), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n800), .B1(new_n718), .B2(new_n829), .C1(new_n787), .C2(new_n714), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n796), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(G384));
  NOR2_X1   g0632(.A1(new_n772), .A2(new_n261), .ZN(new_n833));
  AOI21_X1  g0633(.A(KEYINPUT16), .B1(new_n322), .B2(new_n311), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n298), .B1(new_n361), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n652), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n353), .B2(new_n368), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n652), .B(new_n335), .C1(new_n341), .C2(new_n342), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n365), .A2(new_n366), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(KEYINPUT37), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT101), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n842), .A2(KEYINPUT101), .A3(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n345), .A2(KEYINPUT37), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n324), .A2(new_n652), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n848), .A2(new_n365), .A3(new_n366), .A4(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT102), .B1(new_n847), .B2(new_n851), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n842), .A2(KEYINPUT101), .A3(KEYINPUT37), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT101), .B1(new_n842), .B2(KEYINPUT37), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n851), .B(KEYINPUT102), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n839), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT38), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n851), .B1(new_n853), .B2(new_n854), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT102), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n838), .B1(new_n862), .B2(new_n855), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT38), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n382), .A2(new_n654), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n411), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n403), .A2(new_n410), .A3(new_n866), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n696), .A2(new_n787), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT40), .B1(new_n865), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n368), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n849), .B1(new_n873), .B2(new_n352), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n345), .B(new_n849), .C1(new_n324), .C2(new_n358), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT37), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n851), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n864), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n696), .A2(new_n870), .A3(KEYINPUT40), .A4(new_n787), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n872), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n437), .A2(new_n696), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n648), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n883), .B2(new_n884), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n836), .B1(new_n350), .B2(new_n351), .ZN(new_n887));
  INV_X1    g0687(.A(new_n870), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n790), .B1(new_n704), .B2(new_n645), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT100), .B1(new_n889), .B2(new_n785), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT100), .ZN(new_n891));
  INV_X1    g0691(.A(new_n785), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n792), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n888), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n887), .B1(new_n894), .B2(new_n865), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n859), .A2(KEYINPUT39), .A3(new_n864), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n858), .B(new_n838), .C1(new_n862), .C2(new_n855), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n897), .B1(new_n898), .B2(new_n878), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n410), .A2(new_n654), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n896), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n895), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n627), .B1(new_n710), .B2(new_n437), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n902), .B(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n833), .B1(new_n886), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n904), .B2(new_n886), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n249), .A2(new_n439), .A3(new_n254), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n535), .B(KEYINPUT98), .Z(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT35), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n910), .B2(new_n909), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n912), .B(KEYINPUT36), .Z(new_n913));
  NOR2_X1   g0713(.A1(new_n201), .A2(new_n220), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n203), .B(new_n216), .C1(G58), .C2(G68), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n914), .B1(new_n915), .B2(KEYINPUT99), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(KEYINPUT99), .B2(new_n915), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(G1), .A3(new_n257), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n906), .A2(new_n913), .A3(new_n918), .ZN(G367));
  OR2_X1    g0719(.A1(new_n639), .A2(new_n655), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n565), .B(new_n557), .C1(new_n537), .C2(new_n655), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n630), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n654), .B1(new_n923), .B2(new_n565), .ZN(new_n924));
  INV_X1    g0724(.A(new_n669), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT87), .B1(new_n616), .B2(new_n655), .ZN(new_n926));
  INV_X1    g0726(.A(new_n664), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n925), .B1(new_n928), .B2(new_n661), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n922), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n924), .B1(new_n930), .B2(KEYINPUT42), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n665), .A2(new_n669), .ZN(new_n932));
  INV_X1    g0732(.A(new_n922), .ZN(new_n933));
  OR3_X1    g0733(.A1(new_n932), .A2(KEYINPUT42), .A3(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT103), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n931), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n499), .A2(new_n568), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n654), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n940), .A2(new_n640), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n940), .A2(new_n640), .A3(new_n570), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT43), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n938), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n666), .A2(new_n933), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n934), .B(new_n935), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n950), .A2(new_n945), .A3(new_n944), .A4(new_n931), .ZN(new_n951));
  AND3_X1   g0751(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n949), .B1(new_n948), .B2(new_n951), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n673), .B(KEYINPUT41), .Z(new_n955));
  INV_X1    g0755(.A(new_n667), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n932), .A2(new_n956), .A3(new_n922), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT45), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n670), .A2(KEYINPUT45), .A3(new_n922), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI211_X1 g0761(.A(KEYINPUT44), .B(new_n933), .C1(new_n929), .C2(new_n667), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT44), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n670), .B2(new_n922), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n666), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n961), .A2(new_n965), .A3(new_n666), .ZN(new_n969));
  INV_X1    g0769(.A(new_n710), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n928), .A2(new_n661), .A3(new_n925), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n780), .B1(new_n972), .B2(new_n929), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n971), .A2(new_n932), .A3(new_n659), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n970), .A2(new_n973), .A3(new_n794), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT104), .ZN(new_n976));
  INV_X1    g0776(.A(new_n974), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n659), .B1(new_n971), .B2(new_n932), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT104), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n979), .A2(new_n980), .A3(new_n711), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n968), .A2(new_n969), .A3(new_n976), .A4(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n955), .B1(new_n982), .B2(new_n711), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT105), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n773), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI211_X1 g0785(.A(KEYINPUT105), .B(new_n955), .C1(new_n982), .C2(new_n711), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n954), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n237), .A2(new_n767), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n763), .B1(new_n672), .B2(new_n495), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n776), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n715), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n723), .A2(G97), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G294), .B2(new_n823), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n734), .A2(KEYINPUT46), .A3(G116), .ZN(new_n994));
  INV_X1    g0794(.A(G317), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n994), .B1(new_n995), .B2(new_n745), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n752), .A2(new_n439), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n303), .B1(new_n414), .B2(new_n739), .C1(new_n997), .C2(KEYINPUT46), .ZN(new_n998));
  INV_X1    g0798(.A(G283), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n750), .A2(new_n999), .B1(new_n825), .B2(new_n735), .ZN(new_n1000));
  NOR3_X1   g0800(.A1(new_n996), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n993), .B(new_n1001), .C1(new_n815), .C2(new_n726), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n729), .A2(new_n201), .B1(new_n736), .B2(G150), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n803), .B2(new_n745), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n739), .A2(new_n220), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n270), .B1(new_n752), .B2(new_n754), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n823), .A2(G159), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n727), .A2(new_n801), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n723), .A2(G77), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1002), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT47), .Z(new_n1013));
  OAI221_X1 g0813(.A(new_n990), .B1(new_n991), .B2(new_n943), .C1(new_n1013), .C2(new_n718), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT106), .Z(new_n1015));
  NAND2_X1  g0815(.A1(new_n987), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT107), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1016), .B(new_n1017), .ZN(G387));
  OAI22_X1  g0818(.A1(new_n977), .A2(new_n978), .B1(new_n697), .B2(new_n710), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n975), .A2(new_n1019), .A3(new_n673), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n739), .A2(new_n422), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G50), .B2(new_n736), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT111), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n725), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n729), .A2(G68), .B1(new_n1024), .B2(G159), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n251), .B2(new_n742), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n270), .B1(new_n752), .B2(new_n203), .C1(new_n745), .C2(new_n804), .ZN(new_n1027));
  OR4_X1    g0827(.A1(new_n992), .A2(new_n1023), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n727), .A2(G322), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n729), .A2(G303), .B1(new_n736), .B2(G317), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1029), .B(new_n1030), .C1(new_n822), .C2(new_n815), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT48), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n810), .A2(G283), .B1(new_n731), .B2(G294), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(KEYINPUT112), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT112), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1033), .A2(new_n1039), .A3(new_n1036), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1038), .A2(KEYINPUT49), .A3(new_n1040), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n723), .A2(G116), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n270), .B(new_n1042), .C1(G326), .C2(new_n746), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(KEYINPUT49), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1028), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n717), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n928), .A2(new_n661), .A3(new_n715), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n675), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n765), .A2(new_n1049), .B1(new_n414), .B2(new_n672), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n234), .A2(new_n279), .ZN(new_n1051));
  XOR2_X1   g0851(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n1052));
  OR3_X1    g0852(.A1(new_n1052), .A2(G50), .A3(new_n251), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n279), .B1(new_n220), .B2(new_n203), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n675), .B2(KEYINPUT108), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n675), .A2(KEYINPUT108), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1052), .B1(G50), .B2(new_n251), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n767), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1050), .B1(new_n1051), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT110), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1062), .A2(new_n762), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n776), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AND3_X1   g0865(.A1(new_n1047), .A2(new_n1048), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n979), .B2(new_n774), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1020), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT113), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1020), .A2(new_n1067), .A3(KEYINPUT113), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(G393));
  AND3_X1   g0872(.A1(new_n961), .A2(new_n965), .A3(new_n666), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n666), .B1(new_n961), .B2(new_n965), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n975), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n982), .A2(new_n1075), .A3(new_n673), .ZN(new_n1076));
  OAI21_X1  g0876(.A(KEYINPUT114), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT114), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n968), .A2(new_n1078), .A3(new_n969), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1077), .A2(new_n1079), .A3(new_n774), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n922), .A2(new_n991), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT115), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n242), .A2(new_n768), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n762), .B1(new_n446), .B2(new_n207), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n775), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n815), .A2(new_n735), .B1(new_n725), .B2(new_n995), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1086), .B(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n823), .A2(G303), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n303), .B1(new_n752), .B2(new_n999), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n746), .B2(G322), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G294), .A2(new_n729), .B1(new_n810), .B2(G116), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1089), .A2(new_n749), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n823), .A2(new_n201), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n270), .B1(new_n752), .B2(new_n220), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n746), .B2(new_n801), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n424), .A2(new_n729), .B1(new_n810), .B2(G77), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1094), .A2(new_n818), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n804), .A2(new_n725), .B1(new_n735), .B2(new_n757), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT51), .Z(new_n1100));
  OAI22_X1  g0900(.A1(new_n1088), .A2(new_n1093), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1085), .B1(new_n1101), .B2(new_n717), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1082), .A2(new_n1102), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n1080), .A2(KEYINPUT117), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT117), .B1(new_n1080), .B2(new_n1103), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1076), .B1(new_n1104), .B2(new_n1105), .ZN(G390));
  NAND4_X1  g0906(.A1(new_n696), .A2(new_n870), .A3(G330), .A4(new_n787), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n891), .B1(new_n792), .B2(new_n892), .ZN(new_n1109));
  AOI211_X1 g0909(.A(KEYINPUT100), .B(new_n785), .C1(new_n698), .C2(new_n791), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n870), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n900), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n899), .A2(new_n896), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n786), .A2(new_n432), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n785), .B1(new_n709), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1115), .A2(new_n888), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n878), .B1(new_n863), .B2(KEYINPUT38), .ZN(new_n1117));
  NOR3_X1   g0917(.A1(new_n1116), .A2(new_n1117), .A3(new_n900), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1108), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n880), .B(new_n1112), .C1(new_n888), .C2(new_n1115), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n896), .A2(new_n899), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n894), .A2(new_n900), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1107), .B(new_n1120), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1119), .A2(new_n1123), .A3(new_n774), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n775), .B1(new_n798), .B2(new_n424), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n735), .A2(new_n808), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n731), .A2(G150), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT53), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1126), .B(new_n1128), .C1(G128), .C2(new_n1024), .ZN(new_n1129));
  INV_X1    g0929(.A(G125), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n745), .A2(new_n1130), .B1(new_n739), .B2(new_n757), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT54), .B(G143), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n303), .B(new_n1131), .C1(new_n729), .C2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n823), .A2(G137), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n723), .A2(new_n201), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1129), .A2(new_n1134), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n739), .A2(new_n203), .B1(new_n735), .B2(new_n439), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n723), .A2(G68), .B1(KEYINPUT119), .B2(new_n1138), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(KEYINPUT119), .B2(new_n1138), .C1(new_n414), .C2(new_n822), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n270), .B1(new_n734), .B2(G87), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n729), .A2(G97), .B1(new_n1024), .B2(G283), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(new_n604), .C2(new_n745), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1137), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1125), .B1(new_n1144), .B2(new_n717), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n1121), .B2(new_n714), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n697), .A2(new_n437), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n628), .B(new_n1147), .C1(new_n438), .C2(new_n970), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n696), .A2(G330), .A3(new_n787), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n888), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1150), .A2(new_n1107), .B1(new_n893), .B2(new_n890), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1150), .A2(new_n1107), .A3(new_n1115), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1148), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1119), .A2(new_n1123), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT118), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(new_n1156), .A3(new_n673), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1119), .A2(new_n1123), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1148), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1157), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1156), .B1(new_n1155), .B2(new_n673), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1124), .B(new_n1146), .C1(new_n1163), .C2(new_n1164), .ZN(G378));
  NAND2_X1  g0965(.A1(new_n1155), .A2(new_n1160), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n264), .A2(new_n836), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n296), .B(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1168), .B(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(G330), .B1(new_n1117), .B2(new_n881), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n872), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1169), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1168), .B(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n863), .A2(KEYINPUT38), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n871), .B1(new_n1175), .B2(new_n898), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT40), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n648), .B1(new_n880), .B2(new_n882), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1174), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n902), .B1(new_n1172), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1170), .B1(new_n872), .B2(new_n1171), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n895), .A2(new_n901), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1178), .A2(new_n1174), .A3(new_n1179), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1181), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1166), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT57), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1188), .B1(new_n1155), .B2(new_n1160), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT121), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n1181), .B2(new_n1185), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1185), .A2(new_n1191), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1190), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1189), .A2(new_n1195), .A3(new_n673), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1186), .A2(new_n774), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n797), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n775), .B1(new_n201), .B2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n270), .A2(G41), .ZN(new_n1200));
  AOI211_X1 g1000(.A(G50), .B(new_n1200), .C1(new_n507), .C2(new_n278), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n723), .A2(G58), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n750), .A2(new_n422), .B1(new_n742), .B2(new_n446), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G116), .B2(new_n1024), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1200), .B1(new_n752), .B2(new_n203), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1205), .A2(new_n1005), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n746), .A2(G283), .B1(new_n736), .B2(G107), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1202), .A2(new_n1204), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT58), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1201), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G137), .A2(new_n729), .B1(new_n810), .B2(G150), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n819), .A2(G132), .B1(new_n1024), .B2(G125), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n736), .A2(G128), .B1(new_n731), .B2(new_n1133), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n723), .A2(G159), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1217));
  AOI211_X1 g1017(.A(G33), .B(G41), .C1(new_n746), .C2(G124), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1210), .B1(new_n1209), .B2(new_n1208), .C1(new_n1215), .C2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1199), .B1(new_n1220), .B2(new_n717), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n1170), .B2(new_n714), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT120), .Z(new_n1223));
  AND2_X1   g1023(.A1(new_n1197), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1196), .A2(new_n1224), .ZN(G375));
  INV_X1    g1025(.A(new_n955), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1152), .A2(new_n1148), .A3(new_n1153), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1161), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n888), .A2(new_n713), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n775), .B1(new_n798), .B2(G68), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n823), .A2(new_n1133), .ZN(new_n1231));
  INV_X1    g1031(.A(G128), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n745), .A2(new_n1232), .B1(new_n803), .B2(new_n735), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(G150), .B2(new_n729), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n739), .A2(new_n260), .B1(new_n725), .B2(new_n808), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n303), .B(new_n1235), .C1(new_n734), .C2(G159), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1231), .A2(new_n1202), .A3(new_n1234), .A4(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1010), .A2(new_n303), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1238), .A2(KEYINPUT123), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(KEYINPUT123), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n733), .A2(new_n446), .B1(new_n825), .B2(new_n745), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1021), .B(new_n1241), .C1(G283), .C2(new_n736), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1239), .A2(new_n1240), .A3(new_n1242), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n729), .A2(G107), .B1(new_n1024), .B2(G294), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n822), .B2(new_n439), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT122), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1237), .B1(new_n1243), .B2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1230), .B1(new_n1247), .B2(new_n717), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1159), .A2(new_n774), .B1(new_n1229), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1228), .A2(new_n1249), .ZN(G381));
  NAND3_X1  g1050(.A1(new_n1070), .A2(new_n783), .A3(new_n1071), .ZN(new_n1251));
  OR4_X1    g1051(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1251), .ZN(new_n1252));
  OR4_X1    g1052(.A1(G387), .A2(new_n1252), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1053(.A(G378), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n653), .ZN(new_n1255));
  OAI211_X1 g1055(.A(G407), .B(G213), .C1(G375), .C2(new_n1255), .ZN(G409));
  AND2_X1   g1056(.A1(new_n987), .A2(new_n1015), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n783), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT107), .B1(new_n1259), .B2(new_n1251), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(G390), .A2(new_n1260), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1070), .A2(new_n783), .A3(new_n1071), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1262), .A2(new_n1258), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1080), .A2(new_n1103), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT117), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1080), .A2(KEYINPUT117), .A3(new_n1103), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1263), .B1(new_n1268), .B2(new_n1076), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1257), .B1(new_n1261), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1263), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(G390), .A2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1017), .B1(new_n1262), .B2(new_n1258), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1268), .A2(new_n1076), .A3(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1272), .A2(new_n1016), .A3(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1270), .A2(new_n1275), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1150), .A2(new_n1107), .A3(new_n1115), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1277), .A2(new_n1151), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT60), .B1(new_n1278), .B2(new_n1148), .ZN(new_n1279));
  OAI21_X1  g1079(.A(KEYINPUT125), .B1(new_n1279), .B2(new_n1154), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT60), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1227), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT125), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1282), .A2(new_n1161), .A3(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1152), .A2(new_n1148), .A3(KEYINPUT60), .A4(new_n1153), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1285), .A2(new_n673), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1280), .A2(new_n1284), .A3(new_n1286), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1287), .A2(G384), .A3(new_n1249), .ZN(new_n1288));
  AOI21_X1  g1088(.A(G384), .B1(new_n1287), .B2(new_n1249), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n653), .A2(G213), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(G2897), .ZN(new_n1293));
  OR2_X1    g1093(.A1(new_n1291), .A2(KEYINPUT126), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1290), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1287), .A2(new_n1249), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n831), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1287), .A2(G384), .A3(new_n1249), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1297), .A2(new_n1298), .A3(new_n1294), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1293), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1295), .A2(new_n1301), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1196), .A2(G378), .A3(new_n1224), .ZN(new_n1303));
  OAI21_X1  g1103(.A(KEYINPUT124), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1183), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1306));
  OAI21_X1  g1106(.A(KEYINPUT121), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT124), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1307), .A2(new_n1308), .A3(new_n1193), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1304), .A2(new_n1309), .A3(new_n774), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1166), .A2(new_n1226), .A3(new_n1186), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1311), .A2(new_n1223), .ZN(new_n1312));
  AOI21_X1  g1112(.A(G378), .B1(new_n1310), .B2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1291), .B1(new_n1303), .B2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(KEYINPUT61), .B1(new_n1302), .B2(new_n1314), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1291), .B(new_n1290), .C1(new_n1303), .C2(new_n1313), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(KEYINPUT62), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1315), .A2(new_n1317), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1316), .A2(KEYINPUT62), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1276), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT61), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1254), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1196), .A2(G378), .A3(new_n1224), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1292), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1295), .A2(new_n1301), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1321), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT63), .ZN(new_n1328));
  NOR3_X1   g1128(.A1(new_n1288), .A2(new_n1289), .A3(new_n1328), .ZN(new_n1329));
  OAI211_X1 g1129(.A(new_n1291), .B(new_n1329), .C1(new_n1303), .C2(new_n1313), .ZN(new_n1330));
  AND3_X1   g1130(.A1(new_n1272), .A2(new_n1016), .A3(new_n1274), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1016), .B1(new_n1274), .B2(new_n1272), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1330), .A2(new_n1333), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1327), .A2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1316), .A2(new_n1328), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT127), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1276), .B1(new_n1325), .B2(new_n1329), .ZN(new_n1338));
  AND4_X1   g1138(.A1(KEYINPUT127), .A2(new_n1315), .A3(new_n1338), .A4(new_n1336), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1320), .B1(new_n1337), .B2(new_n1339), .ZN(G405));
  XNOR2_X1  g1140(.A(G375), .B(G378), .ZN(new_n1341));
  XNOR2_X1  g1141(.A(new_n1341), .B(new_n1290), .ZN(new_n1342));
  XNOR2_X1  g1142(.A(new_n1342), .B(new_n1333), .ZN(G402));
endmodule


