//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n629, new_n630,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AND2_X1   g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n456), .A2(KEYINPUT66), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n453), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(KEYINPUT66), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OR2_X1    g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(new_n462), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n463), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n462), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n469), .A2(new_n472), .ZN(G160));
  OAI21_X1  g048(.A(KEYINPUT68), .B1(G100), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NOR3_X1   g050(.A1(KEYINPUT68), .A2(G100), .A3(G2105), .ZN(new_n476));
  OAI221_X1 g051(.A(G2104), .B1(G112), .B2(new_n462), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT69), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n464), .A2(new_n465), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(new_n462), .ZN(new_n480));
  OR2_X1    g055(.A1(new_n480), .A2(KEYINPUT67), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(KEYINPUT67), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n479), .A2(G2105), .ZN(new_n486));
  AOI211_X1 g061(.A(new_n478), .B(new_n485), .C1(G136), .C2(new_n486), .ZN(G162));
  NAND2_X1  g062(.A1(new_n480), .A2(G126), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n462), .A2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  OR2_X1    g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT4), .B1(new_n467), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n486), .A2(new_n495), .A3(G138), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n492), .B1(new_n494), .B2(new_n496), .ZN(G164));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(KEYINPUT5), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT71), .B1(new_n500), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(new_n498), .A3(KEYINPUT5), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(KEYINPUT6), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT70), .B1(new_n507), .B2(G651), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(new_n505), .A3(KEYINPUT6), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n506), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n504), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n517), .A2(new_n505), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n516), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n521));
  AOI211_X1 g096(.A(new_n521), .B(new_n499), .C1(new_n501), .C2(new_n503), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n501), .A2(new_n503), .ZN(new_n523));
  INV_X1    g098(.A(new_n499), .ZN(new_n524));
  AOI21_X1  g099(.A(KEYINPUT72), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(G63), .A2(G651), .ZN(new_n526));
  NOR3_X1   g101(.A1(new_n522), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n511), .A2(G51), .A3(G543), .ZN(new_n528));
  OR2_X1    g103(.A1(KEYINPUT73), .A2(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(KEYINPUT73), .A2(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n529), .A2(new_n532), .A3(new_n530), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  OAI211_X1 g112(.A(new_n528), .B(new_n536), .C1(new_n512), .C2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n527), .A2(new_n538), .ZN(G168));
  AOI21_X1  g114(.A(new_n502), .B1(KEYINPUT5), .B2(new_n498), .ZN(new_n540));
  NOR3_X1   g115(.A1(new_n500), .A2(KEYINPUT71), .A3(G543), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n524), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(new_n521), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n504), .A2(KEYINPUT72), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n543), .A2(G64), .A3(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(G77), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n498), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n505), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n504), .A2(new_n511), .ZN(new_n550));
  XOR2_X1   g125(.A(KEYINPUT74), .B(G90), .Z(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(G52), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n553), .B2(new_n514), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n549), .A2(new_n554), .ZN(G171));
  NAND3_X1  g130(.A1(new_n543), .A2(G56), .A3(new_n544), .ZN(new_n556));
  AND2_X1   g131(.A1(G68), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n505), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(G81), .ZN(new_n560));
  INV_X1    g135(.A(G43), .ZN(new_n561));
  OAI22_X1  g136(.A1(new_n512), .A2(new_n560), .B1(new_n514), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  INV_X1    g143(.A(new_n514), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n569), .A2(new_n570), .A3(G53), .ZN(new_n571));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT9), .B1(new_n514), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n550), .A2(G91), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n504), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n576));
  OAI211_X1 g151(.A(new_n574), .B(new_n575), .C1(new_n505), .C2(new_n576), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  AND2_X1   g153(.A1(new_n528), .A2(new_n536), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n550), .A2(G89), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n543), .A2(new_n544), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n526), .ZN(G286));
  INV_X1    g157(.A(G87), .ZN(new_n583));
  INV_X1    g158(.A(G49), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n512), .A2(new_n583), .B1(new_n514), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(G74), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n585), .B1(new_n587), .B2(G651), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G288));
  INV_X1    g164(.A(G86), .ZN(new_n590));
  INV_X1    g165(.A(G48), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n512), .A2(new_n590), .B1(new_n514), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n504), .A2(G61), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT75), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n505), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G305));
  NOR2_X1   g173(.A1(new_n522), .A2(new_n525), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n505), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  INV_X1    g177(.A(G47), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n512), .A2(new_n602), .B1(new_n514), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G290));
  OR2_X1    g181(.A1(new_n514), .A2(KEYINPUT77), .ZN(new_n607));
  INV_X1    g182(.A(G54), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(new_n514), .B2(KEYINPUT77), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT78), .Z(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT79), .B(G66), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n542), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n607), .A2(new_n609), .B1(new_n613), .B2(G651), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n504), .A2(new_n511), .A3(G92), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(KEYINPUT76), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT76), .ZN(new_n618));
  NAND4_X1  g193(.A1(new_n504), .A2(new_n511), .A3(new_n618), .A4(G92), .ZN(new_n619));
  AND3_X1   g194(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n617), .B1(new_n616), .B2(new_n619), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n614), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G868), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(new_n623), .B2(G171), .ZN(G284));
  OAI21_X1  g200(.A(new_n624), .B1(new_n623), .B2(G171), .ZN(G321));
  NAND2_X1  g201(.A1(G286), .A2(G868), .ZN(new_n627));
  INV_X1    g202(.A(G91), .ZN(new_n628));
  OAI22_X1  g203(.A1(new_n576), .A2(new_n505), .B1(new_n512), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(new_n573), .B2(new_n571), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n627), .B1(G868), .B2(new_n630), .ZN(G297));
  OAI21_X1  g206(.A(new_n627), .B1(G868), .B2(new_n630), .ZN(G280));
  INV_X1    g207(.A(new_n622), .ZN(new_n633));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(G860), .ZN(G148));
  NOR2_X1   g210(.A1(new_n563), .A2(G868), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n633), .A2(new_n634), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n636), .B1(new_n637), .B2(G868), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT80), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g215(.A1(new_n486), .A2(G135), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n462), .A2(G111), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  INV_X1    g218(.A(G123), .ZN(new_n644));
  OAI221_X1 g219(.A(new_n641), .B1(new_n642), .B2(new_n643), .C1(new_n483), .C2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT81), .B(G2096), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT13), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2100), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n647), .A2(new_n651), .ZN(G156));
  XNOR2_X1  g227(.A(G2427), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(KEYINPUT14), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT82), .Z(new_n666));
  OAI21_X1  g241(.A(G14), .B1(new_n663), .B2(new_n664), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(G401));
  XOR2_X1   g243(.A(G2067), .B(G2678), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT83), .ZN(new_n670));
  NOR2_X1   g245(.A1(G2072), .A2(G2078), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n442), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2084), .B(G2090), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT18), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n672), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n672), .B(KEYINPUT17), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n676), .B(new_n673), .C1(new_n670), .C2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n673), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n670), .A2(new_n679), .A3(new_n677), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n675), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT84), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT85), .ZN(new_n684));
  XOR2_X1   g259(.A(G2096), .B(G2100), .Z(new_n685));
  OR2_X1    g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(G227));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  XOR2_X1   g264(.A(G1961), .B(G1966), .Z(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(KEYINPUT86), .ZN(new_n693));
  XOR2_X1   g268(.A(G1971), .B(G1976), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT19), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT86), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n693), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT20), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n689), .A2(new_n690), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT87), .ZN(new_n702));
  OR3_X1    g277(.A1(new_n695), .A2(new_n692), .A3(new_n700), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n699), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT88), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1991), .B(G1996), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n706), .A2(new_n709), .ZN(new_n712));
  AND3_X1   g287(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n711), .B1(new_n710), .B2(new_n712), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(G229));
  AND2_X1   g290(.A1(new_n466), .A2(G127), .ZN(new_n716));
  AND2_X1   g291(.A1(G115), .A2(G2104), .ZN(new_n717));
  OAI21_X1  g292(.A(G2105), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(KEYINPUT96), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(KEYINPUT96), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT25), .ZN(new_n721));
  NAND2_X1  g296(.A1(G103), .A2(G2104), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(G2105), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n462), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n486), .A2(G139), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n719), .A2(new_n720), .A3(new_n725), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT97), .Z(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n728), .B2(G33), .ZN(new_n730));
  INV_X1    g305(.A(G2072), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n732), .A2(KEYINPUT100), .ZN(new_n733));
  NOR2_X1   g308(.A1(G29), .A2(G35), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G162), .B2(G29), .ZN(new_n735));
  INV_X1    g310(.A(G2090), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT105), .B(KEYINPUT29), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n732), .A2(KEYINPUT100), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n733), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n730), .A2(new_n731), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT98), .Z(new_n743));
  NOR2_X1   g318(.A1(G27), .A2(G29), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G164), .B2(G29), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(G2078), .ZN(new_n746));
  AND2_X1   g321(.A1(KEYINPUT24), .A2(G34), .ZN(new_n747));
  NOR2_X1   g322(.A1(KEYINPUT24), .A2(G34), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n728), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT99), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G160), .B2(G29), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n751), .A2(G2084), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT104), .Z(new_n753));
  AOI211_X1 g328(.A(new_n746), .B(new_n753), .C1(G2084), .C2(new_n751), .ZN(new_n754));
  NOR2_X1   g329(.A1(G5), .A2(G16), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT102), .ZN(new_n756));
  INV_X1    g331(.A(G16), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(G301), .B2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G1961), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n757), .A2(G20), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT23), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n630), .B2(new_n757), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(G1956), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n728), .A2(G32), .ZN(new_n765));
  AND3_X1   g340(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n766));
  NAND3_X1  g341(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT26), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n766), .B(new_n768), .C1(G141), .C2(new_n486), .ZN(new_n769));
  INV_X1    g344(.A(G129), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n483), .B2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n765), .B1(new_n772), .B2(new_n728), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT27), .B(G1996), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G2078), .B2(new_n745), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n754), .A2(new_n760), .A3(new_n764), .A4(new_n776), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n741), .A2(new_n743), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n757), .A2(G4), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n633), .B2(new_n757), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1348), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n728), .A2(G26), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT28), .ZN(new_n783));
  OAI21_X1  g358(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n784));
  INV_X1    g359(.A(G116), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(G2105), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(G140), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n467), .B2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT94), .ZN(new_n790));
  INV_X1    g365(.A(G128), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n483), .B2(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n481), .A2(new_n482), .A3(KEYINPUT94), .A4(G128), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n789), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n783), .B1(new_n794), .B2(new_n728), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G2067), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n757), .A2(G19), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n563), .B2(new_n757), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1341), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n781), .A2(new_n796), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT95), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT30), .B(G28), .ZN(new_n802));
  OR2_X1    g377(.A1(KEYINPUT31), .A2(G11), .ZN(new_n803));
  NAND2_X1  g378(.A1(KEYINPUT31), .A2(G11), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n802), .A2(new_n728), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n645), .B2(new_n728), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT101), .Z(new_n807));
  NAND2_X1  g382(.A1(new_n757), .A2(G21), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G168), .B2(new_n757), .ZN(new_n809));
  INV_X1    g384(.A(G1966), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n807), .B(new_n811), .C1(new_n759), .C2(new_n758), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT103), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n778), .A2(new_n801), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n757), .A2(G24), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n605), .B2(new_n757), .ZN(new_n816));
  INV_X1    g391(.A(G1986), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n484), .A2(G119), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n486), .A2(G131), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT89), .Z(new_n821));
  INV_X1    g396(.A(G95), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n822), .A2(new_n462), .A3(KEYINPUT90), .ZN(new_n823));
  AOI21_X1  g398(.A(KEYINPUT90), .B1(new_n822), .B2(new_n462), .ZN(new_n824));
  OAI221_X1 g399(.A(G2104), .B1(G107), .B2(new_n462), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n819), .A2(new_n821), .A3(new_n825), .ZN(new_n826));
  MUX2_X1   g401(.A(G25), .B(new_n826), .S(G29), .Z(new_n827));
  XOR2_X1   g402(.A(KEYINPUT35), .B(G1991), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n757), .A2(G23), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n588), .B2(new_n757), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT33), .B(G1976), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT91), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n831), .B(new_n833), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT92), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n831), .B(new_n833), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT92), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n757), .A2(G22), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(G303), .B2(G16), .ZN(new_n840));
  INV_X1    g415(.A(G1971), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(G6), .A2(G16), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n597), .B2(G16), .ZN(new_n844));
  XNOR2_X1  g419(.A(KEYINPUT32), .B(G1981), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  AND3_X1   g422(.A1(new_n835), .A2(new_n838), .A3(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n818), .B(new_n829), .C1(new_n849), .C2(KEYINPUT34), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT93), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(KEYINPUT34), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(KEYINPUT36), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT36), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n851), .A2(new_n855), .A3(new_n852), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n814), .B1(new_n854), .B2(new_n856), .ZN(G311));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n856), .ZN(new_n858));
  INV_X1    g433(.A(new_n814), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(G150));
  NAND2_X1  g435(.A1(new_n633), .A2(G559), .ZN(new_n861));
  XOR2_X1   g436(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n862));
  XOR2_X1   g437(.A(new_n861), .B(new_n862), .Z(new_n863));
  NAND2_X1  g438(.A1(new_n556), .A2(new_n558), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(G651), .ZN(new_n865));
  INV_X1    g440(.A(G67), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n522), .A2(new_n525), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(G80), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n868), .A2(new_n498), .ZN(new_n869));
  OAI21_X1  g444(.A(G651), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n562), .ZN(new_n871));
  INV_X1    g446(.A(G93), .ZN(new_n872));
  INV_X1    g447(.A(G55), .ZN(new_n873));
  OAI22_X1  g448(.A1(new_n512), .A2(new_n872), .B1(new_n514), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n865), .A2(new_n870), .A3(new_n871), .A4(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n543), .A2(G67), .A3(new_n544), .ZN(new_n877));
  INV_X1    g452(.A(new_n869), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n505), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI22_X1  g454(.A1(new_n559), .A2(new_n562), .B1(new_n879), .B2(new_n874), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n863), .B(new_n881), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n882), .A2(KEYINPUT39), .ZN(new_n883));
  INV_X1    g458(.A(G860), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(KEYINPUT39), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n879), .A2(new_n874), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n887), .A2(new_n884), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT37), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n886), .A2(new_n889), .ZN(G145));
  XNOR2_X1  g465(.A(new_n645), .B(G160), .ZN(new_n891));
  XNOR2_X1  g466(.A(G162), .B(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n484), .A2(G130), .ZN(new_n893));
  OAI21_X1  g468(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n894));
  INV_X1    g469(.A(G118), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n894), .B1(new_n895), .B2(G2105), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n896), .B1(new_n486), .B2(G142), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n494), .A2(new_n496), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(new_n491), .A3(new_n488), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n901), .B(new_n769), .C1(new_n770), .C2(new_n483), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n771), .A2(G164), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n794), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT107), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n794), .A2(new_n902), .A3(new_n903), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n907), .B1(new_n906), .B2(new_n908), .ZN(new_n911));
  OAI211_X1 g486(.A(KEYINPUT108), .B(new_n727), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n908), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n794), .B1(new_n902), .B2(new_n903), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n726), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n727), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT107), .B1(new_n913), .B2(new_n914), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n918), .B1(new_n919), .B2(new_n909), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n920), .A2(KEYINPUT108), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n899), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n920), .A2(KEYINPUT108), .B1(new_n726), .B2(new_n915), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n727), .B1(new_n910), .B2(new_n911), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(new_n898), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n826), .B(new_n649), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n922), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n928), .B1(new_n922), .B2(new_n927), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n892), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n928), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n917), .A2(new_n921), .A3(new_n899), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n898), .B1(new_n923), .B2(new_n926), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n892), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n922), .A2(new_n927), .A3(new_n928), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G37), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n931), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n940), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n942));
  NAND2_X1  g517(.A1(G290), .A2(G288), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n605), .A2(new_n588), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(G305), .B(G303), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n943), .A2(new_n942), .A3(new_n944), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n946), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n948), .B1(new_n950), .B2(new_n945), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT42), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n637), .B(new_n881), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT41), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n622), .A2(G299), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n616), .A2(new_n619), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT10), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n630), .B1(new_n960), .B2(new_n614), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n955), .B1(new_n956), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n622), .A2(G299), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n960), .A2(new_n630), .A3(new_n614), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(new_n964), .A3(KEYINPUT41), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n954), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n956), .A2(new_n961), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n967), .B1(new_n954), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n953), .A2(KEYINPUT110), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(KEYINPUT110), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n969), .A2(KEYINPUT110), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n971), .B1(new_n952), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(G868), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n887), .A2(G868), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(G295));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n979), .B1(new_n975), .B2(new_n977), .ZN(new_n980));
  AOI211_X1 g555(.A(KEYINPUT111), .B(new_n976), .C1(new_n974), .C2(G868), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(G331));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n983));
  OAI21_X1  g558(.A(G286), .B1(new_n549), .B2(new_n554), .ZN(new_n984));
  INV_X1    g559(.A(G64), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n522), .A2(new_n525), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(G651), .B1(new_n986), .B2(new_n547), .ZN(new_n987));
  AOI22_X1  g562(.A1(G52), .A2(new_n569), .B1(new_n550), .B2(new_n551), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(G168), .A3(new_n988), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n984), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n990), .A2(KEYINPUT112), .A3(new_n880), .A4(new_n876), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT112), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n984), .A2(new_n989), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n992), .B1(new_n881), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n881), .A2(new_n993), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n991), .A2(new_n994), .A3(new_n968), .A4(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n881), .A2(new_n993), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n880), .A2(new_n876), .B1(new_n984), .B2(new_n989), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n962), .B(new_n965), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  OR2_X1    g575(.A1(new_n951), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n991), .A2(new_n995), .A3(new_n994), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n1002), .A2(new_n962), .A3(new_n965), .ZN(new_n1003));
  NOR4_X1   g578(.A1(new_n997), .A2(new_n998), .A3(new_n961), .A4(new_n956), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n951), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1001), .A2(new_n939), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n983), .B1(new_n1006), .B2(KEYINPUT43), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1000), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n996), .A2(new_n999), .A3(KEYINPUT113), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(new_n951), .A3(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1011), .A2(KEYINPUT114), .A3(new_n939), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n1001), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT114), .B1(new_n1011), .B2(new_n939), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1007), .B1(new_n1015), .B2(KEYINPUT43), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT43), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1018));
  OR2_X1    g593(.A1(new_n1006), .A2(KEYINPUT43), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1017), .B1(new_n1020), .B2(new_n983), .ZN(new_n1021));
  AOI211_X1 g596(.A(KEYINPUT115), .B(KEYINPUT44), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1016), .B1(new_n1021), .B2(new_n1022), .ZN(G397));
  INV_X1    g598(.A(KEYINPUT45), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(G164), .B2(G1384), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G160), .A2(G40), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1028), .A2(G1996), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(KEYINPUT46), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n794), .B(G2067), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1028), .B1(new_n1031), .B2(new_n772), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g608(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1034));
  XNOR2_X1  g609(.A(new_n1033), .B(new_n1034), .ZN(new_n1035));
  XOR2_X1   g610(.A(new_n771), .B(G1996), .Z(new_n1036));
  AND2_X1   g611(.A1(new_n1031), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n828), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n826), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G2067), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n794), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1028), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n1043), .B(KEYINPUT125), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n826), .B(new_n828), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1037), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n605), .A2(new_n817), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1047), .B(KEYINPUT116), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n1027), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT48), .ZN(new_n1050));
  OAI22_X1  g625(.A1(new_n1046), .A2(new_n1028), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1051), .B1(new_n1050), .B2(new_n1049), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1035), .A2(new_n1044), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(G303), .A2(G8), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1054), .B(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1054), .B(KEYINPUT55), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT118), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT50), .ZN(new_n1061));
  INV_X1    g636(.A(G1384), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n901), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1026), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1063), .A2(new_n1064), .A3(new_n736), .A4(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n901), .A2(KEYINPUT45), .A3(new_n1062), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(new_n1025), .A3(new_n1065), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1066), .B1(new_n1069), .B2(G1971), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1058), .A2(new_n1060), .A3(new_n1070), .A4(G8), .ZN(new_n1071));
  INV_X1    g646(.A(G8), .ZN(new_n1072));
  NOR2_X1   g647(.A1(G164), .A2(G1384), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1072), .B1(new_n1073), .B2(new_n1065), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n588), .A2(G1976), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT52), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT49), .ZN(new_n1078));
  INV_X1    g653(.A(G1981), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n597), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n597), .A2(new_n1079), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1078), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1082), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(KEYINPUT49), .A3(new_n1080), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1083), .A2(new_n1085), .A3(new_n1074), .ZN(new_n1086));
  INV_X1    g661(.A(G1976), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT52), .B1(G288), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1088), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1077), .A2(new_n1086), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1074), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n588), .A2(new_n1087), .ZN(new_n1092));
  XOR2_X1   g667(.A(new_n1092), .B(KEYINPUT119), .Z(new_n1093));
  NAND2_X1  g668(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1081), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI22_X1  g670(.A1(new_n1071), .A2(new_n1090), .B1(new_n1091), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1090), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1071), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1070), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1059), .B1(new_n1099), .B2(new_n1072), .ZN(new_n1100));
  NAND2_X1  g675(.A1(KEYINPUT121), .A2(KEYINPUT63), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(G168), .B(G8), .C1(KEYINPUT121), .C2(KEYINPUT63), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n901), .A2(new_n1062), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1026), .B1(new_n1104), .B2(new_n1024), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1067), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1073), .A2(KEYINPUT120), .A3(KEYINPUT45), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1105), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n810), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1063), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G2084), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1103), .B1(new_n1110), .B2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1098), .A2(new_n1100), .A3(new_n1102), .A4(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1100), .A2(new_n1071), .A3(new_n1097), .A4(new_n1116), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n1101), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1096), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n630), .B(KEYINPUT57), .ZN(new_n1121));
  XOR2_X1   g696(.A(KEYINPUT56), .B(G2072), .Z(new_n1122));
  OAI221_X1 g697(.A(new_n1121), .B1(new_n1068), .B2(new_n1122), .C1(new_n1113), .C2(G1956), .ZN(new_n1123));
  INV_X1    g698(.A(G1348), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1104), .A2(new_n1026), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n1041), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1123), .A2(new_n633), .A3(new_n1128), .ZN(new_n1129));
  OAI22_X1  g704(.A1(new_n1113), .A2(G1956), .B1(new_n1068), .B2(new_n1122), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1121), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1132), .A2(KEYINPUT61), .A3(new_n1123), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1134), .B(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT60), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n633), .B1(new_n1128), .B2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1125), .A2(KEYINPUT60), .A3(new_n622), .A4(new_n1127), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1138), .A2(new_n1139), .B1(new_n1137), .B2(new_n1128), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT61), .B1(new_n1132), .B2(new_n1123), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT58), .B(G1341), .ZN(new_n1142));
  OAI22_X1  g717(.A1(new_n1068), .A2(G1996), .B1(new_n1126), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT59), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1143), .A2(new_n1144), .A3(new_n563), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1144), .B1(new_n1143), .B2(new_n563), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1140), .A2(new_n1141), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1133), .B1(new_n1136), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1110), .A2(G168), .A3(new_n1115), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(G8), .ZN(new_n1151));
  OR2_X1    g726(.A1(new_n1151), .A2(KEYINPUT51), .ZN(new_n1152));
  AOI21_X1  g727(.A(G168), .B1(new_n1110), .B2(new_n1115), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT51), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1100), .A2(new_n1071), .A3(new_n1097), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT53), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1068), .B2(G2078), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1157), .A2(G2078), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1105), .A2(new_n1107), .A3(new_n1108), .A4(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n759), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1158), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(G171), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1069), .A2(new_n1159), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1164), .A2(new_n1158), .A3(G301), .A4(new_n1161), .ZN(new_n1165));
  AOI21_X1  g740(.A(KEYINPUT54), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1156), .A2(new_n1166), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1162), .A2(G171), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n1164), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1168), .B(KEYINPUT54), .C1(new_n1169), .C2(G301), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1155), .A2(new_n1167), .A3(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1120), .B1(new_n1149), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT123), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT123), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1120), .B(new_n1174), .C1(new_n1149), .C2(new_n1171), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT124), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1155), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1176), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1155), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1156), .A2(new_n1163), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1173), .A2(new_n1175), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(G290), .A2(G1986), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(KEYINPUT117), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1048), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1046), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  AND2_X1   g763(.A1(new_n1188), .A2(new_n1027), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1053), .B1(new_n1184), .B2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g765(.A(G227), .ZN(new_n1192));
  INV_X1    g766(.A(new_n666), .ZN(new_n1193));
  INV_X1    g767(.A(new_n667), .ZN(new_n1194));
  AOI21_X1  g768(.A(new_n460), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g769(.A(G229), .ZN(new_n1196));
  NAND3_X1  g770(.A1(new_n1192), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g771(.A1(new_n1197), .A2(KEYINPUT127), .ZN(new_n1198));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n1199));
  NAND4_X1  g773(.A1(new_n1192), .A2(new_n1195), .A3(new_n1199), .A4(new_n1196), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  AND3_X1   g775(.A1(new_n1201), .A2(new_n940), .A3(new_n1020), .ZN(G308));
  NAND3_X1  g776(.A1(new_n1201), .A2(new_n940), .A3(new_n1020), .ZN(G225));
endmodule


