//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n548, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n561, new_n563, new_n564, new_n565, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1175, new_n1176;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT64), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT66), .Z(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G137), .ZN(new_n470));
  NAND2_X1  g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n467), .A2(new_n469), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n474), .A2(new_n461), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G124), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n478), .A2(KEYINPUT67), .A3(G124), .ZN(new_n484));
  AND4_X1   g059(.A1(new_n476), .A2(new_n481), .A3(new_n483), .A4(new_n484), .ZN(G162));
  NAND4_X1  g060(.A1(new_n467), .A2(new_n469), .A3(G126), .A4(G2105), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n487), .A2(new_n489), .A3(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n467), .A2(new_n469), .A3(G138), .A4(new_n461), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n462), .A2(KEYINPUT4), .A3(G138), .A4(new_n461), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n486), .A2(KEYINPUT68), .A3(new_n490), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n493), .A2(new_n496), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(KEYINPUT69), .A3(G543), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n503), .A2(new_n505), .B1(KEYINPUT5), .B2(new_n502), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT6), .B(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n509), .A2(G88), .B1(G50), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n503), .A2(new_n505), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n502), .A2(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n522), .A2(KEYINPUT70), .A3(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n512), .A2(new_n516), .A3(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(G166));
  NAND2_X1  g100(.A1(new_n509), .A2(G89), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n511), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n530));
  AND3_X1   g105(.A1(new_n529), .A2(KEYINPUT71), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(KEYINPUT71), .B1(new_n529), .B2(new_n530), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n526), .B(new_n528), .C1(new_n531), .C2(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  AOI22_X1  g109(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n515), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n508), .A2(new_n537), .B1(new_n538), .B2(new_n510), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  AOI22_X1  g115(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n515), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT72), .B(G81), .ZN(new_n543));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n508), .A2(new_n543), .B1(new_n544), .B2(new_n510), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(G188));
  AOI22_X1  g127(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(KEYINPUT73), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(KEYINPUT73), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n554), .A2(G651), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n509), .A2(G91), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n511), .A2(G53), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT9), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(G299));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n561));
  XNOR2_X1  g136(.A(G171), .B(new_n561), .ZN(G301));
  NAND2_X1  g137(.A1(new_n524), .A2(KEYINPUT75), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n512), .A2(new_n516), .A3(new_n523), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(G303));
  NAND2_X1  g141(.A1(new_n509), .A2(G87), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n511), .A2(G49), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(G288));
  NAND3_X1  g145(.A1(new_n506), .A2(G86), .A3(new_n507), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n507), .A2(G48), .A3(G543), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n504), .A2(KEYINPUT69), .A3(G543), .ZN(new_n574));
  AOI21_X1  g149(.A(KEYINPUT69), .B1(new_n504), .B2(G543), .ZN(new_n575));
  OAI211_X1 g150(.A(G61), .B(new_n519), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n518), .A2(KEYINPUT76), .A3(G61), .A4(new_n519), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n573), .B1(new_n581), .B2(G651), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n509), .A2(G85), .B1(G47), .B2(new_n511), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT78), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n584), .B(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n515), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT77), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n586), .A2(new_n589), .ZN(G290));
  INV_X1    g165(.A(G92), .ZN(new_n591));
  OR3_X1    g166(.A1(new_n508), .A2(KEYINPUT10), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(KEYINPUT10), .B1(new_n508), .B2(new_n591), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n511), .A2(G54), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(new_n515), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g176(.A(G171), .B(KEYINPUT74), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(KEYINPUT79), .Z(G284));
  XNOR2_X1  g179(.A(new_n603), .B(KEYINPUT80), .ZN(G321));
  NAND2_X1  g180(.A1(G286), .A2(G868), .ZN(new_n606));
  INV_X1    g181(.A(G299), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(G297));
  OAI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(G280));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n598), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n598), .A2(new_n610), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OR3_X1    g188(.A1(new_n613), .A2(KEYINPUT81), .A3(new_n600), .ZN(new_n614));
  OAI21_X1  g189(.A(KEYINPUT81), .B1(new_n613), .B2(new_n600), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n614), .B(new_n615), .C1(G868), .C2(new_n546), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n475), .A2(G2104), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT12), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2100), .Z(new_n621));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n622));
  INV_X1    g197(.A(G123), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n479), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n475), .A2(G135), .ZN(new_n625));
  OR2_X1    g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n626), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n478), .A2(KEYINPUT82), .A3(G123), .ZN(new_n628));
  NAND4_X1  g203(.A1(new_n624), .A2(new_n625), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n621), .A2(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2435), .ZN(new_n633));
  XOR2_X1   g208(.A(G2427), .B(G2438), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(KEYINPUT14), .ZN(new_n636));
  XOR2_X1   g211(.A(G2451), .B(G2454), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n636), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G1341), .B(G1348), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(G14), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n643), .A2(new_n644), .ZN(G401));
  XNOR2_X1  g220(.A(G2084), .B(G2090), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT83), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2072), .B(G2078), .ZN(new_n648));
  XOR2_X1   g223(.A(G2067), .B(G2678), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n647), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT84), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n648), .B(KEYINPUT17), .Z(new_n653));
  OAI21_X1  g228(.A(new_n652), .B1(new_n653), .B2(new_n649), .ZN(new_n654));
  INV_X1    g229(.A(new_n647), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n655), .A2(new_n648), .A3(new_n650), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT18), .Z(new_n657));
  NAND3_X1  g232(.A1(new_n655), .A2(new_n653), .A3(new_n649), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n654), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT85), .B(G2096), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2100), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n659), .B(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n665), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n670), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n667), .A2(new_n669), .A3(new_n671), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n674), .B(new_n675), .C1(new_n673), .C2(new_n672), .ZN(new_n676));
  XOR2_X1   g251(.A(G1991), .B(G1996), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT86), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n680), .B(new_n682), .Z(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G229));
  INV_X1    g259(.A(KEYINPUT23), .ZN(new_n685));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G20), .ZN(new_n687));
  AOI22_X1  g262(.A1(G299), .A2(G16), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(new_n685), .B2(new_n687), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1956), .ZN(new_n690));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n691), .A2(G33), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT93), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT25), .ZN(new_n695));
  NAND2_X1  g270(.A1(G115), .A2(G2104), .ZN(new_n696));
  INV_X1    g271(.A(G127), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n474), .B2(new_n697), .ZN(new_n698));
  AOI22_X1  g273(.A1(new_n698), .A2(G2105), .B1(new_n475), .B2(G139), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n692), .B1(new_n700), .B2(G29), .ZN(new_n701));
  INV_X1    g276(.A(G2072), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT94), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n701), .A2(new_n702), .ZN(new_n706));
  OAI21_X1  g281(.A(G29), .B1(new_n465), .B2(new_n472), .ZN(new_n707));
  INV_X1    g282(.A(G2084), .ZN(new_n708));
  INV_X1    g283(.A(G34), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n709), .A2(KEYINPUT24), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(KEYINPUT24), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n691), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n707), .A2(new_n708), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n706), .B1(KEYINPUT100), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(KEYINPUT100), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT30), .B(G28), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n715), .B1(new_n691), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n705), .A2(new_n714), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(G168), .A2(KEYINPUT97), .A3(G16), .ZN(new_n720));
  OAI21_X1  g295(.A(KEYINPUT97), .B1(G16), .B2(G21), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G286), .B2(new_n686), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n720), .A2(G1966), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n720), .A2(new_n722), .ZN(new_n724));
  INV_X1    g299(.A(G1966), .ZN(new_n725));
  AOI21_X1  g300(.A(KEYINPUT98), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AND3_X1   g301(.A1(new_n724), .A2(KEYINPUT98), .A3(new_n725), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n719), .B(new_n723), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n708), .B1(new_n707), .B2(new_n712), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n691), .A2(G27), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G164), .B2(new_n691), .ZN(new_n732));
  MUX2_X1   g307(.A(new_n731), .B(new_n732), .S(KEYINPUT101), .Z(new_n733));
  INV_X1    g308(.A(G2078), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n629), .A2(new_n691), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT99), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G5), .B2(G16), .ZN(new_n738));
  OR3_X1    g313(.A1(new_n737), .A2(G5), .A3(G16), .ZN(new_n739));
  INV_X1    g314(.A(G171), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n738), .B(new_n739), .C1(new_n740), .C2(new_n686), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G1961), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n478), .A2(G129), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT95), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n475), .A2(G141), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT26), .Z(new_n748));
  NAND4_X1  g323(.A1(new_n743), .A2(new_n745), .A3(new_n746), .A4(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n749), .A2(new_n691), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(KEYINPUT96), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT96), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G29), .B2(G32), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n751), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT27), .B(G1996), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT31), .B(G11), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n742), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n730), .A2(new_n735), .A3(new_n736), .A4(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT102), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n690), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(G25), .A2(G29), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n478), .A2(G119), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT87), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n475), .A2(G131), .ZN(new_n766));
  NOR2_X1   g341(.A1(G95), .A2(G2105), .ZN(new_n767));
  OAI21_X1  g342(.A(G2104), .B1(new_n461), .B2(G107), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT88), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n763), .B1(new_n771), .B2(G29), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT35), .B(G1991), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  MUX2_X1   g349(.A(G24), .B(G290), .S(G16), .Z(new_n775));
  NOR2_X1   g350(.A1(new_n775), .A2(G1986), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n775), .A2(G1986), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n774), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n686), .A2(G22), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G166), .B2(new_n686), .ZN(new_n780));
  INV_X1    g355(.A(G1971), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G16), .A2(G23), .ZN(new_n783));
  INV_X1    g358(.A(G288), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT33), .B(G1976), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n686), .A2(G6), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n582), .B2(new_n686), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT32), .B(G1981), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n782), .A2(new_n787), .A3(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT34), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n778), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT36), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n728), .A2(new_n758), .A3(new_n729), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n797), .A2(KEYINPUT102), .A3(new_n735), .A4(new_n736), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n691), .A2(G35), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G162), .B2(new_n691), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT29), .B(G2090), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n762), .A2(new_n796), .A3(new_n798), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n691), .A2(G26), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n478), .A2(G128), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT90), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n475), .A2(G140), .ZN(new_n808));
  OAI21_X1  g383(.A(G2104), .B1(new_n461), .B2(G116), .ZN(new_n809));
  NOR2_X1   g384(.A1(G104), .A2(G2105), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT91), .Z(new_n811));
  OAI21_X1  g386(.A(new_n808), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n807), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n804), .B1(new_n813), .B2(new_n691), .ZN(new_n814));
  MUX2_X1   g389(.A(new_n804), .B(new_n814), .S(KEYINPUT28), .Z(new_n815));
  XOR2_X1   g390(.A(KEYINPUT92), .B(G2067), .Z(new_n816));
  XOR2_X1   g391(.A(new_n815), .B(new_n816), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n686), .A2(G4), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n598), .B2(new_n686), .ZN(new_n819));
  INV_X1    g394(.A(G1348), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n686), .A2(G19), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n546), .B2(new_n686), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT89), .Z(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(G1341), .Z(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NOR4_X1   g402(.A1(new_n803), .A2(new_n817), .A3(new_n822), .A4(new_n827), .ZN(G311));
  INV_X1    g403(.A(new_n803), .ZN(new_n829));
  INV_X1    g404(.A(new_n817), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n829), .A2(new_n830), .A3(new_n821), .A4(new_n826), .ZN(G150));
  NAND2_X1  g406(.A1(new_n598), .A2(G559), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT39), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n832), .B(new_n834), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n836), .A2(new_n515), .ZN(new_n837));
  INV_X1    g412(.A(G93), .ZN(new_n838));
  INV_X1    g413(.A(G55), .ZN(new_n839));
  OAI22_X1  g414(.A1(new_n508), .A2(new_n838), .B1(new_n839), .B2(new_n510), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n546), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n835), .B(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n843), .A2(G860), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT104), .Z(new_n845));
  OAI21_X1  g420(.A(G860), .B1(new_n837), .B2(new_n840), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT37), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(G145));
  XNOR2_X1  g423(.A(new_n629), .B(G160), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G162), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n478), .A2(G130), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n475), .A2(G142), .ZN(new_n853));
  NOR2_X1   g428(.A1(G106), .A2(G2105), .ZN(new_n854));
  OAI21_X1  g429(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n852), .B(new_n853), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n770), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT106), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n619), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n496), .A2(new_n497), .A3(new_n486), .A4(new_n490), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n749), .B(new_n861), .Z(new_n862));
  NOR2_X1   g437(.A1(new_n700), .A2(KEYINPUT105), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n813), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT107), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n851), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n859), .A2(new_n619), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n859), .A2(new_n619), .ZN(new_n870));
  OR3_X1    g445(.A1(new_n869), .A2(new_n870), .A3(new_n865), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n860), .A2(new_n865), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(new_n872), .A3(KEYINPUT107), .ZN(new_n873));
  AOI21_X1  g448(.A(G37), .B1(new_n868), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n871), .A2(new_n872), .A3(new_n851), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g452(.A1(G299), .A2(KEYINPUT108), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT108), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n556), .A2(new_n880), .A3(new_n557), .A4(new_n559), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n598), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n879), .A2(new_n882), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n885), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT41), .B1(new_n887), .B2(new_n883), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n884), .A2(new_n885), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT109), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n886), .A2(KEYINPUT109), .A3(KEYINPUT41), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n613), .B(new_n842), .ZN(new_n895));
  MUX2_X1   g470(.A(new_n886), .B(new_n894), .S(new_n895), .Z(new_n896));
  XOR2_X1   g471(.A(G290), .B(KEYINPUT110), .Z(new_n897));
  XNOR2_X1  g472(.A(new_n582), .B(G288), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(G166), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n897), .B(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT42), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n896), .A2(new_n901), .ZN(new_n903));
  OAI21_X1  g478(.A(G868), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(G868), .B2(new_n841), .ZN(G295));
  OAI21_X1  g480(.A(new_n904), .B1(G868), .B2(new_n841), .ZN(G331));
  INV_X1    g481(.A(new_n842), .ZN(new_n907));
  NAND2_X1  g482(.A1(G301), .A2(G168), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT111), .ZN(new_n909));
  NAND2_X1  g484(.A1(G286), .A2(G171), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n909), .B1(new_n908), .B2(new_n910), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n907), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT112), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n602), .A2(G286), .ZN(new_n915));
  INV_X1    g490(.A(new_n910), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT111), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n842), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n913), .A2(new_n914), .A3(new_n919), .ZN(new_n920));
  OAI211_X1 g495(.A(KEYINPUT112), .B(new_n907), .C1(new_n911), .C2(new_n912), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n892), .A2(new_n920), .A3(new_n893), .A4(new_n921), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n913), .A2(new_n885), .A3(new_n919), .A4(new_n884), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n900), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(G37), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n900), .B1(new_n922), .B2(new_n923), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT43), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n900), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n886), .B1(new_n920), .B2(new_n921), .ZN(new_n930));
  AOI22_X1  g505(.A1(new_n888), .A2(new_n890), .B1(new_n913), .B2(new_n919), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n932), .A2(new_n924), .A3(new_n933), .A4(new_n925), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n928), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n933), .B1(new_n926), .B2(new_n927), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n932), .A2(new_n924), .A3(KEYINPUT43), .A4(new_n925), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  MUX2_X1   g513(.A(new_n935), .B(new_n938), .S(KEYINPUT44), .Z(G397));
  OAI21_X1  g514(.A(KEYINPUT113), .B1(G290), .B2(G1986), .ZN(new_n940));
  NAND2_X1  g515(.A1(G290), .A2(G1986), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n940), .B(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G1384), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n861), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT45), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(G160), .A2(G40), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n942), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n813), .B(G2067), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n749), .A2(G1996), .ZN(new_n951));
  INV_X1    g526(.A(new_n749), .ZN(new_n952));
  INV_X1    g527(.A(G1996), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n950), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n770), .B(new_n773), .Z(new_n956));
  OAI21_X1  g531(.A(new_n948), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n949), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(G305), .A2(G1981), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT117), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n581), .A2(G651), .ZN(new_n961));
  INV_X1    g536(.A(G1981), .ZN(new_n962));
  INV_X1    g537(.A(new_n573), .ZN(new_n963));
  AND4_X1   g538(.A1(new_n960), .A2(new_n961), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n960), .B1(new_n582), .B2(new_n962), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n959), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT49), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n947), .A2(new_n944), .ZN(new_n969));
  INV_X1    g544(.A(G8), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI211_X1 g546(.A(KEYINPUT49), .B(new_n959), .C1(new_n964), .C2(new_n965), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n968), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1976), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(new_n974), .A3(new_n784), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n964), .A2(new_n965), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n971), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n499), .A2(new_n943), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n979), .A2(KEYINPUT114), .A3(new_n945), .ZN(new_n980));
  INV_X1    g555(.A(G40), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n465), .A2(new_n981), .A3(new_n472), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n861), .A2(KEYINPUT45), .A3(new_n943), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT45), .B1(new_n499), .B2(new_n943), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n984), .B1(new_n985), .B2(KEYINPUT114), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n781), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT115), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n499), .B2(new_n943), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n496), .A2(new_n497), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n989), .B(new_n943), .C1(new_n991), .C2(new_n491), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n982), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G2090), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT116), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n997));
  NOR4_X1   g572(.A1(new_n990), .A2(new_n993), .A3(new_n997), .A4(G2090), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n947), .B1(new_n985), .B2(KEYINPUT114), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n486), .A2(KEYINPUT68), .A3(new_n490), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT68), .B1(new_n486), .B2(new_n490), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n991), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1384), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1001), .B1(new_n1006), .B2(KEYINPUT45), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1000), .A2(new_n1007), .A3(new_n984), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(new_n1009), .A3(new_n781), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n988), .A2(new_n999), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(G303), .B2(G8), .ZN(new_n1013));
  AOI211_X1 g588(.A(KEYINPUT55), .B(new_n970), .C1(new_n563), .C2(new_n565), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1011), .A2(new_n1015), .A3(G8), .ZN(new_n1016));
  INV_X1    g591(.A(new_n971), .ZN(new_n1017));
  NOR2_X1   g592(.A1(G288), .A2(new_n974), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT52), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT52), .B1(G288), .B2(new_n974), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n971), .B(new_n1020), .C1(new_n974), .C2(G288), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n973), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1016), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n978), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1011), .A2(new_n1015), .A3(G8), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n973), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1017), .B1(new_n975), .B2(new_n976), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT118), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1025), .A2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n946), .B(new_n982), .C1(new_n979), .C2(new_n945), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n725), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n994), .A2(new_n708), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(G168), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n970), .A2(KEYINPUT122), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1036), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1039));
  AOI211_X1 g614(.A(new_n970), .B(G168), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1000), .A2(new_n734), .A3(new_n1007), .A4(new_n984), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n994), .A2(G1961), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n734), .A2(KEYINPUT53), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1032), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  AND4_X1   g624(.A1(G301), .A2(new_n1044), .A3(new_n1046), .A4(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1045), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n982), .A2(KEYINPUT123), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1047), .B1(new_n982), .B2(KEYINPUT123), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1052), .A2(new_n1053), .A3(new_n946), .A4(new_n984), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n740), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT54), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1051), .A2(G301), .A3(new_n1054), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n1058));
  AOI211_X1 g633(.A(new_n1045), .B(new_n1048), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1057), .B(new_n1058), .C1(new_n1059), .C2(G301), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1041), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n979), .A2(KEYINPUT50), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n992), .A2(new_n982), .ZN(new_n1063));
  AOI21_X1  g638(.A(G1348), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT60), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n982), .A2(new_n943), .A3(new_n861), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(G2067), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1065), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT121), .B1(new_n1070), .B2(new_n598), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n820), .B1(new_n990), .B2(new_n993), .ZN(new_n1072));
  INV_X1    g647(.A(G2067), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n969), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT60), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n1076));
  NOR3_X1   g651(.A1(new_n1075), .A2(new_n1076), .A3(new_n599), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1069), .B1(new_n1071), .B2(new_n1077), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT58), .B(G1341), .Z(new_n1079));
  NAND2_X1  g654(.A1(new_n1066), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1008), .B2(G1996), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1081), .A2(KEYINPUT120), .A3(KEYINPUT59), .A4(new_n546), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1070), .A2(KEYINPUT121), .A3(new_n598), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1076), .B1(new_n1075), .B2(new_n599), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1083), .A2(new_n1068), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n983), .A2(new_n986), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1087), .A2(new_n953), .B1(new_n1066), .B2(new_n1079), .ZN(new_n1088));
  INV_X1    g663(.A(new_n546), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1086), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1078), .A2(new_n1082), .A3(new_n1085), .A4(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n607), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n944), .A2(KEYINPUT50), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n982), .B(new_n1096), .C1(new_n979), .C2(KEYINPUT50), .ZN(new_n1097));
  INV_X1    g672(.A(G1956), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1087), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1095), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1101), .A2(new_n1099), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1104), .A2(new_n599), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1102), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1091), .A2(new_n1106), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1097), .A2(G2090), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(new_n1008), .B2(new_n781), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1108), .B1(new_n970), .B2(new_n1110), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1022), .A2(new_n1026), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT61), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1102), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1095), .A2(KEYINPUT61), .A3(new_n1099), .A4(new_n1101), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1106), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1061), .A2(new_n1107), .A3(new_n1112), .A4(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n1041), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1041), .A2(new_n1118), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1059), .A2(G301), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1119), .A2(new_n1112), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1031), .A2(new_n1117), .A3(new_n1122), .ZN(new_n1123));
  AOI211_X1 g698(.A(new_n970), .B(G286), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1112), .A2(KEYINPUT119), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT63), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1022), .A2(new_n1026), .A3(new_n1111), .A4(new_n1124), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1125), .A2(new_n1126), .A3(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1016), .A2(new_n1027), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1011), .A2(G8), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1126), .B1(new_n1132), .B2(new_n1108), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1131), .A2(new_n1124), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1130), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n958), .B1(new_n1123), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n950), .A2(new_n952), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1137), .A2(new_n948), .B1(KEYINPUT125), .B2(KEYINPUT46), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n948), .A2(new_n953), .ZN(new_n1139));
  NOR2_X1   g714(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n1139), .B(new_n1140), .Z(new_n1141));
  NAND2_X1  g716(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT47), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1142), .B(new_n1143), .ZN(new_n1144));
  NOR4_X1   g719(.A1(G290), .A2(G1986), .A3(new_n946), .A4(new_n947), .ZN(new_n1145));
  OR2_X1    g720(.A1(new_n1145), .A2(KEYINPUT48), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(KEYINPUT48), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1146), .A2(new_n957), .A3(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1144), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n773), .B1(new_n955), .B2(new_n948), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n771), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n813), .A2(new_n1073), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT124), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT124), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1151), .A2(new_n1155), .A3(new_n1152), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1154), .A2(new_n948), .A3(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1149), .A2(new_n1157), .A3(KEYINPUT126), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT126), .B1(new_n1149), .B2(new_n1157), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT127), .B1(new_n1136), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n958), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1134), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1127), .B(KEYINPUT119), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1164), .B1(new_n1165), .B2(new_n1126), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1031), .A2(new_n1117), .A3(new_n1122), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1163), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1160), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n1158), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1168), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1162), .A2(new_n1172), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g748(.A(new_n662), .B1(new_n643), .B2(new_n644), .ZN(new_n1175));
  AOI21_X1  g749(.A(new_n1175), .B1(new_n874), .B2(new_n875), .ZN(new_n1176));
  NAND4_X1  g750(.A1(new_n935), .A2(new_n1176), .A3(G319), .A4(new_n683), .ZN(G225));
  INV_X1    g751(.A(G225), .ZN(G308));
endmodule


