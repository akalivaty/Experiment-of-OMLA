//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n547, new_n549, new_n550, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n564, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n602, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT66), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT67), .Z(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n460), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  OR2_X1    g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(G137), .ZN(new_n464));
  NAND2_X1  g039(.A1(G101), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(new_n462), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(G160));
  OR2_X1    g044(.A1(G100), .A2(G2105), .ZN(new_n470));
  OAI211_X1 g045(.A(new_n470), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n471));
  AND3_X1   g046(.A1(new_n460), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n472));
  AOI21_X1  g047(.A(KEYINPUT69), .B1(new_n460), .B2(G2105), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G124), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n460), .A2(new_n462), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n476), .B(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G136), .ZN(new_n479));
  OAI221_X1 g054(.A(new_n471), .B1(new_n474), .B2(new_n475), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n480), .B(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  NAND3_X1  g058(.A1(new_n460), .A2(KEYINPUT4), .A3(G138), .ZN(new_n484));
  NAND2_X1  g059(.A1(G102), .A2(G2104), .ZN(new_n485));
  AOI21_X1  g060(.A(G2105), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(G114), .A2(G2104), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n460), .B2(G126), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT4), .B1(new_n489), .B2(new_n462), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n460), .A2(G138), .A3(new_n462), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n486), .B1(new_n490), .B2(new_n491), .ZN(G164));
  INV_X1    g067(.A(G651), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT6), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G543), .ZN(new_n495));
  AND2_X1   g070(.A1(KEYINPUT71), .A2(KEYINPUT6), .ZN(new_n496));
  NOR2_X1   g071(.A1(KEYINPUT71), .A2(KEYINPUT6), .ZN(new_n497));
  OAI21_X1  g072(.A(G651), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT72), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT72), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(G651), .C1(new_n496), .C2(new_n497), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n495), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G50), .ZN(new_n503));
  NAND2_X1  g078(.A1(G75), .A2(G543), .ZN(new_n504));
  XNOR2_X1  g079(.A(new_n504), .B(KEYINPUT74), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  AND3_X1   g084(.A1(new_n507), .A2(new_n509), .A3(G62), .ZN(new_n510));
  OAI21_X1  g085(.A(G651), .B1(new_n505), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT75), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n511), .B(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n507), .A2(new_n509), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT71), .B(KEYINPUT6), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n500), .B1(new_n516), .B2(G651), .ZN(new_n517));
  INV_X1    g092(.A(new_n501), .ZN(new_n518));
  OAI211_X1 g093(.A(new_n515), .B(new_n494), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n499), .A2(new_n501), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n522), .A2(KEYINPUT73), .A3(new_n515), .A4(new_n494), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  OAI211_X1 g100(.A(new_n503), .B(new_n513), .C1(new_n524), .C2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND3_X1  g102(.A1(new_n521), .A2(G89), .A3(new_n523), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n502), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n528), .A2(new_n529), .A3(new_n531), .A4(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  INV_X1    g109(.A(new_n524), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G90), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(new_n493), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n502), .A2(G52), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(G171));
  NAND3_X1  g115(.A1(new_n521), .A2(G81), .A3(new_n523), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n493), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n502), .A2(G43), .ZN(new_n544));
  AND3_X1   g119(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(G188));
  NAND2_X1  g126(.A1(new_n515), .A2(G65), .ZN(new_n552));
  NAND2_X1  g127(.A1(G78), .A2(G543), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n493), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n495), .ZN(new_n555));
  OAI211_X1 g130(.A(G53), .B(new_n555), .C1(new_n517), .C2(new_n518), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT9), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n502), .A2(new_n558), .A3(G53), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n554), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n521), .A2(G91), .A3(new_n523), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(G299));
  NAND3_X1  g137(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(G301));
  NAND3_X1  g138(.A1(new_n521), .A2(G87), .A3(new_n523), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n502), .A2(G49), .ZN(new_n566));
  AND3_X1   g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G288));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n569));
  AND3_X1   g144(.A1(new_n502), .A2(new_n569), .A3(G48), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n569), .B1(new_n502), .B2(G48), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n573), .A2(new_n493), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n521), .A2(G86), .A3(new_n523), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(G305));
  AOI22_X1  g151(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  XOR2_X1   g152(.A(new_n577), .B(KEYINPUT77), .Z(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(G651), .B1(G47), .B2(new_n502), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n535), .A2(G85), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(G290));
  NAND2_X1  g156(.A1(G301), .A2(G868), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT10), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n535), .A2(new_n583), .A3(G92), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n515), .A2(G66), .ZN(new_n585));
  NAND2_X1  g160(.A1(G79), .A2(G543), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT78), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n493), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(G54), .B2(new_n502), .ZN(new_n589));
  INV_X1    g164(.A(G92), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT10), .B1(new_n524), .B2(new_n590), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n584), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n582), .B1(new_n592), .B2(G868), .ZN(G284));
  XNOR2_X1  g168(.A(G284), .B(KEYINPUT79), .ZN(G321));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NOR2_X1   g170(.A1(G168), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(KEYINPUT80), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(G299), .B2(new_n595), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n597), .B1(new_n596), .B2(new_n599), .ZN(G297));
  OAI21_X1  g175(.A(new_n597), .B1(new_n596), .B2(new_n599), .ZN(G280));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n592), .B1(new_n602), .B2(G860), .ZN(G148));
  NAND2_X1  g178(.A1(new_n592), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g182(.A1(G99), .A2(G2105), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n608), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n609));
  INV_X1    g184(.A(G123), .ZN(new_n610));
  INV_X1    g185(.A(G135), .ZN(new_n611));
  OAI221_X1 g186(.A(new_n609), .B1(new_n474), .B2(new_n610), .C1(new_n478), .C2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT82), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(G2096), .Z(new_n617));
  INV_X1    g192(.A(G2104), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n476), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT12), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XOR2_X1   g196(.A(KEYINPUT81), .B(G2100), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n617), .A2(new_n623), .ZN(G156));
  XNOR2_X1  g199(.A(G2443), .B(G2446), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT15), .B(G2435), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2438), .ZN(new_n628));
  XOR2_X1   g203(.A(G2427), .B(G2430), .Z(new_n629));
  OAI21_X1  g204(.A(KEYINPUT14), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT83), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n628), .A2(new_n629), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n633), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n636), .A2(new_n638), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n626), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n643), .A2(new_n625), .A3(new_n639), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n642), .A2(new_n644), .A3(G14), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(G401));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2072), .B(G2078), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT84), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT18), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n648), .B(KEYINPUT85), .Z(new_n653));
  OAI21_X1  g228(.A(KEYINPUT17), .B1(new_n653), .B2(new_n647), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(new_n649), .Z(new_n655));
  AND2_X1   g230(.A1(new_n653), .A2(new_n647), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n652), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT86), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2096), .B(G2100), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(G227));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT87), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1956), .B(G2474), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G1971), .B(G1976), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT89), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n666), .A2(new_n662), .A3(new_n663), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT90), .Z(new_n672));
  NAND2_X1  g247(.A1(new_n662), .A2(new_n663), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n664), .A2(new_n666), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  INV_X1    g252(.A(G1981), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n676), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT91), .B(G1986), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n682), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G229));
  NAND2_X1  g261(.A1(new_n592), .A2(G16), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G4), .B2(G16), .ZN(new_n688));
  INV_X1    g263(.A(G1348), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(G168), .A2(G16), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G16), .B2(G21), .ZN(new_n692));
  INV_X1    g267(.A(G1966), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G19), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(new_n545), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G1341), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n690), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n616), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT28), .ZN(new_n702));
  INV_X1    g277(.A(G26), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(G29), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(G29), .ZN(new_n705));
  OR2_X1    g280(.A1(G104), .A2(G2105), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n706), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT96), .ZN(new_n708));
  INV_X1    g283(.A(G128), .ZN(new_n709));
  INV_X1    g284(.A(G140), .ZN(new_n710));
  OAI221_X1 g285(.A(new_n708), .B1(new_n474), .B2(new_n709), .C1(new_n478), .C2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n705), .B1(new_n711), .B2(G29), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n704), .B1(new_n712), .B2(new_n702), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n701), .A2(G29), .B1(new_n713), .B2(G2067), .ZN(new_n714));
  NAND2_X1  g289(.A1(G171), .A2(G16), .ZN(new_n715));
  OR2_X1    g290(.A1(G5), .A2(G16), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT98), .B(G1961), .Z(new_n717));
  AND3_X1   g292(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n717), .B1(new_n715), .B2(new_n716), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT31), .B(G11), .Z(new_n720));
  NOR3_X1   g295(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n713), .A2(G2067), .ZN(new_n722));
  OR2_X1    g297(.A1(G29), .A2(G32), .ZN(new_n723));
  INV_X1    g298(.A(new_n478), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G141), .ZN(new_n725));
  INV_X1    g300(.A(new_n474), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G129), .ZN(new_n727));
  NAND3_X1  g302(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT26), .Z(new_n729));
  NAND3_X1  g304(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n725), .A2(new_n727), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n723), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT27), .B(G1996), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n722), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n732), .A2(G27), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G164), .B2(new_n732), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT99), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G2078), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT25), .Z(new_n743));
  AOI22_X1  g318(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n744));
  INV_X1    g319(.A(G139), .ZN(new_n745));
  OAI221_X1 g320(.A(new_n743), .B1(new_n462), .B2(new_n744), .C1(new_n478), .C2(new_n745), .ZN(new_n746));
  MUX2_X1   g321(.A(G33), .B(new_n746), .S(G29), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G2072), .ZN(new_n748));
  NOR3_X1   g323(.A1(new_n737), .A2(new_n741), .A3(new_n748), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n700), .A2(new_n714), .A3(new_n721), .A4(new_n749), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n732), .A2(G35), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n482), .B2(G29), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT29), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G2090), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT100), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n754), .A2(G2090), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT30), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(G28), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(G28), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n759), .A2(new_n760), .A3(new_n732), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT24), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(G34), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(G34), .ZN(new_n764));
  AOI21_X1  g339(.A(G29), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n468), .B2(G29), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G2084), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n757), .A2(new_n761), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n688), .A2(new_n689), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  NOR4_X1   g345(.A1(new_n750), .A2(new_n756), .A3(new_n768), .A4(new_n770), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n692), .A2(new_n693), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT97), .Z(new_n773));
  NAND2_X1  g348(.A1(G299), .A2(G16), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n695), .A2(KEYINPUT23), .A3(G20), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT23), .ZN(new_n776));
  INV_X1    g351(.A(G20), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(G16), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n774), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1956), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n697), .A2(G1341), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n771), .A2(new_n773), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT94), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(KEYINPUT36), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT95), .ZN(new_n787));
  NOR2_X1   g362(.A1(G16), .A2(G23), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n567), .B2(G16), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT33), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1976), .ZN(new_n791));
  MUX2_X1   g366(.A(G6), .B(G305), .S(G16), .Z(new_n792));
  XOR2_X1   g367(.A(KEYINPUT32), .B(G1981), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G16), .A2(G22), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G166), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT93), .B(G1971), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n791), .A2(new_n794), .A3(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT34), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n695), .A2(G24), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G290), .B2(G16), .ZN(new_n805));
  INV_X1    g380(.A(G1986), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n732), .A2(G25), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n724), .A2(G131), .B1(new_n726), .B2(G119), .ZN(new_n809));
  OR2_X1    g384(.A1(G95), .A2(G2105), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n810), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n808), .B1(new_n813), .B2(new_n732), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT35), .B(G1991), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT92), .Z(new_n816));
  OR2_X1    g391(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n805), .A2(new_n806), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n814), .A2(new_n816), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n807), .A2(new_n817), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n787), .B1(new_n803), .B2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n787), .ZN(new_n823));
  AOI211_X1 g398(.A(new_n820), .B(new_n823), .C1(new_n801), .C2(new_n802), .ZN(new_n824));
  NOR3_X1   g399(.A1(new_n784), .A2(new_n822), .A3(new_n824), .ZN(G311));
  NOR3_X1   g400(.A1(new_n750), .A2(new_n768), .A3(new_n770), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n755), .B(KEYINPUT100), .Z(new_n827));
  AND4_X1   g402(.A1(new_n781), .A2(new_n826), .A3(new_n783), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n803), .A2(new_n821), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(new_n823), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n803), .A2(new_n821), .A3(new_n787), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n828), .A2(new_n830), .A3(new_n773), .A4(new_n831), .ZN(G150));
  NAND2_X1  g407(.A1(G80), .A2(G543), .ZN(new_n833));
  INV_X1    g408(.A(G67), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n514), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G651), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT101), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n502), .A2(G55), .ZN(new_n838));
  INV_X1    g413(.A(G93), .ZN(new_n839));
  OAI211_X1 g414(.A(new_n837), .B(new_n838), .C1(new_n839), .C2(new_n524), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n545), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n545), .A2(new_n840), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT38), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n592), .A2(G559), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT102), .ZN(new_n848));
  AOI21_X1  g423(.A(G860), .B1(new_n846), .B2(KEYINPUT39), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n840), .A2(G860), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT37), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(G145));
  XNOR2_X1  g428(.A(new_n711), .B(new_n620), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n468), .A3(new_n615), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n468), .B1(new_n614), .B2(new_n615), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n482), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n858), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n860), .A2(G162), .A3(new_n856), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n746), .B(G164), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n859), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n862), .B1(new_n859), .B2(new_n861), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n724), .A2(G142), .B1(new_n726), .B2(G130), .ZN(new_n866));
  NOR2_X1   g441(.A1(G106), .A2(G2105), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n812), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n731), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n864), .A2(new_n865), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n731), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n870), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n859), .A2(new_n861), .ZN(new_n875));
  INV_X1    g450(.A(new_n862), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n874), .B1(new_n877), .B2(new_n863), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n855), .B1(new_n872), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n871), .B1(new_n864), .B2(new_n865), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n877), .A2(new_n874), .A3(new_n863), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(new_n854), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n879), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n567), .A2(G305), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n567), .A2(G305), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n887), .A2(G290), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(G290), .B1(new_n887), .B2(new_n888), .ZN(new_n890));
  NOR3_X1   g465(.A1(new_n889), .A2(new_n890), .A3(G303), .ZN(new_n891));
  INV_X1    g466(.A(new_n888), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n567), .A2(G305), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n580), .B(new_n579), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n887), .A2(G290), .A3(new_n888), .ZN(new_n895));
  AOI21_X1  g470(.A(G166), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n886), .B1(new_n891), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(G303), .B1(new_n889), .B2(new_n890), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n894), .A2(G166), .A3(new_n895), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT104), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT42), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n891), .A2(new_n896), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n902), .B1(KEYINPUT42), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n905));
  NAND2_X1  g480(.A1(G299), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n560), .A2(KEYINPUT103), .A3(new_n561), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n592), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n584), .A2(new_n589), .A3(new_n591), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n909), .A2(new_n905), .A3(G299), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(KEYINPUT41), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n908), .A2(new_n914), .A3(new_n910), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n843), .B(new_n604), .ZN(new_n917));
  MUX2_X1   g492(.A(new_n912), .B(new_n916), .S(new_n917), .Z(new_n918));
  AND2_X1   g493(.A1(new_n904), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n904), .A2(new_n918), .ZN(new_n920));
  OAI21_X1  g495(.A(G868), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n840), .A2(new_n595), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(G295));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n922), .ZN(G331));
  AND3_X1   g499(.A1(new_n841), .A2(G301), .A3(new_n842), .ZN(new_n925));
  AOI21_X1  g500(.A(G301), .B1(new_n841), .B2(new_n842), .ZN(new_n926));
  OAI21_X1  g501(.A(G286), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n843), .A2(G171), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n841), .A2(G301), .A3(new_n842), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(G168), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n916), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n927), .A2(new_n930), .A3(new_n912), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n932), .A2(new_n897), .A3(new_n900), .A4(new_n933), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n934), .A2(new_n880), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n932), .A2(new_n933), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n901), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT43), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n934), .A2(new_n880), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n911), .A2(KEYINPUT105), .A3(KEYINPUT41), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n931), .B(new_n940), .C1(new_n916), .C2(KEYINPUT105), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n941), .A2(new_n933), .B1(new_n900), .B2(new_n897), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT43), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n939), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT44), .B1(new_n938), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n943), .B1(new_n935), .B2(new_n937), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n939), .A2(new_n942), .A3(KEYINPUT43), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n945), .A2(new_n949), .ZN(G397));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(G164), .B2(G1384), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n463), .A2(new_n467), .A3(G40), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(G1996), .A3(new_n731), .ZN(new_n957));
  XOR2_X1   g532(.A(new_n957), .B(KEYINPUT107), .Z(new_n958));
  XNOR2_X1  g533(.A(new_n711), .B(G2067), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n955), .A2(G1996), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT106), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n958), .B(new_n960), .C1(new_n731), .C2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(G290), .A2(G1986), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n579), .A2(new_n580), .A3(new_n806), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n955), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OR2_X1    g541(.A1(new_n812), .A2(new_n816), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n812), .A2(new_n816), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n955), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n963), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT49), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n572), .A2(new_n972), .A3(new_n575), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n972), .B1(new_n572), .B2(new_n575), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n678), .B1(new_n975), .B2(new_n574), .ZN(new_n976));
  XOR2_X1   g551(.A(KEYINPUT110), .B(G1981), .Z(new_n977));
  NAND4_X1  g552(.A1(new_n572), .A2(new_n575), .A3(new_n574), .A4(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT111), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n971), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  XOR2_X1   g555(.A(new_n978), .B(KEYINPUT111), .Z(new_n981));
  NAND2_X1  g556(.A1(new_n572), .A2(new_n575), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT112), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n572), .A2(new_n972), .A3(new_n575), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(new_n574), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(G1981), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n981), .A2(KEYINPUT49), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n618), .A2(KEYINPUT3), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT3), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(G2104), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n988), .A2(new_n990), .A3(G126), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n462), .B1(new_n991), .B2(new_n487), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT4), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n491), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n484), .A2(new_n485), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n462), .ZN(new_n996));
  AOI21_X1  g571(.A(G1384), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n954), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT109), .B(G8), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n980), .A2(new_n987), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n567), .A2(G1976), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n1002), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT52), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n1008));
  AND3_X1   g583(.A1(G303), .A2(new_n1008), .A3(G8), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1008), .B1(G303), .B2(G8), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G8), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n463), .A2(new_n467), .A3(G40), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n994), .A2(new_n996), .ZN(new_n1014));
  INV_X1    g589(.A(G1384), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1013), .B1(new_n1016), .B2(KEYINPUT50), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1014), .A2(new_n1018), .A3(new_n1015), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT108), .ZN(new_n1020));
  INV_X1    g595(.A(G2090), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT108), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n997), .A2(new_n1022), .A3(new_n1018), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1017), .A2(new_n1020), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1014), .A2(KEYINPUT45), .A3(new_n1015), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n952), .A2(new_n954), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1971), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1012), .B1(new_n1024), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1011), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1017), .A2(new_n1021), .A3(new_n1019), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1001), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n1011), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G1976), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT52), .B1(G288), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1035), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1007), .A2(new_n1030), .A3(new_n1033), .A4(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT121), .ZN(new_n1038));
  AND2_X1   g613(.A1(G286), .A2(new_n1000), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1039), .A2(KEYINPUT51), .ZN(new_n1040));
  INV_X1    g615(.A(G2084), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1017), .A2(new_n1020), .A3(new_n1041), .A4(new_n1023), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1026), .A2(new_n693), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1038), .B(new_n1040), .C1(new_n1044), .C2(new_n1001), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1012), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT51), .B1(new_n1046), .B2(new_n1039), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1001), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT51), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(G168), .B2(new_n1001), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT121), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1045), .A2(new_n1047), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1048), .A2(G286), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G2078), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n952), .A2(new_n1055), .A3(new_n954), .A4(new_n1025), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1017), .A2(new_n1020), .A3(new_n1023), .ZN(new_n1059));
  INV_X1    g634(.A(G1961), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT123), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1063), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1056), .A2(new_n1063), .A3(new_n1057), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1062), .B(G301), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT53), .B1(new_n1013), .B2(KEYINPUT125), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1067), .B1(KEYINPUT125), .B2(new_n1013), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1068), .A2(new_n1055), .A3(new_n952), .A4(new_n1025), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1069), .B(new_n1061), .C1(new_n1065), .C2(new_n1064), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G171), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1066), .A2(new_n1071), .A3(KEYINPUT54), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1054), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1065), .A2(new_n1064), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1075));
  OAI21_X1  g650(.A(G171), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT124), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1070), .A2(G171), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  XOR2_X1   g656(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1082));
  AOI21_X1  g657(.A(new_n1073), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT61), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n557), .A2(new_n559), .ZN(new_n1085));
  INV_X1    g660(.A(new_n554), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n561), .A2(new_n1085), .A3(KEYINPUT57), .A4(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n560), .A2(new_n561), .A3(KEYINPUT117), .A4(KEYINPUT57), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT115), .B(G1956), .Z(new_n1092));
  OAI21_X1  g667(.A(new_n954), .B1(new_n997), .B2(new_n1018), .ZN(new_n1093));
  NOR3_X1   g668(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1092), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT118), .B(G2072), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1096), .B(KEYINPUT56), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n952), .A2(new_n954), .A3(new_n1025), .A4(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1100), .B1(G299), .B2(new_n1101), .ZN(new_n1102));
  AOI211_X1 g677(.A(KEYINPUT116), .B(KEYINPUT57), .C1(new_n560), .C2(new_n561), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1091), .B(new_n1099), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n521), .A2(G91), .A3(new_n523), .ZN(new_n1106));
  AND4_X1   g681(.A1(new_n558), .A2(new_n522), .A3(G53), .A4(new_n555), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n558), .B1(new_n502), .B2(G53), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1086), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1101), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT116), .ZN(new_n1111));
  NAND3_X1  g686(.A1(G299), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1099), .B1(new_n1113), .B2(new_n1091), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1084), .B1(new_n1105), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n998), .A2(G2067), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1116), .B1(new_n1059), .B2(new_n689), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1117), .A2(new_n909), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(new_n909), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT60), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT58), .B(G1341), .ZN(new_n1121));
  OAI22_X1  g696(.A1(new_n1026), .A2(G1996), .B1(new_n999), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n545), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1123), .A2(KEYINPUT119), .A3(KEYINPUT59), .ZN(new_n1124));
  NAND2_X1  g699(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1122), .A2(new_n545), .A3(new_n1125), .ZN(new_n1126));
  AOI211_X1 g701(.A(KEYINPUT60), .B(new_n1116), .C1(new_n1059), .C2(new_n689), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1124), .A2(new_n1126), .B1(new_n1127), .B2(new_n592), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1090), .ZN(new_n1130));
  OAI22_X1  g705(.A1(new_n1129), .A2(new_n1130), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1099), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1133), .A2(KEYINPUT61), .A3(new_n1104), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1115), .A2(new_n1120), .A3(new_n1128), .A4(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1105), .B1(new_n1133), .B2(new_n1119), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1135), .A2(KEYINPUT120), .A3(new_n1136), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1083), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1054), .B(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1037), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT113), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1148));
  OAI211_X1 g723(.A(G168), .B(new_n1048), .C1(new_n1148), .C2(new_n1029), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1148), .A2(new_n1029), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1151), .A2(new_n1003), .A3(new_n1006), .A4(new_n1036), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT63), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT63), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1154), .B1(new_n1011), .B2(new_n1032), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1048), .A2(G168), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1030), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1003), .A2(new_n1157), .A3(new_n1006), .A4(new_n1036), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n567), .A2(new_n1034), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1159), .B1(new_n980), .B2(new_n987), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1002), .B1(new_n1160), .B2(new_n979), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1153), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT114), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT114), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1153), .A2(new_n1164), .A3(new_n1158), .A4(new_n1161), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n970), .B1(new_n1146), .B2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n965), .A2(new_n955), .ZN(new_n1168));
  XOR2_X1   g743(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1169));
  XNOR2_X1  g744(.A(new_n1168), .B(new_n1169), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n963), .A2(new_n969), .A3(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n956), .B1(new_n959), .B2(new_n731), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n962), .A2(KEYINPUT46), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n962), .A2(KEYINPUT46), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1172), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n1175), .B(KEYINPUT47), .Z(new_n1176));
  OAI22_X1  g751(.A1(new_n963), .A2(new_n967), .B1(G2067), .B2(new_n711), .ZN(new_n1177));
  AOI211_X1 g752(.A(new_n1171), .B(new_n1176), .C1(new_n956), .C2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1167), .A2(new_n1178), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n1181));
  INV_X1    g755(.A(G319), .ZN(new_n1182));
  NOR2_X1   g756(.A1(G227), .A2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g757(.A1(new_n685), .A2(new_n1181), .A3(new_n645), .A4(new_n1183), .ZN(new_n1184));
  NAND2_X1  g758(.A1(new_n884), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g759(.A1(new_n685), .A2(new_n645), .A3(new_n1183), .ZN(new_n1186));
  AND2_X1   g760(.A1(new_n1186), .A2(KEYINPUT127), .ZN(new_n1187));
  NAND3_X1  g761(.A1(new_n937), .A2(new_n880), .A3(new_n934), .ZN(new_n1188));
  NAND2_X1  g762(.A1(new_n1188), .A2(KEYINPUT43), .ZN(new_n1189));
  INV_X1    g763(.A(new_n942), .ZN(new_n1190));
  NAND3_X1  g764(.A1(new_n935), .A2(new_n1190), .A3(new_n943), .ZN(new_n1191));
  AOI211_X1 g765(.A(new_n1185), .B(new_n1187), .C1(new_n1189), .C2(new_n1191), .ZN(G308));
  AOI21_X1  g766(.A(new_n1187), .B1(new_n1191), .B2(new_n1189), .ZN(new_n1193));
  INV_X1    g767(.A(new_n1185), .ZN(new_n1194));
  NAND2_X1  g768(.A1(new_n1193), .A2(new_n1194), .ZN(G225));
endmodule


