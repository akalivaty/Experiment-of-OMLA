

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805;

  BUF_X1 U374 ( .A(n803), .Z(n352) );
  AND2_X1 U375 ( .A1(n805), .A2(n602), .ZN(n603) );
  AND2_X1 U376 ( .A1(n589), .A2(n633), .ZN(n463) );
  BUF_X1 U377 ( .A(n591), .Z(n353) );
  NOR2_X1 U378 ( .A1(n734), .A2(n735), .ZN(n648) );
  NAND2_X1 U379 ( .A1(n617), .A2(n552), .ZN(n553) );
  INV_X1 U380 ( .A(n719), .ZN(n625) );
  NOR2_X1 U381 ( .A1(n599), .A2(n600), .ZN(n704) );
  NOR2_X2 U382 ( .A1(n658), .A2(n546), .ZN(n355) );
  NAND2_X1 U383 ( .A1(n591), .A2(n483), .ZN(n719) );
  INV_X1 U384 ( .A(KEYINPUT19), .ZN(n354) );
  XNOR2_X1 U385 ( .A(G131), .B(G134), .ZN(n440) );
  XNOR2_X1 U386 ( .A(G119), .B(G110), .ZN(n510) );
  XNOR2_X2 U387 ( .A(n355), .B(n354), .ZN(n617) );
  NOR2_X1 U388 ( .A1(n429), .A2(n699), .ZN(n632) );
  NOR2_X1 U389 ( .A1(n704), .A2(n702), .ZN(n736) );
  XOR2_X1 U390 ( .A(G107), .B(G104), .Z(n496) );
  XNOR2_X1 U391 ( .A(n783), .B(KEYINPUT69), .ZN(n528) );
  AND2_X1 U392 ( .A1(n386), .A2(n624), .ZN(n626) );
  AND2_X2 U393 ( .A1(n434), .A2(n371), .ZN(n433) );
  XNOR2_X1 U394 ( .A(n441), .B(n440), .ZN(n439) );
  XNOR2_X1 U395 ( .A(n473), .B(G137), .ZN(n441) );
  NOR2_X2 U396 ( .A1(n759), .A2(G902), .ZN(n418) );
  XNOR2_X2 U397 ( .A(n525), .B(KEYINPUT91), .ZN(n788) );
  INV_X1 U398 ( .A(n713), .ZN(n591) );
  INV_X1 U399 ( .A(n594), .ZN(n717) );
  AND2_X1 U400 ( .A1(n599), .A2(n600), .ZN(n702) );
  XNOR2_X1 U401 ( .A(n524), .B(n523), .ZN(n538) );
  XNOR2_X1 U402 ( .A(n388), .B(G119), .ZN(n524) );
  XNOR2_X1 U403 ( .A(n563), .B(n769), .ZN(n599) );
  XNOR2_X1 U404 ( .A(n539), .B(n538), .ZN(n782) );
  XNOR2_X1 U405 ( .A(G146), .B(G116), .ZN(n519) );
  INV_X1 U406 ( .A(KEYINPUT30), .ZN(n363) );
  AND2_X1 U407 ( .A1(n488), .A2(n486), .ZN(n485) );
  NAND2_X1 U408 ( .A1(n445), .A2(n373), .ZN(n421) );
  BUF_X1 U409 ( .A(n658), .Z(n356) );
  BUF_X1 U410 ( .A(n788), .Z(n413) );
  XNOR2_X1 U411 ( .A(n424), .B(n423), .ZN(n554) );
  INV_X1 U412 ( .A(KEYINPUT66), .ZN(n473) );
  INV_X2 U413 ( .A(G953), .ZN(n795) );
  NOR2_X1 U414 ( .A1(n686), .A2(n777), .ZN(n688) );
  AND2_X1 U415 ( .A1(n392), .A2(n393), .ZN(n358) );
  XNOR2_X1 U416 ( .A(n364), .B(n363), .ZN(n627) );
  NOR2_X1 U417 ( .A1(n612), .A2(n546), .ZN(n364) );
  XNOR2_X1 U418 ( .A(n402), .B(KEYINPUT86), .ZN(n401) );
  BUF_X1 U419 ( .A(n805), .Z(n357) );
  OR2_X1 U420 ( .A1(n581), .A2(n366), .ZN(n447) );
  XNOR2_X1 U421 ( .A(n646), .B(n381), .ZN(n359) );
  BUF_X1 U422 ( .A(n653), .Z(n360) );
  BUF_X1 U423 ( .A(n386), .Z(n361) );
  XNOR2_X1 U424 ( .A(n646), .B(n381), .ZN(n651) );
  BUF_X1 U425 ( .A(n617), .Z(n362) );
  NAND2_X1 U426 ( .A1(n391), .A2(n390), .ZN(n389) );
  AND2_X1 U427 ( .A1(n619), .A2(n362), .ZN(n428) );
  INV_X1 U428 ( .A(KEYINPUT104), .ZN(n431) );
  XNOR2_X1 U429 ( .A(n736), .B(n459), .ZN(n620) );
  INV_X1 U430 ( .A(KEYINPUT73), .ZN(n459) );
  INV_X1 U431 ( .A(KEYINPUT44), .ZN(n398) );
  NOR2_X1 U432 ( .A1(n400), .A2(n398), .ZN(n397) );
  INV_X1 U433 ( .A(n707), .ZN(n641) );
  INV_X1 U434 ( .A(KEYINPUT46), .ZN(n471) );
  INV_X1 U435 ( .A(KEYINPUT65), .ZN(n400) );
  INV_X1 U436 ( .A(KEYINPUT83), .ZN(n668) );
  NAND2_X1 U437 ( .A1(G234), .A2(G237), .ZN(n547) );
  XNOR2_X1 U438 ( .A(n386), .B(n501), .ZN(n581) );
  NOR2_X1 U439 ( .A1(n751), .A2(n753), .ZN(n752) );
  INV_X1 U440 ( .A(KEYINPUT107), .ZN(n615) );
  NOR2_X1 U441 ( .A1(n453), .A2(n777), .ZN(n452) );
  NOR2_X1 U442 ( .A1(n467), .A2(G472), .ZN(n453) );
  NOR2_X1 U443 ( .A1(n767), .A2(n490), .ZN(n489) );
  INV_X1 U444 ( .A(G475), .ZN(n490) );
  NOR2_X1 U445 ( .A1(n487), .A2(n777), .ZN(n486) );
  NAND2_X1 U446 ( .A1(n450), .A2(n767), .ZN(n484) );
  NAND2_X1 U447 ( .A1(n631), .A2(n430), .ZN(n429) );
  NOR2_X1 U448 ( .A1(n394), .A2(n383), .ZN(n393) );
  NOR2_X1 U449 ( .A1(n590), .A2(n395), .ZN(n394) );
  INV_X1 U450 ( .A(n397), .ZN(n395) );
  NOR2_X1 U451 ( .A1(G953), .A2(G237), .ZN(n567) );
  INV_X1 U452 ( .A(KEYINPUT48), .ZN(n469) );
  NAND2_X1 U453 ( .A1(n374), .A2(n365), .ZN(n390) );
  XOR2_X1 U454 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n569) );
  XNOR2_X1 U455 ( .A(G143), .B(G131), .ZN(n564) );
  XOR2_X1 U456 ( .A(KEYINPUT12), .B(G113), .Z(n565) );
  XNOR2_X1 U457 ( .A(G101), .B(G146), .ZN(n495) );
  INV_X1 U458 ( .A(KEYINPUT33), .ZN(n448) );
  NOR2_X1 U459 ( .A1(G237), .A2(G902), .ZN(n541) );
  XNOR2_X1 U460 ( .A(KEYINPUT97), .B(G472), .ZN(n526) );
  XNOR2_X1 U461 ( .A(G101), .B(KEYINPUT68), .ZN(n523) );
  INV_X1 U462 ( .A(G116), .ZN(n536) );
  XNOR2_X1 U463 ( .A(KEYINPUT10), .B(G140), .ZN(n477) );
  INV_X1 U464 ( .A(KEYINPUT8), .ZN(n423) );
  NAND2_X1 U465 ( .A1(n795), .A2(G234), .ZN(n424) );
  XOR2_X1 U466 ( .A(KEYINPUT24), .B(KEYINPUT92), .Z(n511) );
  XOR2_X1 U467 ( .A(n457), .B(G137), .Z(n513) );
  XNOR2_X1 U468 ( .A(G134), .B(G122), .ZN(n555) );
  XOR2_X1 U469 ( .A(KEYINPUT7), .B(KEYINPUT101), .Z(n556) );
  INV_X1 U470 ( .A(G210), .ZN(n681) );
  INV_X1 U471 ( .A(G902), .ZN(n562) );
  INV_X1 U472 ( .A(G469), .ZN(n417) );
  BUF_X1 U473 ( .A(n581), .Z(n720) );
  AND2_X1 U474 ( .A1(n464), .A2(n370), .ZN(n755) );
  XNOR2_X1 U475 ( .A(n425), .B(KEYINPUT42), .ZN(n803) );
  XNOR2_X1 U476 ( .A(n416), .B(n415), .ZN(n705) );
  INV_X1 U477 ( .A(KEYINPUT31), .ZN(n415) );
  AND2_X1 U478 ( .A1(n454), .A2(n452), .ZN(n451) );
  NAND2_X1 U479 ( .A1(n450), .A2(n676), .ZN(n449) );
  INV_X1 U480 ( .A(KEYINPUT60), .ZN(n491) );
  AND2_X1 U481 ( .A1(n679), .A2(n590), .ZN(n365) );
  AND2_X1 U482 ( .A1(n591), .A2(n379), .ZN(n366) );
  NOR2_X1 U483 ( .A1(n597), .A2(n411), .ZN(n367) );
  XOR2_X1 U484 ( .A(n582), .B(KEYINPUT103), .Z(n368) );
  OR2_X1 U485 ( .A1(n791), .A2(n753), .ZN(n369) );
  OR2_X1 U486 ( .A1(n748), .A2(n747), .ZN(n370) );
  AND2_X1 U487 ( .A1(n435), .A2(n577), .ZN(n371) );
  AND2_X1 U488 ( .A1(n720), .A2(n353), .ZN(n372) );
  AND2_X1 U489 ( .A1(n637), .A2(n480), .ZN(n373) );
  NOR2_X1 U490 ( .A1(n800), .A2(KEYINPUT44), .ZN(n374) );
  XNOR2_X1 U491 ( .A(KEYINPUT100), .B(KEYINPUT9), .ZN(n375) );
  AND2_X1 U492 ( .A1(n567), .A2(G210), .ZN(n376) );
  NOR2_X1 U493 ( .A1(n750), .A2(G953), .ZN(n377) );
  AND2_X1 U494 ( .A1(n590), .A2(n400), .ZN(n378) );
  AND2_X1 U495 ( .A1(n483), .A2(KEYINPUT105), .ZN(n379) );
  AND2_X1 U496 ( .A1(n660), .A2(KEYINPUT2), .ZN(n380) );
  XNOR2_X1 U497 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n381) );
  XOR2_X1 U498 ( .A(n580), .B(KEYINPUT22), .Z(n382) );
  AND2_X1 U499 ( .A1(n400), .A2(n398), .ZN(n383) );
  INV_X1 U500 ( .A(KEYINPUT105), .ZN(n481) );
  AND2_X1 U501 ( .A1(n467), .A2(G472), .ZN(n384) );
  AND2_X1 U502 ( .A1(n677), .A2(G953), .ZN(n777) );
  NOR2_X1 U503 ( .A1(n385), .A2(G902), .ZN(n527) );
  XNOR2_X1 U504 ( .A(n385), .B(n675), .ZN(n676) );
  XNOR2_X1 U505 ( .A(n474), .B(n405), .ZN(n385) );
  AND2_X1 U506 ( .A1(n625), .A2(n361), .ZN(n595) );
  NAND2_X1 U507 ( .A1(n614), .A2(n361), .ZN(n616) );
  XNOR2_X2 U508 ( .A(n418), .B(n417), .ZN(n386) );
  XNOR2_X1 U509 ( .A(n788), .B(n528), .ZN(n387) );
  XNOR2_X2 U510 ( .A(n439), .B(n529), .ZN(n525) );
  XNOR2_X1 U511 ( .A(n387), .B(n500), .ZN(n759) );
  XNOR2_X2 U512 ( .A(G113), .B(KEYINPUT3), .ZN(n388) );
  NOR2_X2 U513 ( .A1(n389), .A2(n401), .ZN(n605) );
  NAND2_X1 U514 ( .A1(n358), .A2(n396), .ZN(n391) );
  NAND2_X1 U515 ( .A1(n679), .A2(n378), .ZN(n392) );
  NAND2_X1 U516 ( .A1(n399), .A2(n397), .ZN(n396) );
  INV_X1 U517 ( .A(n679), .ZN(n399) );
  NAND2_X1 U518 ( .A1(n604), .A2(n603), .ZN(n402) );
  INV_X1 U519 ( .A(n476), .ZN(n713) );
  BUF_X1 U520 ( .A(n683), .Z(n403) );
  NOR2_X2 U521 ( .A1(n727), .A2(n411), .ZN(n416) );
  XNOR2_X1 U522 ( .A(n421), .B(n448), .ZN(n404) );
  XNOR2_X1 U523 ( .A(n421), .B(n448), .ZN(n710) );
  AND2_X1 U524 ( .A1(n468), .A2(n660), .ZN(n662) );
  XNOR2_X1 U525 ( .A(n419), .B(n469), .ZN(n468) );
  AND2_X1 U526 ( .A1(n444), .A2(n791), .ZN(n665) );
  BUF_X1 U527 ( .A(n525), .Z(n405) );
  XNOR2_X1 U528 ( .A(n669), .B(n668), .ZN(n670) );
  NAND2_X1 U529 ( .A1(n540), .A2(n782), .ZN(n408) );
  NAND2_X1 U530 ( .A1(n406), .A2(n407), .ZN(n409) );
  NAND2_X1 U531 ( .A1(n409), .A2(n408), .ZN(n683) );
  INV_X1 U532 ( .A(n540), .ZN(n406) );
  INV_X1 U533 ( .A(n782), .ZN(n407) );
  NOR2_X1 U534 ( .A1(n711), .A2(n649), .ZN(n425) );
  XNOR2_X1 U535 ( .A(n553), .B(KEYINPUT0), .ZN(n410) );
  XNOR2_X1 U536 ( .A(n553), .B(KEYINPUT0), .ZN(n411) );
  XNOR2_X1 U537 ( .A(n553), .B(KEYINPUT0), .ZN(n596) );
  XNOR2_X2 U538 ( .A(n585), .B(n584), .ZN(n679) );
  INV_X1 U539 ( .A(n768), .ZN(n765) );
  OR2_X1 U540 ( .A1(n356), .A2(n546), .ZN(n412) );
  XNOR2_X1 U541 ( .A(n516), .B(n515), .ZN(n773) );
  XNOR2_X1 U542 ( .A(n442), .B(n531), .ZN(n532) );
  XOR2_X1 U543 ( .A(G143), .B(G128), .Z(n414) );
  BUF_X1 U544 ( .A(G128), .Z(n457) );
  NAND2_X1 U545 ( .A1(n437), .A2(n436), .ZN(n432) );
  XNOR2_X1 U546 ( .A(n443), .B(n382), .ZN(n589) );
  INV_X1 U547 ( .A(n612), .ZN(n622) );
  NOR2_X1 U548 ( .A1(n410), .A2(KEYINPUT34), .ZN(n436) );
  NAND2_X1 U549 ( .A1(n470), .A2(n472), .ZN(n419) );
  NOR2_X2 U550 ( .A1(n627), .A2(n420), .ZN(n628) );
  NAND2_X1 U551 ( .A1(n626), .A2(n625), .ZN(n420) );
  OR2_X2 U552 ( .A1(n601), .A2(n736), .ZN(n602) );
  XNOR2_X2 U553 ( .A(n592), .B(KEYINPUT102), .ZN(n805) );
  XNOR2_X1 U554 ( .A(n494), .B(n789), .ZN(n516) );
  XNOR2_X1 U555 ( .A(n422), .B(KEYINPUT67), .ZN(n472) );
  NAND2_X1 U556 ( .A1(n642), .A2(n641), .ZN(n422) );
  XNOR2_X1 U557 ( .A(n517), .B(n518), .ZN(n476) );
  XNOR2_X2 U558 ( .A(KEYINPUT15), .B(G902), .ZN(n663) );
  NAND2_X1 U559 ( .A1(n749), .A2(n661), .ZN(n478) );
  XNOR2_X2 U560 ( .A(n605), .B(KEYINPUT45), .ZN(n749) );
  NAND2_X1 U561 ( .A1(n426), .A2(KEYINPUT47), .ZN(n430) );
  NAND2_X1 U562 ( .A1(n427), .A2(n428), .ZN(n426) );
  INV_X1 U563 ( .A(n649), .ZN(n427) );
  NOR2_X2 U564 ( .A1(n649), .A2(n618), .ZN(n700) );
  AND2_X1 U565 ( .A1(n643), .A2(n630), .ZN(n699) );
  XNOR2_X2 U566 ( .A(n586), .B(n431), .ZN(n612) );
  XNOR2_X2 U567 ( .A(n527), .B(n526), .ZN(n586) );
  NAND2_X2 U568 ( .A1(n433), .A2(n432), .ZN(n438) );
  NAND2_X1 U569 ( .A1(n710), .A2(KEYINPUT34), .ZN(n434) );
  NAND2_X1 U570 ( .A1(n410), .A2(KEYINPUT34), .ZN(n435) );
  INV_X1 U571 ( .A(n404), .ZN(n437) );
  XNOR2_X2 U572 ( .A(n438), .B(KEYINPUT35), .ZN(n800) );
  XNOR2_X2 U573 ( .A(n559), .B(KEYINPUT4), .ZN(n529) );
  XNOR2_X2 U574 ( .A(G143), .B(G128), .ZN(n559) );
  XNOR2_X1 U575 ( .A(n442), .B(n477), .ZN(n789) );
  XNOR2_X2 U576 ( .A(n509), .B(G146), .ZN(n442) );
  NAND2_X1 U577 ( .A1(n463), .A2(n372), .ZN(n592) );
  NOR2_X2 U578 ( .A1(n596), .A2(n579), .ZN(n443) );
  NAND2_X1 U579 ( .A1(n444), .A2(KEYINPUT2), .ZN(n666) );
  NAND2_X1 U580 ( .A1(n664), .A2(n663), .ZN(n444) );
  NAND2_X1 U581 ( .A1(n447), .A2(n446), .ZN(n445) );
  NAND2_X1 U582 ( .A1(n581), .A2(KEYINPUT105), .ZN(n446) );
  NAND2_X1 U583 ( .A1(n451), .A2(n449), .ZN(n455) );
  INV_X1 U584 ( .A(n674), .ZN(n450) );
  NAND2_X1 U585 ( .A1(n674), .A2(n384), .ZN(n454) );
  XNOR2_X1 U586 ( .A(n455), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U587 ( .A(n534), .B(n456), .ZN(n540) );
  XNOR2_X1 U588 ( .A(n532), .B(n533), .ZN(n456) );
  NAND2_X2 U589 ( .A1(n653), .A2(n702), .ZN(n646) );
  NAND2_X1 U590 ( .A1(n458), .A2(n665), .ZN(n667) );
  NAND2_X1 U591 ( .A1(n479), .A2(n478), .ZN(n458) );
  NAND2_X1 U592 ( .A1(n468), .A2(n380), .ZN(n669) );
  XNOR2_X1 U593 ( .A(n461), .B(n460), .ZN(n770) );
  XNOR2_X1 U594 ( .A(n557), .B(n375), .ZN(n460) );
  XNOR2_X1 U595 ( .A(n462), .B(n561), .ZN(n461) );
  NAND2_X1 U596 ( .A1(n554), .A2(G217), .ZN(n462) );
  NAND2_X1 U597 ( .A1(n463), .A2(n368), .ZN(n585) );
  INV_X1 U598 ( .A(n750), .ZN(n751) );
  NAND2_X1 U599 ( .A1(n466), .A2(n465), .ZN(n464) );
  AND2_X1 U600 ( .A1(n754), .A2(n369), .ZN(n465) );
  XNOR2_X1 U601 ( .A(n752), .B(KEYINPUT81), .ZN(n466) );
  XNOR2_X1 U602 ( .A(n359), .B(G131), .ZN(n802) );
  INV_X1 U603 ( .A(n676), .ZN(n467) );
  XNOR2_X1 U604 ( .A(n652), .B(n471), .ZN(n470) );
  XNOR2_X1 U605 ( .A(n538), .B(n475), .ZN(n474) );
  XNOR2_X1 U606 ( .A(n522), .B(n376), .ZN(n475) );
  OR2_X2 U607 ( .A1(n749), .A2(n606), .ZN(n479) );
  OR2_X1 U608 ( .A1(n581), .A2(n719), .ZN(n482) );
  NAND2_X1 U609 ( .A1(n719), .A2(n481), .ZN(n480) );
  INV_X1 U610 ( .A(n482), .ZN(n593) );
  INV_X1 U611 ( .A(n578), .ZN(n483) );
  NAND2_X1 U612 ( .A1(n765), .A2(n489), .ZN(n488) );
  NAND2_X1 U613 ( .A1(n485), .A2(n484), .ZN(n492) );
  NOR2_X1 U614 ( .A1(n493), .A2(G475), .ZN(n487) );
  XNOR2_X1 U615 ( .A(n492), .B(n491), .ZN(G60) );
  INV_X1 U616 ( .A(n767), .ZN(n493) );
  NOR2_X1 U617 ( .A1(n612), .A2(n634), .ZN(n613) );
  AND2_X1 U618 ( .A1(G221), .A2(n554), .ZN(n494) );
  INV_X1 U619 ( .A(n803), .ZN(n650) );
  INV_X2 U620 ( .A(G125), .ZN(n509) );
  NOR2_X2 U621 ( .A1(n670), .A2(n749), .ZN(n671) );
  BUF_X1 U622 ( .A(n662), .Z(n791) );
  BUF_X1 U623 ( .A(n404), .Z(n741) );
  BUF_X1 U624 ( .A(n759), .Z(n761) );
  BUF_X1 U625 ( .A(n800), .Z(n801) );
  XNOR2_X2 U626 ( .A(KEYINPUT76), .B(G110), .ZN(n783) );
  XNOR2_X1 U627 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U628 ( .A(G140), .B(n497), .Z(n499) );
  NAND2_X1 U629 ( .A1(G227), .A2(n795), .ZN(n498) );
  XNOR2_X1 U630 ( .A(n499), .B(n498), .ZN(n500) );
  INV_X1 U631 ( .A(KEYINPUT1), .ZN(n501) );
  NAND2_X1 U632 ( .A1(n663), .A2(G234), .ZN(n502) );
  XNOR2_X1 U633 ( .A(n502), .B(KEYINPUT20), .ZN(n505) );
  NAND2_X1 U634 ( .A1(G221), .A2(n505), .ZN(n504) );
  XOR2_X1 U635 ( .A(KEYINPUT95), .B(KEYINPUT21), .Z(n503) );
  XNOR2_X1 U636 ( .A(n504), .B(n503), .ZN(n714) );
  XNOR2_X1 U637 ( .A(n714), .B(KEYINPUT96), .ZN(n578) );
  XOR2_X1 U638 ( .A(KEYINPUT25), .B(KEYINPUT94), .Z(n507) );
  NAND2_X1 U639 ( .A1(n505), .A2(G217), .ZN(n506) );
  XNOR2_X1 U640 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U641 ( .A(KEYINPUT93), .B(n508), .ZN(n518) );
  XNOR2_X1 U642 ( .A(n510), .B(KEYINPUT23), .ZN(n512) );
  XNOR2_X1 U643 ( .A(n512), .B(n511), .ZN(n514) );
  XNOR2_X1 U644 ( .A(n514), .B(n513), .ZN(n515) );
  NOR2_X1 U645 ( .A1(G902), .A2(n773), .ZN(n517) );
  INV_X1 U646 ( .A(n519), .ZN(n521) );
  XNOR2_X1 U647 ( .A(KEYINPUT75), .B(KEYINPUT5), .ZN(n520) );
  XNOR2_X1 U648 ( .A(n521), .B(n520), .ZN(n522) );
  INV_X1 U649 ( .A(n586), .ZN(n594) );
  XNOR2_X1 U650 ( .A(n717), .B(KEYINPUT6), .ZN(n633) );
  XNOR2_X1 U651 ( .A(n529), .B(n528), .ZN(n534) );
  NAND2_X1 U652 ( .A1(n795), .A2(G224), .ZN(n530) );
  XNOR2_X1 U653 ( .A(n530), .B(KEYINPUT87), .ZN(n533) );
  XNOR2_X1 U654 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n531) );
  XNOR2_X2 U655 ( .A(G122), .B(G104), .ZN(n570) );
  XNOR2_X1 U656 ( .A(KEYINPUT71), .B(KEYINPUT16), .ZN(n535) );
  XNOR2_X1 U657 ( .A(n570), .B(n535), .ZN(n537) );
  XNOR2_X1 U658 ( .A(n536), .B(G107), .ZN(n558) );
  XNOR2_X1 U659 ( .A(n537), .B(n558), .ZN(n539) );
  NAND2_X1 U660 ( .A1(n683), .A2(n663), .ZN(n543) );
  XNOR2_X1 U661 ( .A(n541), .B(KEYINPUT74), .ZN(n545) );
  OR2_X1 U662 ( .A1(n545), .A2(n681), .ZN(n542) );
  XNOR2_X2 U663 ( .A(n543), .B(n542), .ZN(n658) );
  INV_X1 U664 ( .A(G214), .ZN(n544) );
  OR2_X1 U665 ( .A1(n545), .A2(n544), .ZN(n731) );
  INV_X1 U666 ( .A(n731), .ZN(n546) );
  XNOR2_X1 U667 ( .A(n547), .B(KEYINPUT88), .ZN(n548) );
  XNOR2_X1 U668 ( .A(KEYINPUT14), .B(n548), .ZN(n550) );
  NAND2_X1 U669 ( .A1(G902), .A2(n550), .ZN(n607) );
  XNOR2_X1 U670 ( .A(G898), .B(KEYINPUT89), .ZN(n780) );
  NAND2_X1 U671 ( .A1(G953), .A2(n780), .ZN(n784) );
  NOR2_X1 U672 ( .A1(n607), .A2(n784), .ZN(n549) );
  XNOR2_X1 U673 ( .A(n549), .B(KEYINPUT90), .ZN(n551) );
  NAND2_X1 U674 ( .A1(G952), .A2(n550), .ZN(n748) );
  NOR2_X1 U675 ( .A1(n748), .A2(G953), .ZN(n610) );
  OR2_X1 U676 ( .A1(n551), .A2(n610), .ZN(n552) );
  XNOR2_X1 U677 ( .A(n556), .B(n555), .ZN(n557) );
  INV_X1 U678 ( .A(n558), .ZN(n560) );
  XNOR2_X1 U679 ( .A(n560), .B(n414), .ZN(n561) );
  NAND2_X1 U680 ( .A1(n770), .A2(n562), .ZN(n563) );
  INV_X1 U681 ( .A(G478), .ZN(n769) );
  XNOR2_X1 U682 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U683 ( .A(n789), .B(n566), .ZN(n574) );
  NAND2_X1 U684 ( .A1(G214), .A2(n567), .ZN(n568) );
  XNOR2_X1 U685 ( .A(n569), .B(n568), .ZN(n572) );
  XOR2_X1 U686 ( .A(KEYINPUT11), .B(n570), .Z(n571) );
  XNOR2_X1 U687 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U688 ( .A(n574), .B(n573), .ZN(n766) );
  NOR2_X1 U689 ( .A1(G902), .A2(n766), .ZN(n576) );
  XOR2_X1 U690 ( .A(KEYINPUT13), .B(G475), .Z(n575) );
  XNOR2_X1 U691 ( .A(n576), .B(n575), .ZN(n598) );
  OR2_X1 U692 ( .A1(n599), .A2(n598), .ZN(n629) );
  INV_X1 U693 ( .A(n629), .ZN(n577) );
  NAND2_X1 U694 ( .A1(n599), .A2(n598), .ZN(n734) );
  OR2_X1 U695 ( .A1(n734), .A2(n578), .ZN(n579) );
  INV_X1 U696 ( .A(KEYINPUT70), .ZN(n580) );
  NOR2_X1 U697 ( .A1(n720), .A2(n353), .ZN(n582) );
  INV_X1 U698 ( .A(KEYINPUT79), .ZN(n583) );
  XNOR2_X1 U699 ( .A(n583), .B(KEYINPUT32), .ZN(n584) );
  NOR2_X1 U700 ( .A1(n353), .A2(n622), .ZN(n587) );
  AND2_X1 U701 ( .A1(n720), .A2(n587), .ZN(n588) );
  AND2_X1 U702 ( .A1(n589), .A2(n588), .ZN(n696) );
  INV_X1 U703 ( .A(n696), .ZN(n590) );
  NAND2_X1 U704 ( .A1(n800), .A2(KEYINPUT44), .ZN(n604) );
  NAND2_X1 U705 ( .A1(n593), .A2(n717), .ZN(n727) );
  NAND2_X1 U706 ( .A1(n595), .A2(n594), .ZN(n597) );
  NOR2_X1 U707 ( .A1(n705), .A2(n367), .ZN(n601) );
  INV_X1 U708 ( .A(n598), .ZN(n600) );
  NOR2_X1 U709 ( .A1(n663), .A2(KEYINPUT82), .ZN(n606) );
  INV_X1 U710 ( .A(KEYINPUT82), .ZN(n661) );
  OR2_X1 U711 ( .A1(n795), .A2(n607), .ZN(n608) );
  NOR2_X1 U712 ( .A1(G900), .A2(n608), .ZN(n609) );
  NOR2_X1 U713 ( .A1(n610), .A2(n609), .ZN(n623) );
  NOR2_X1 U714 ( .A1(n714), .A2(n623), .ZN(n611) );
  NAND2_X1 U715 ( .A1(n611), .A2(n713), .ZN(n634) );
  XNOR2_X1 U716 ( .A(n613), .B(KEYINPUT28), .ZN(n614) );
  XNOR2_X2 U717 ( .A(n616), .B(n615), .ZN(n649) );
  INV_X1 U718 ( .A(n362), .ZN(n618) );
  NOR2_X1 U719 ( .A1(n736), .A2(KEYINPUT73), .ZN(n619) );
  NOR2_X1 U720 ( .A1(KEYINPUT47), .A2(n620), .ZN(n621) );
  NAND2_X1 U721 ( .A1(n700), .A2(n621), .ZN(n631) );
  INV_X1 U722 ( .A(n623), .ZN(n624) );
  XNOR2_X1 U723 ( .A(n628), .B(KEYINPUT78), .ZN(n643) );
  NOR2_X1 U724 ( .A1(n356), .A2(n629), .ZN(n630) );
  XNOR2_X1 U725 ( .A(n632), .B(KEYINPUT72), .ZN(n642) );
  INV_X1 U726 ( .A(n633), .ZN(n637) );
  INV_X1 U727 ( .A(n702), .ZN(n635) );
  NOR2_X1 U728 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U729 ( .A1(n637), .A2(n636), .ZN(n655) );
  NOR2_X1 U730 ( .A1(n655), .A2(n412), .ZN(n639) );
  XOR2_X1 U731 ( .A(KEYINPUT36), .B(n639), .Z(n640) );
  NOR2_X1 U732 ( .A1(n720), .A2(n640), .ZN(n707) );
  XNOR2_X1 U733 ( .A(n658), .B(KEYINPUT38), .ZN(n732) );
  NAND2_X1 U734 ( .A1(n643), .A2(n732), .ZN(n645) );
  XOR2_X1 U735 ( .A(KEYINPUT85), .B(KEYINPUT39), .Z(n644) );
  XNOR2_X2 U736 ( .A(n645), .B(n644), .ZN(n653) );
  NAND2_X1 U737 ( .A1(n732), .A2(n731), .ZN(n735) );
  XNOR2_X1 U738 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n647) );
  XNOR2_X1 U739 ( .A(n648), .B(n647), .ZN(n729) );
  INV_X1 U740 ( .A(n729), .ZN(n711) );
  NAND2_X1 U741 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U742 ( .A1(n704), .A2(n360), .ZN(n709) );
  NAND2_X1 U743 ( .A1(n720), .A2(n731), .ZN(n654) );
  NOR2_X1 U744 ( .A1(n655), .A2(n654), .ZN(n657) );
  XNOR2_X1 U745 ( .A(KEYINPUT43), .B(KEYINPUT106), .ZN(n656) );
  XOR2_X1 U746 ( .A(n657), .B(n656), .Z(n659) );
  NAND2_X1 U747 ( .A1(n659), .A2(n356), .ZN(n678) );
  AND2_X1 U748 ( .A1(n709), .A2(n678), .ZN(n660) );
  NAND2_X1 U749 ( .A1(n662), .A2(n661), .ZN(n664) );
  NAND2_X1 U750 ( .A1(n667), .A2(n666), .ZN(n672) );
  XNOR2_X1 U751 ( .A(n671), .B(KEYINPUT77), .ZN(n754) );
  NAND2_X1 U752 ( .A1(n672), .A2(n754), .ZN(n673) );
  XNOR2_X2 U753 ( .A(n673), .B(KEYINPUT64), .ZN(n768) );
  INV_X1 U754 ( .A(n768), .ZN(n674) );
  XNOR2_X1 U755 ( .A(KEYINPUT110), .B(KEYINPUT62), .ZN(n675) );
  INV_X1 U756 ( .A(G952), .ZN(n677) );
  XNOR2_X1 U757 ( .A(n678), .B(G140), .ZN(G42) );
  XOR2_X1 U758 ( .A(G119), .B(KEYINPUT124), .Z(n680) );
  XOR2_X1 U759 ( .A(n680), .B(n679), .Z(G21) );
  NOR2_X1 U760 ( .A1(n768), .A2(n681), .ZN(n685) );
  XOR2_X1 U761 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n682) );
  XNOR2_X1 U762 ( .A(n403), .B(n682), .ZN(n684) );
  XNOR2_X1 U763 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U764 ( .A(KEYINPUT84), .B(KEYINPUT56), .ZN(n687) );
  XNOR2_X1 U765 ( .A(n688), .B(n687), .ZN(G51) );
  XOR2_X1 U766 ( .A(G104), .B(KEYINPUT111), .Z(n690) );
  NAND2_X1 U767 ( .A1(n367), .A2(n702), .ZN(n689) );
  XNOR2_X1 U768 ( .A(n690), .B(n689), .ZN(G6) );
  XOR2_X1 U769 ( .A(KEYINPUT113), .B(KEYINPUT27), .Z(n692) );
  XNOR2_X1 U770 ( .A(G107), .B(KEYINPUT26), .ZN(n691) );
  XNOR2_X1 U771 ( .A(n692), .B(n691), .ZN(n693) );
  XOR2_X1 U772 ( .A(KEYINPUT112), .B(n693), .Z(n695) );
  NAND2_X1 U773 ( .A1(n367), .A2(n704), .ZN(n694) );
  XNOR2_X1 U774 ( .A(n695), .B(n694), .ZN(G9) );
  XOR2_X1 U775 ( .A(G110), .B(n696), .Z(G12) );
  XOR2_X1 U776 ( .A(n457), .B(KEYINPUT29), .Z(n698) );
  NAND2_X1 U777 ( .A1(n700), .A2(n704), .ZN(n697) );
  XNOR2_X1 U778 ( .A(n698), .B(n697), .ZN(G30) );
  XOR2_X1 U779 ( .A(G143), .B(n699), .Z(G45) );
  NAND2_X1 U780 ( .A1(n700), .A2(n702), .ZN(n701) );
  XNOR2_X1 U781 ( .A(n701), .B(G146), .ZN(G48) );
  NAND2_X1 U782 ( .A1(n705), .A2(n702), .ZN(n703) );
  XNOR2_X1 U783 ( .A(n703), .B(G113), .ZN(G15) );
  NAND2_X1 U784 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U785 ( .A(n706), .B(G116), .ZN(G18) );
  XNOR2_X1 U786 ( .A(G125), .B(n707), .ZN(n708) );
  XNOR2_X1 U787 ( .A(n708), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U788 ( .A(G134), .B(n709), .ZN(G36) );
  XOR2_X1 U789 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n758) );
  NOR2_X1 U790 ( .A1(n741), .A2(n711), .ZN(n712) );
  NOR2_X1 U791 ( .A1(G953), .A2(n712), .ZN(n756) );
  NAND2_X1 U792 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U793 ( .A(KEYINPUT49), .B(n715), .ZN(n716) );
  NOR2_X1 U794 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U795 ( .A(KEYINPUT114), .B(n718), .ZN(n725) );
  XOR2_X1 U796 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n722) );
  NAND2_X1 U797 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U798 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U799 ( .A(KEYINPUT115), .B(n723), .ZN(n724) );
  NAND2_X1 U800 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U801 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U802 ( .A(KEYINPUT51), .B(n728), .Z(n730) );
  NAND2_X1 U803 ( .A1(n730), .A2(n729), .ZN(n744) );
  NOR2_X1 U804 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U805 ( .A1(n734), .A2(n733), .ZN(n738) );
  NOR2_X1 U806 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U807 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U808 ( .A(KEYINPUT117), .B(n739), .Z(n740) );
  NOR2_X1 U809 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U810 ( .A(KEYINPUT118), .B(n742), .Z(n743) );
  NAND2_X1 U811 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U812 ( .A(n745), .B(KEYINPUT52), .ZN(n746) );
  XNOR2_X1 U813 ( .A(n746), .B(KEYINPUT119), .ZN(n747) );
  BUF_X1 U814 ( .A(n749), .Z(n750) );
  XNOR2_X1 U815 ( .A(KEYINPUT2), .B(KEYINPUT80), .ZN(n753) );
  NAND2_X1 U816 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U817 ( .A(n758), .B(n757), .ZN(G75) );
  NAND2_X1 U818 ( .A1(n765), .A2(G469), .ZN(n763) );
  XOR2_X1 U819 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n760) );
  XNOR2_X1 U820 ( .A(n761), .B(n760), .ZN(n762) );
  XNOR2_X1 U821 ( .A(n763), .B(n762), .ZN(n764) );
  NOR2_X1 U822 ( .A1(n764), .A2(n777), .ZN(G54) );
  XOR2_X1 U823 ( .A(n766), .B(KEYINPUT59), .Z(n767) );
  NOR2_X1 U824 ( .A1(n450), .A2(n769), .ZN(n771) );
  XNOR2_X1 U825 ( .A(n771), .B(n770), .ZN(n772) );
  NOR2_X1 U826 ( .A1(n772), .A2(n777), .ZN(G63) );
  NAND2_X1 U827 ( .A1(n765), .A2(G217), .ZN(n775) );
  XOR2_X1 U828 ( .A(n773), .B(KEYINPUT121), .Z(n774) );
  XNOR2_X1 U829 ( .A(n775), .B(n774), .ZN(n776) );
  NOR2_X1 U830 ( .A1(n777), .A2(n776), .ZN(G66) );
  NAND2_X1 U831 ( .A1(G953), .A2(G224), .ZN(n778) );
  XOR2_X1 U832 ( .A(KEYINPUT61), .B(n778), .Z(n779) );
  NOR2_X1 U833 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U834 ( .A1(n377), .A2(n781), .ZN(n787) );
  XOR2_X1 U835 ( .A(n783), .B(n782), .Z(n785) );
  NAND2_X1 U836 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U837 ( .A(n787), .B(n786), .ZN(G69) );
  XOR2_X1 U838 ( .A(n413), .B(n789), .Z(n790) );
  XOR2_X1 U839 ( .A(KEYINPUT122), .B(n790), .Z(n793) );
  XNOR2_X1 U840 ( .A(n793), .B(n791), .ZN(n792) );
  NAND2_X1 U841 ( .A1(n792), .A2(n795), .ZN(n798) );
  XOR2_X1 U842 ( .A(G227), .B(n793), .Z(n794) );
  NOR2_X1 U843 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U844 ( .A1(G900), .A2(n796), .ZN(n797) );
  NAND2_X1 U845 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U846 ( .A(KEYINPUT123), .B(n799), .ZN(G72) );
  XOR2_X1 U847 ( .A(n801), .B(G122), .Z(G24) );
  XNOR2_X1 U848 ( .A(KEYINPUT126), .B(n802), .ZN(G33) );
  XNOR2_X1 U849 ( .A(G137), .B(KEYINPUT125), .ZN(n804) );
  XNOR2_X1 U850 ( .A(n804), .B(n352), .ZN(G39) );
  XNOR2_X1 U851 ( .A(n357), .B(G101), .ZN(G3) );
endmodule

