//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1023,
    new_n1024, new_n1025, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1061, new_n1062, new_n1063;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT11), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G197gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(KEYINPUT12), .ZN(new_n208));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(KEYINPUT92), .A2(G1gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT16), .ZN(new_n211));
  AND2_X1   g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(G1gat), .B1(new_n209), .B2(KEYINPUT92), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT93), .ZN(new_n214));
  OAI22_X1  g013(.A1(new_n212), .A2(new_n213), .B1(new_n214), .B2(G8gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(G8gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n215), .B(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT14), .ZN(new_n219));
  INV_X1    g018(.A(G29gat), .ZN(new_n220));
  INV_X1    g019(.A(G36gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G29gat), .A2(G36gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT15), .ZN(new_n227));
  OR2_X1    g026(.A1(G43gat), .A2(G50gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(G43gat), .A2(G50gat), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n222), .A2(KEYINPUT89), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT89), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n223), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n232), .B1(new_n222), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G43gat), .B(G50gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT15), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n225), .B(KEYINPUT90), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n228), .A2(new_n227), .A3(new_n229), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n231), .B1(new_n235), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT17), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT17), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n241), .A2(KEYINPUT91), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT91), .B1(new_n241), .B2(new_n244), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n218), .B(new_n243), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT94), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n241), .A2(new_n244), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT91), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n241), .A2(KEYINPUT91), .A3(new_n244), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT94), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n253), .A2(new_n254), .A3(new_n218), .A4(new_n243), .ZN(new_n255));
  NAND2_X1  g054(.A1(G229gat), .A2(G233gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n215), .B(new_n216), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(new_n241), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n248), .A2(new_n255), .A3(new_n256), .A4(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT95), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT18), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n258), .A2(KEYINPUT96), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n218), .A2(new_n242), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT96), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n265), .B1(new_n266), .B2(new_n264), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n256), .B(KEYINPUT13), .Z(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n261), .B1(new_n259), .B2(new_n260), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n208), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n259), .A2(new_n260), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT18), .ZN(new_n274));
  INV_X1    g073(.A(new_n208), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n274), .A2(new_n262), .A3(new_n269), .A4(new_n275), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT80), .ZN(new_n278));
  NAND2_X1  g077(.A1(G225gat), .A2(G233gat), .ZN(new_n279));
  INV_X1    g078(.A(G141gat), .ZN(new_n280));
  INV_X1    g079(.A(G148gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT2), .ZN(new_n283));
  NAND2_X1  g082(.A1(G141gat), .A2(G148gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G162gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G155gat), .ZN(new_n287));
  INV_X1    g086(.A(G155gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G162gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  XOR2_X1   g090(.A(KEYINPUT78), .B(KEYINPUT3), .Z(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT77), .B(G162gat), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n283), .B1(new_n293), .B2(G155gat), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n282), .A2(new_n287), .A3(new_n289), .A4(new_n284), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n291), .B(new_n292), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G134gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G127gat), .ZN(new_n298));
  INV_X1    g097(.A(G127gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G134gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G113gat), .B(G120gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n301), .B1(new_n302), .B2(KEYINPUT1), .ZN(new_n303));
  INV_X1    g102(.A(G113gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G120gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(KEYINPUT68), .A2(G120gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(KEYINPUT68), .A2(G120gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n306), .B1(new_n309), .B2(G113gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT1), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n298), .A2(new_n300), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n303), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  AND2_X1   g112(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n315));
  OAI21_X1  g114(.A(G155gat), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT2), .ZN(new_n317));
  AND4_X1   g116(.A1(new_n282), .A2(new_n287), .A3(new_n289), .A4(new_n284), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n317), .A2(new_n318), .B1(new_n285), .B2(new_n290), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n296), .B(new_n313), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT4), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n291), .B1(new_n294), .B2(new_n295), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n322), .B1(new_n313), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n308), .ZN(new_n325));
  NAND2_X1  g124(.A1(KEYINPUT68), .A2(G120gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(G113gat), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n305), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n298), .A2(new_n300), .A3(new_n311), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n304), .A2(G120gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n311), .B1(new_n306), .B2(new_n330), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n328), .A2(new_n329), .B1(new_n331), .B2(new_n301), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n332), .A2(new_n319), .A3(KEYINPUT4), .ZN(new_n333));
  AND4_X1   g132(.A1(new_n279), .A2(new_n321), .A3(new_n324), .A4(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT5), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n278), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n279), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n313), .A2(new_n323), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n317), .A2(new_n318), .ZN(new_n339));
  NOR3_X1   g138(.A1(new_n307), .A2(new_n308), .A3(new_n304), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n329), .B1(new_n340), .B2(new_n306), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n291), .A2(new_n339), .B1(new_n341), .B2(new_n303), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n337), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n321), .A2(new_n324), .A3(new_n279), .A4(new_n333), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n313), .A2(new_n323), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n339), .A2(new_n341), .A3(new_n291), .A4(new_n303), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n279), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT79), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n345), .A2(KEYINPUT5), .A3(new_n346), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT80), .B1(new_n346), .B2(KEYINPUT5), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n335), .B1(new_n343), .B2(new_n344), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n353), .A2(new_n346), .A3(new_n350), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  XOR2_X1   g155(.A(G1gat), .B(G29gat), .Z(new_n357));
  XNOR2_X1  g156(.A(new_n357), .B(KEYINPUT0), .ZN(new_n358));
  XNOR2_X1  g157(.A(G57gat), .B(G85gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT6), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT81), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n360), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n364), .B1(new_n352), .B2(new_n355), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT81), .B1(new_n365), .B2(KEYINPUT6), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT82), .B1(new_n356), .B2(new_n360), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT82), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n352), .A2(new_n355), .A3(new_n368), .A4(new_n364), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n363), .A2(new_n366), .A3(new_n367), .A4(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n356), .A2(new_n360), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT6), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G8gat), .B(G36gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(G64gat), .B(G92gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G183gat), .A2(G190gat), .ZN(new_n378));
  INV_X1    g177(.A(G176gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n204), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT67), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT26), .ZN(new_n382));
  NAND2_X1  g181(.A1(G169gat), .A2(G176gat), .ZN(new_n383));
  OR3_X1    g182(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT67), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n378), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G190gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT64), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT64), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(G190gat), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT28), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT27), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT27), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(KEYINPUT65), .A3(G183gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT64), .B(G190gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT27), .B(G183gat), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n395), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n402), .A2(new_n405), .A3(KEYINPUT66), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT66), .ZN(new_n407));
  INV_X1    g206(.A(G183gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT27), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n399), .A2(G183gat), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n392), .A2(new_n394), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT28), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n403), .A2(new_n395), .A3(new_n398), .A4(new_n400), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n407), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n390), .B1(new_n406), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT23), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n416), .A2(G169gat), .A3(G176gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n383), .A2(KEYINPUT23), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n417), .B1(new_n380), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(G183gat), .A2(G190gat), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT24), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n378), .B(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n419), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT25), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI211_X1 g224(.A(new_n424), .B(new_n417), .C1(new_n380), .C2(new_n418), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n403), .A2(new_n408), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n378), .B(KEYINPUT24), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(G226gat), .ZN(new_n432));
  INV_X1    g231(.A(G233gat), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n415), .A2(new_n431), .A3(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(KEYINPUT29), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT66), .B1(new_n402), .B2(new_n405), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n412), .A2(new_n407), .A3(new_n413), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n389), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n424), .A2(new_n423), .B1(new_n426), .B2(new_n429), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n436), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(G211gat), .B(G218gat), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT73), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(G211gat), .A2(G218gat), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(G211gat), .A2(G218gat), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(KEYINPUT73), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(G197gat), .B(G204gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT72), .B(KEYINPUT22), .ZN(new_n451));
  AND2_X1   g250(.A1(G211gat), .A2(G218gat), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n442), .B(new_n450), .C1(new_n451), .C2(new_n452), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT74), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n449), .A2(new_n456), .A3(new_n453), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n435), .A2(new_n441), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n460), .B1(new_n435), .B2(new_n441), .ZN(new_n462));
  OAI211_X1 g261(.A(KEYINPUT30), .B(new_n377), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n460), .ZN(new_n464));
  INV_X1    g263(.A(new_n436), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n465), .B1(new_n415), .B2(new_n431), .ZN(new_n466));
  INV_X1    g265(.A(new_n434), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n439), .A2(new_n440), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n464), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n435), .A2(new_n441), .A3(new_n460), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(new_n376), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n463), .A2(new_n471), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n472), .A2(KEYINPUT75), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n376), .B1(new_n469), .B2(new_n470), .ZN(new_n474));
  XOR2_X1   g273(.A(KEYINPUT76), .B(KEYINPUT30), .Z(new_n475));
  OR2_X1    g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n472), .A2(KEYINPUT75), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n473), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n373), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(G78gat), .B(G106gat), .ZN(new_n481));
  XOR2_X1   g280(.A(new_n481), .B(KEYINPUT83), .Z(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G228gat), .A2(G233gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(KEYINPUT84), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT22), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT72), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT72), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT22), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n452), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n452), .A2(new_n445), .ZN(new_n491));
  INV_X1    g290(.A(G204gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(G197gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n206), .A2(G204gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n490), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n453), .A2(new_n491), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT85), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n453), .A2(KEYINPUT85), .A3(new_n491), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT29), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n292), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n323), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT29), .B1(new_n319), .B2(new_n292), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n460), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n485), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n484), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n507), .B1(new_n460), .B2(new_n504), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT29), .ZN(new_n509));
  INV_X1    g308(.A(new_n459), .ZN(new_n510));
  AOI22_X1  g309(.A1(new_n449), .A2(new_n453), .B1(new_n455), .B2(new_n456), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(new_n320), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n508), .B1(new_n513), .B2(new_n323), .ZN(new_n514));
  OAI21_X1  g313(.A(G22gat), .B1(new_n506), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n485), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n497), .A2(new_n498), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(new_n500), .A3(new_n455), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n509), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n319), .B1(new_n519), .B2(new_n292), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n460), .A2(new_n504), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n516), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(G22gat), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT3), .B1(new_n460), .B2(new_n509), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n505), .B(new_n507), .C1(new_n524), .C2(new_n319), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  XOR2_X1   g325(.A(KEYINPUT31), .B(G50gat), .Z(new_n527));
  AND3_X1   g326(.A1(new_n515), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n527), .B1(new_n515), .B2(new_n526), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n483), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n527), .ZN(new_n531));
  NOR3_X1   g330(.A1(new_n506), .A2(new_n514), .A3(G22gat), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n523), .B1(new_n522), .B2(new_n525), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n515), .A2(new_n526), .A3(new_n527), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(new_n482), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT86), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n530), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n537), .B1(new_n530), .B2(new_n536), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n480), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n415), .A2(new_n313), .A3(new_n431), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n332), .B1(new_n439), .B2(new_n440), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G227gat), .A2(G233gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT70), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT34), .ZN(new_n547));
  OAI211_X1 g346(.A(new_n544), .B(new_n545), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n545), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n542), .A2(new_n543), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT32), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT69), .B(KEYINPUT33), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(G15gat), .B(G43gat), .Z(new_n554));
  XNOR2_X1  g353(.A(G71gat), .B(G99gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n551), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n544), .A2(new_n545), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n547), .B1(new_n545), .B2(new_n546), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n556), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n550), .B(KEYINPUT32), .C1(new_n552), .C2(new_n561), .ZN(new_n562));
  AND4_X1   g361(.A1(new_n548), .A2(new_n557), .A3(new_n560), .A4(new_n562), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n557), .A2(new_n562), .B1(new_n548), .B2(new_n560), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(KEYINPUT71), .A2(KEYINPUT36), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(KEYINPUT71), .B(KEYINPUT36), .Z(new_n568));
  AOI21_X1  g367(.A(new_n567), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT87), .ZN(new_n570));
  AND3_X1   g369(.A1(new_n352), .A2(new_n570), .A3(new_n355), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n570), .B1(new_n352), .B2(new_n355), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n364), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(new_n361), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT37), .B1(new_n461), .B2(new_n462), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT37), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n469), .A2(new_n576), .A3(new_n470), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT38), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n377), .B1(new_n461), .B2(new_n462), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n578), .A2(new_n376), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI211_X1 g380(.A(KEYINPUT38), .B(new_n377), .C1(new_n575), .C2(new_n577), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n574), .A2(new_n372), .A3(new_n583), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n463), .B(new_n471), .C1(new_n474), .C2(new_n475), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n321), .A2(new_n324), .A3(new_n333), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(new_n337), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n347), .A2(new_n348), .A3(new_n279), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n588), .A2(KEYINPUT39), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n364), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT39), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n586), .A2(new_n591), .A3(new_n337), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n590), .A2(KEYINPUT40), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT40), .B1(new_n590), .B2(new_n592), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n573), .A2(new_n585), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(new_n536), .A3(new_n530), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT88), .B1(new_n584), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n530), .A2(new_n536), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n336), .A2(new_n351), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT5), .B1(new_n349), .B2(KEYINPUT79), .ZN(new_n601));
  AOI211_X1 g400(.A(new_n344), .B(new_n279), .C1(new_n347), .C2(new_n348), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n353), .B1(new_n603), .B2(new_n346), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT87), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n352), .A2(new_n570), .A3(new_n355), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n360), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n585), .A2(new_n595), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n599), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT88), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n574), .A2(new_n372), .A3(new_n583), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n541), .A2(new_n569), .A3(new_n598), .A4(new_n613), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n565), .A2(new_n536), .A3(new_n530), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n373), .A2(new_n615), .A3(new_n479), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT35), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n565), .A2(new_n530), .A3(new_n536), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n573), .A2(new_n361), .B1(KEYINPUT6), .B2(new_n371), .ZN(new_n619));
  INV_X1    g418(.A(new_n585), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT35), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR3_X1   g421(.A1(new_n618), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n617), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n277), .B1(new_n614), .B2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G127gat), .B(G155gat), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n627), .B(KEYINPUT20), .Z(new_n628));
  XOR2_X1   g427(.A(G71gat), .B(G78gat), .Z(new_n629));
  XNOR2_X1  g428(.A(G57gat), .B(G64gat), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT9), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT97), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(G57gat), .B(G64gat), .Z(new_n636));
  XNOR2_X1  g435(.A(G71gat), .B(G78gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n632), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT21), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G231gat), .A2(G233gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT98), .B(KEYINPUT19), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n642), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n641), .B(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n644), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n628), .B1(new_n645), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n645), .A2(new_n649), .A3(new_n628), .ZN(new_n652));
  XOR2_X1   g451(.A(G183gat), .B(G211gat), .Z(new_n653));
  NAND3_X1  g452(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n653), .ZN(new_n655));
  INV_X1    g454(.A(new_n652), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n655), .B1(new_n656), .B2(new_n650), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n637), .B1(new_n636), .B2(KEYINPUT9), .ZN(new_n658));
  INV_X1    g457(.A(new_n635), .ZN(new_n659));
  INV_X1    g458(.A(new_n638), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n257), .B1(KEYINPUT21), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT99), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n654), .A2(new_n657), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n663), .B1(new_n654), .B2(new_n657), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(G99gat), .A2(G106gat), .ZN(new_n668));
  INV_X1    g467(.A(G85gat), .ZN(new_n669));
  INV_X1    g468(.A(G92gat), .ZN(new_n670));
  AOI22_X1  g469(.A1(KEYINPUT8), .A2(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT7), .ZN(new_n672));
  OAI22_X1  g471(.A1(new_n669), .A2(new_n670), .B1(new_n672), .B2(KEYINPUT101), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT101), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n674), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n671), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g475(.A(G99gat), .B(G106gat), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n243), .B(new_n678), .C1(new_n245), .C2(new_n246), .ZN(new_n679));
  INV_X1    g478(.A(new_n677), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n676), .B(new_n680), .ZN(new_n681));
  AND2_X1   g480(.A1(G232gat), .A2(G233gat), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n681), .A2(new_n241), .B1(KEYINPUT41), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(G190gat), .B(G218gat), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n685), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n687), .B1(new_n679), .B2(new_n683), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n682), .A2(KEYINPUT41), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT100), .ZN(new_n691));
  XOR2_X1   g490(.A(G134gat), .B(G162gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(new_n688), .B2(KEYINPUT102), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n689), .A2(new_n694), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(G120gat), .B(G148gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(G176gat), .B(G204gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n676), .A2(KEYINPUT103), .A3(new_n677), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n677), .B1(new_n676), .B2(KEYINPUT103), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n661), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n681), .A2(new_n639), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(G230gat), .A2(G233gat), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT10), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n678), .A2(new_n661), .ZN(new_n711));
  INV_X1    g510(.A(new_n704), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n639), .B1(new_n712), .B2(new_n702), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n710), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n678), .A2(new_n710), .A3(new_n639), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  AOI211_X1 g516(.A(new_n701), .B(new_n709), .C1(new_n717), .C2(new_n708), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n708), .B(KEYINPUT104), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n720), .B1(new_n714), .B2(new_n716), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n701), .B1(new_n721), .B2(new_n709), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n626), .A2(new_n667), .A3(new_n698), .A4(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n373), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g528(.A1(new_n725), .A2(new_n620), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT16), .B(G8gat), .Z(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(KEYINPUT105), .A3(KEYINPUT42), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT105), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT42), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n732), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n730), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n736), .B1(new_n738), .B2(G8gat), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n734), .B(new_n737), .C1(new_n733), .C2(new_n739), .ZN(G1325gat));
  OAI21_X1  g539(.A(G15gat), .B1(new_n725), .B2(new_n569), .ZN(new_n741));
  INV_X1    g540(.A(new_n565), .ZN(new_n742));
  OR2_X1    g541(.A1(new_n742), .A2(G15gat), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n725), .B2(new_n743), .ZN(G1326gat));
  NAND2_X1  g543(.A1(new_n599), .A2(KEYINPUT86), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n530), .A2(new_n536), .A3(new_n537), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n725), .A2(new_n747), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT43), .B(G22gat), .Z(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1327gat));
  INV_X1    g549(.A(new_n698), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n666), .A2(new_n751), .A3(new_n724), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT106), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n626), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n754), .A2(new_n220), .A3(new_n727), .ZN(new_n755));
  XOR2_X1   g554(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n623), .B1(new_n616), .B2(KEYINPUT35), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n530), .A2(new_n536), .ZN(new_n760));
  AND4_X1   g559(.A1(new_n611), .A2(new_n612), .A3(new_n760), .A4(new_n596), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n611), .B1(new_n610), .B2(new_n612), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n565), .A2(new_n568), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n565), .B2(new_n566), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n765), .B1(new_n480), .B2(new_n540), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n759), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT108), .B1(new_n696), .B2(new_n697), .ZN(new_n768));
  INV_X1    g567(.A(new_n697), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT108), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n769), .A2(new_n770), .A3(new_n695), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n758), .B1(new_n767), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n598), .A2(new_n613), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n478), .B1(new_n370), .B2(new_n372), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n569), .B1(new_n747), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n621), .B1(new_n775), .B2(new_n615), .ZN(new_n777));
  OAI22_X1  g576(.A1(new_n774), .A2(new_n776), .B1(new_n777), .B2(new_n623), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n778), .A2(KEYINPUT44), .A3(new_n751), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n773), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n666), .A2(new_n724), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n277), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(G29gat), .B1(new_n783), .B2(new_n373), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n757), .A2(new_n784), .ZN(G1328gat));
  NAND3_X1  g584(.A1(new_n754), .A2(new_n221), .A3(new_n585), .ZN(new_n786));
  XOR2_X1   g585(.A(new_n786), .B(KEYINPUT46), .Z(new_n787));
  OAI21_X1  g586(.A(G36gat), .B1(new_n783), .B2(new_n620), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(G1329gat));
  NAND4_X1  g588(.A1(new_n773), .A2(new_n765), .A3(new_n779), .A4(new_n782), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G43gat), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n272), .A2(new_n276), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n742), .A2(G43gat), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n778), .A2(new_n792), .A3(new_n753), .A4(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n791), .A2(KEYINPUT47), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n626), .A2(KEYINPUT109), .A3(new_n753), .A4(new_n793), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n791), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT110), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT110), .ZN(new_n803));
  AOI211_X1 g602(.A(new_n803), .B(KEYINPUT47), .C1(new_n791), .C2(new_n799), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n795), .B1(new_n802), .B2(new_n804), .ZN(G1330gat));
  NAND3_X1  g604(.A1(new_n780), .A2(new_n540), .A3(new_n782), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n747), .A2(G50gat), .ZN(new_n807));
  AOI22_X1  g606(.A1(new_n806), .A2(G50gat), .B1(new_n754), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n773), .A2(new_n599), .A3(new_n779), .A4(new_n782), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G50gat), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT48), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n754), .B2(new_n807), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n810), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(new_n810), .B2(new_n812), .ZN(new_n815));
  OAI22_X1  g614(.A1(new_n808), .A2(KEYINPUT48), .B1(new_n814), .B2(new_n815), .ZN(G1331gat));
  NAND2_X1  g615(.A1(new_n667), .A2(new_n698), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n817), .A2(new_n792), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n723), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n767), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n727), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g621(.A1(new_n820), .A2(KEYINPUT112), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n824), .B1(new_n767), .B2(new_n819), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n620), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n823), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n828));
  XOR2_X1   g627(.A(new_n827), .B(new_n828), .Z(G1333gat));
  NAND2_X1  g628(.A1(new_n823), .A2(new_n825), .ZN(new_n830));
  OAI21_X1  g629(.A(G71gat), .B1(new_n830), .B2(new_n569), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT50), .ZN(new_n832));
  INV_X1    g631(.A(G71gat), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n820), .A2(KEYINPUT113), .A3(new_n565), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT113), .B1(new_n820), .B2(new_n565), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n831), .A2(new_n832), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n832), .B1(new_n831), .B2(new_n836), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n837), .A2(new_n838), .ZN(G1334gat));
  NOR2_X1   g638(.A1(new_n830), .A2(new_n747), .ZN(new_n840));
  XOR2_X1   g639(.A(KEYINPUT114), .B(G78gat), .Z(new_n841));
  XNOR2_X1  g640(.A(new_n840), .B(new_n841), .ZN(G1335gat));
  NOR2_X1   g641(.A1(new_n667), .A2(new_n792), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n778), .A2(new_n751), .A3(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n778), .A2(KEYINPUT51), .A3(new_n751), .A4(new_n843), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n724), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(new_n669), .A3(new_n727), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n667), .A2(new_n792), .A3(new_n724), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n780), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n850), .B1(new_n852), .B2(new_n373), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(G85gat), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n852), .A2(new_n850), .A3(new_n373), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n849), .B1(new_n854), .B2(new_n855), .ZN(G1336gat));
  NOR2_X1   g655(.A1(new_n620), .A2(new_n670), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n780), .A2(new_n851), .A3(new_n857), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n848), .A2(new_n585), .ZN(new_n859));
  OAI211_X1 g658(.A(KEYINPUT52), .B(new_n858), .C1(new_n859), .C2(G92gat), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n861));
  INV_X1    g660(.A(new_n858), .ZN(new_n862));
  AOI21_X1  g661(.A(G92gat), .B1(new_n848), .B2(new_n585), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n860), .A2(new_n864), .ZN(G1337gat));
  INV_X1    g664(.A(G99gat), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n848), .A2(new_n866), .A3(new_n565), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n868), .B1(new_n852), .B2(new_n569), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(G99gat), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n852), .A2(new_n868), .A3(new_n569), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n867), .B1(new_n870), .B2(new_n871), .ZN(G1338gat));
  OAI21_X1  g671(.A(G106gat), .B1(new_n852), .B2(new_n760), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n846), .A2(new_n847), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n760), .A2(G106gat), .A3(new_n724), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT53), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n780), .A2(new_n540), .A3(new_n851), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n875), .B(KEYINPUT117), .ZN(new_n879));
  AOI22_X1  g678(.A1(new_n878), .A2(G106gat), .B1(new_n874), .B2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n877), .B1(new_n880), .B2(new_n881), .ZN(G1339gat));
  NAND2_X1  g681(.A1(new_n818), .A2(new_n724), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT10), .B1(new_n705), .B2(new_n706), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n708), .B1(new_n884), .B2(new_n715), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n714), .A2(new_n716), .A3(new_n720), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT54), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT118), .A4(KEYINPUT54), .ZN(new_n890));
  INV_X1    g689(.A(new_n701), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(new_n721), .B2(new_n892), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n889), .A2(KEYINPUT55), .A3(new_n890), .A4(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n893), .A2(new_n890), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n897), .A2(KEYINPUT119), .A3(KEYINPUT55), .A4(new_n889), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n889), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT55), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n718), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n248), .A2(new_n255), .A3(new_n258), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(G229gat), .A3(G233gat), .ZN(new_n904));
  INV_X1    g703(.A(new_n268), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n265), .B(new_n905), .C1(new_n266), .C2(new_n264), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n207), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n899), .A2(new_n902), .A3(new_n276), .A4(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(new_n772), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n276), .A2(new_n908), .A3(new_n723), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n899), .A2(new_n902), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n277), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n910), .B1(new_n913), .B2(new_n772), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n883), .B1(new_n914), .B2(new_n667), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n373), .A2(new_n585), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n917), .A2(new_n618), .ZN(new_n918));
  AOI21_X1  g717(.A(G113gat), .B1(new_n918), .B2(new_n792), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n540), .A2(new_n742), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n277), .A2(new_n304), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(G1340gat));
  INV_X1    g723(.A(new_n922), .ZN(new_n925));
  OAI21_X1  g724(.A(G120gat), .B1(new_n925), .B2(new_n724), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n918), .A2(new_n309), .A3(new_n723), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1341gat));
  OAI21_X1  g727(.A(G127gat), .B1(new_n925), .B2(new_n666), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n918), .A2(new_n299), .A3(new_n667), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1342gat));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n751), .A3(new_n916), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n932), .A2(G134gat), .A3(new_n618), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT56), .ZN(new_n934));
  OAI21_X1  g733(.A(G134gat), .B1(new_n932), .B2(new_n921), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1343gat));
  NOR3_X1   g735(.A1(new_n817), .A2(new_n792), .A3(new_n723), .ZN(new_n937));
  INV_X1    g736(.A(new_n909), .ZN(new_n938));
  INV_X1    g737(.A(new_n772), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n893), .A2(new_n890), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n892), .B1(new_n717), .B2(new_n708), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT118), .B1(new_n942), .B2(new_n886), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n901), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n719), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n945), .B1(new_n896), .B2(new_n898), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n270), .A2(new_n271), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n907), .B1(new_n947), .B2(new_n275), .ZN(new_n948));
  AOI22_X1  g747(.A1(new_n792), .A2(new_n946), .B1(new_n948), .B2(new_n723), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n940), .B1(new_n949), .B2(new_n751), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n937), .B1(new_n950), .B2(new_n666), .ZN(new_n951));
  OAI21_X1  g750(.A(KEYINPUT57), .B1(new_n951), .B2(new_n747), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT57), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n915), .A2(new_n953), .A3(new_n599), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n765), .A2(new_n373), .A3(new_n585), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n952), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n956), .A2(G141gat), .A3(new_n792), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n569), .A2(new_n599), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n917), .A2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n280), .B1(new_n960), .B2(new_n277), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n957), .A2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT58), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n957), .A2(new_n961), .A3(KEYINPUT58), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1344gat));
  NAND4_X1  g765(.A1(new_n952), .A2(new_n723), .A3(new_n954), .A4(new_n955), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT59), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n915), .A2(new_n599), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(KEYINPUT57), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n913), .A2(new_n698), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n938), .A2(new_n751), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(new_n666), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(new_n883), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n540), .A2(new_n953), .ZN(new_n977));
  INV_X1    g776(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  XOR2_X1   g778(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n980));
  OR2_X1    g779(.A1(new_n955), .A2(KEYINPUT121), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n955), .A2(KEYINPUT121), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND4_X1  g782(.A1(new_n971), .A2(new_n979), .A3(new_n723), .A4(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n281), .B1(new_n969), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n980), .A2(G148gat), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n986), .B1(new_n960), .B2(new_n724), .ZN(new_n987));
  INV_X1    g786(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g787(.A(KEYINPUT122), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT122), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n953), .B1(new_n915), .B2(new_n599), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n977), .B1(new_n975), .B2(new_n883), .ZN(new_n992));
  NOR3_X1   g791(.A1(new_n991), .A2(new_n992), .A3(new_n724), .ZN(new_n993));
  AOI22_X1  g792(.A1(new_n993), .A2(new_n983), .B1(new_n967), .B2(new_n968), .ZN(new_n994));
  OAI211_X1 g793(.A(new_n990), .B(new_n987), .C1(new_n994), .C2(new_n281), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n989), .A2(new_n995), .ZN(G1345gat));
  NAND3_X1  g795(.A1(new_n959), .A2(new_n288), .A3(new_n667), .ZN(new_n997));
  AND2_X1   g796(.A1(new_n956), .A2(new_n667), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n997), .B1(new_n998), .B2(new_n288), .ZN(G1346gat));
  NAND3_X1  g798(.A1(new_n956), .A2(new_n293), .A3(new_n939), .ZN(new_n1000));
  INV_X1    g799(.A(new_n293), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n1001), .B1(new_n932), .B2(new_n958), .ZN(new_n1002));
  AND2_X1   g801(.A1(new_n1000), .A2(new_n1002), .ZN(G1347gat));
  AND2_X1   g802(.A1(new_n915), .A2(new_n373), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n618), .A2(new_n620), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g805(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g806(.A(G169gat), .B1(new_n1007), .B2(new_n792), .ZN(new_n1008));
  NOR2_X1   g807(.A1(new_n727), .A2(new_n620), .ZN(new_n1009));
  AND3_X1   g808(.A1(new_n915), .A2(new_n920), .A3(new_n1009), .ZN(new_n1010));
  NOR2_X1   g809(.A1(new_n277), .A2(new_n204), .ZN(new_n1011));
  AOI21_X1  g810(.A(new_n1008), .B1(new_n1010), .B2(new_n1011), .ZN(G1348gat));
  NAND3_X1  g811(.A1(new_n1007), .A2(new_n379), .A3(new_n723), .ZN(new_n1013));
  AND2_X1   g812(.A1(new_n1010), .A2(new_n723), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1013), .B1(new_n379), .B2(new_n1014), .ZN(G1349gat));
  NAND2_X1  g814(.A1(new_n667), .A2(new_n404), .ZN(new_n1016));
  INV_X1    g815(.A(KEYINPUT60), .ZN(new_n1017));
  OAI22_X1  g816(.A1(new_n1006), .A2(new_n1016), .B1(KEYINPUT123), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g817(.A(new_n408), .B1(new_n1010), .B2(new_n667), .ZN(new_n1019));
  NOR2_X1   g818(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AND2_X1   g819(.A1(new_n1017), .A2(KEYINPUT123), .ZN(new_n1021));
  XNOR2_X1  g820(.A(new_n1020), .B(new_n1021), .ZN(G1350gat));
  AOI21_X1  g821(.A(new_n391), .B1(new_n1010), .B2(new_n751), .ZN(new_n1023));
  XOR2_X1   g822(.A(new_n1023), .B(KEYINPUT61), .Z(new_n1024));
  NAND3_X1  g823(.A1(new_n1007), .A2(new_n403), .A3(new_n939), .ZN(new_n1025));
  NAND2_X1  g824(.A1(new_n1024), .A2(new_n1025), .ZN(G1351gat));
  NOR2_X1   g825(.A1(new_n958), .A2(new_n620), .ZN(new_n1027));
  XNOR2_X1  g826(.A(new_n1027), .B(KEYINPUT124), .ZN(new_n1028));
  NAND2_X1  g827(.A1(new_n1004), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1029), .A2(KEYINPUT125), .ZN(new_n1030));
  INV_X1    g829(.A(KEYINPUT125), .ZN(new_n1031));
  NAND3_X1  g830(.A1(new_n1004), .A2(new_n1031), .A3(new_n1028), .ZN(new_n1032));
  AND2_X1   g831(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g832(.A1(new_n1033), .A2(new_n206), .A3(new_n792), .ZN(new_n1034));
  NAND2_X1  g833(.A1(new_n971), .A2(new_n979), .ZN(new_n1035));
  NAND2_X1  g834(.A1(new_n1009), .A2(new_n569), .ZN(new_n1036));
  OR2_X1    g835(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g836(.A(G197gat), .B1(new_n1037), .B2(new_n277), .ZN(new_n1038));
  NAND2_X1  g837(.A1(new_n1034), .A2(new_n1038), .ZN(G1352gat));
  INV_X1    g838(.A(KEYINPUT126), .ZN(new_n1040));
  NOR2_X1   g839(.A1(new_n724), .A2(G204gat), .ZN(new_n1041));
  INV_X1    g840(.A(new_n1041), .ZN(new_n1042));
  OAI21_X1  g841(.A(new_n1040), .B1(new_n1029), .B2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g842(.A1(new_n1004), .A2(new_n1028), .A3(KEYINPUT126), .A4(new_n1041), .ZN(new_n1044));
  AND3_X1   g843(.A1(new_n1043), .A2(KEYINPUT62), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g844(.A(KEYINPUT62), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1046));
  NOR3_X1   g845(.A1(new_n1035), .A2(new_n724), .A3(new_n1036), .ZN(new_n1047));
  OAI22_X1  g846(.A1(new_n1045), .A2(new_n1046), .B1(new_n492), .B2(new_n1047), .ZN(G1353gat));
  NOR2_X1   g847(.A1(new_n666), .A2(G211gat), .ZN(new_n1049));
  NAND3_X1  g848(.A1(new_n1030), .A2(new_n1032), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g849(.A1(new_n1050), .A2(KEYINPUT127), .ZN(new_n1051));
  INV_X1    g850(.A(KEYINPUT127), .ZN(new_n1052));
  NAND4_X1  g851(.A1(new_n1030), .A2(new_n1052), .A3(new_n1032), .A4(new_n1049), .ZN(new_n1053));
  NAND2_X1  g852(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g853(.A(KEYINPUT63), .ZN(new_n1055));
  OAI211_X1 g854(.A(new_n1055), .B(G211gat), .C1(new_n1037), .C2(new_n666), .ZN(new_n1056));
  NOR3_X1   g855(.A1(new_n1035), .A2(new_n666), .A3(new_n1036), .ZN(new_n1057));
  INV_X1    g856(.A(G211gat), .ZN(new_n1058));
  OAI21_X1  g857(.A(KEYINPUT63), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g858(.A1(new_n1054), .A2(new_n1056), .A3(new_n1059), .ZN(G1354gat));
  INV_X1    g859(.A(G218gat), .ZN(new_n1061));
  NAND3_X1  g860(.A1(new_n1033), .A2(new_n1061), .A3(new_n939), .ZN(new_n1062));
  OAI21_X1  g861(.A(G218gat), .B1(new_n1037), .B2(new_n698), .ZN(new_n1063));
  NAND2_X1  g862(.A1(new_n1062), .A2(new_n1063), .ZN(G1355gat));
endmodule


