//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n191), .A3(new_n195), .A4(new_n192), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(KEYINPUT64), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n193), .A2(new_n198), .A3(G131), .ZN(new_n199));
  XNOR2_X1  g013(.A(G143), .B(G146), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT0), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n200), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  XOR2_X1   g017(.A(KEYINPUT0), .B(G128), .Z(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n200), .B2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n197), .A2(new_n199), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n207), .A2(G143), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n211), .A2(new_n202), .B1(KEYINPUT1), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n200), .A2(new_n214), .A3(G128), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n192), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n188), .A2(G137), .ZN(new_n218));
  OAI21_X1  g032(.A(G131), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n196), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n206), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT30), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(KEYINPUT65), .A2(G119), .ZN(new_n224));
  NOR2_X1   g038(.A1(KEYINPUT65), .A2(G119), .ZN(new_n225));
  OAI21_X1  g039(.A(G116), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G116), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G119), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT2), .B(G113), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n230), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(new_n226), .A3(new_n228), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n206), .A2(KEYINPUT30), .A3(new_n220), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n223), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT31), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n231), .A2(KEYINPUT66), .A3(new_n233), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n239), .A2(new_n206), .A3(new_n240), .A4(new_n220), .ZN(new_n241));
  NOR2_X1   g055(.A1(G237), .A2(G953), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G210), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n243), .B(G101), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n236), .A2(new_n237), .A3(new_n241), .A4(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n247), .B(KEYINPUT67), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n236), .A2(new_n241), .A3(new_n246), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT31), .ZN(new_n250));
  XOR2_X1   g064(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n221), .A2(new_n234), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(new_n241), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT28), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n241), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n250), .B1(new_n246), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT69), .B1(new_n248), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(G472), .A2(G902), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n247), .B(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n263));
  INV_X1    g077(.A(new_n257), .ZN(new_n264));
  INV_X1    g078(.A(new_n246), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n264), .A2(new_n265), .B1(new_n249), .B2(KEYINPUT31), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n262), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n259), .A2(new_n260), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT32), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n259), .A2(new_n267), .A3(KEYINPUT32), .A4(new_n260), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n264), .A2(new_n246), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n236), .A2(new_n241), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n265), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT29), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n239), .A2(new_n240), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n221), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n241), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n256), .B1(new_n278), .B2(KEYINPUT28), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(KEYINPUT29), .A3(new_n246), .ZN(new_n280));
  INV_X1    g094(.A(G902), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(G472), .B1(new_n275), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n270), .A2(new_n271), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G234), .ZN(new_n285));
  OAI21_X1  g099(.A(G217), .B1(new_n285), .B2(G902), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n286), .B(KEYINPUT70), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G140), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G125), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(KEYINPUT16), .ZN(new_n291));
  XNOR2_X1  g105(.A(G125), .B(G140), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n291), .B1(new_n292), .B2(KEYINPUT16), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G146), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT75), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n292), .A2(KEYINPUT16), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n297), .B(new_n207), .C1(new_n298), .C2(new_n291), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT75), .B1(new_n293), .B2(G146), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n293), .A2(KEYINPUT74), .A3(G146), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n296), .A2(new_n299), .A3(new_n300), .A4(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(G128), .B1(new_n224), .B2(new_n225), .ZN(new_n303));
  INV_X1    g117(.A(G119), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n303), .B1(new_n304), .B2(G128), .ZN(new_n305));
  XOR2_X1   g119(.A(KEYINPUT24), .B(G110), .Z(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OR2_X1    g121(.A1(KEYINPUT65), .A2(G119), .ZN(new_n308));
  NAND2_X1  g122(.A1(KEYINPUT65), .A2(G119), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n202), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OR2_X1    g124(.A1(KEYINPUT71), .A2(KEYINPUT23), .ZN(new_n311));
  NAND2_X1  g125(.A1(KEYINPUT71), .A2(KEYINPUT23), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT72), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  OR4_X1    g128(.A1(KEYINPUT73), .A2(new_n224), .A3(new_n225), .A4(G128), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n308), .A2(new_n309), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT73), .B1(new_n316), .B2(G128), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT72), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n303), .A2(new_n318), .A3(new_n311), .A4(new_n312), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n314), .A2(new_n315), .A3(new_n317), .A4(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n202), .A2(KEYINPUT23), .A3(G119), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G110), .ZN(new_n323));
  OAI221_X1 g137(.A(new_n302), .B1(new_n305), .B2(new_n307), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n320), .A2(new_n323), .A3(new_n321), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n305), .A2(new_n307), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n292), .A2(new_n207), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n294), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n325), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  AOI211_X1 g146(.A(KEYINPUT76), .B(new_n330), .C1(new_n326), .C2(new_n327), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n324), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT22), .B(G137), .ZN(new_n335));
  INV_X1    g149(.A(G221), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n336), .A2(new_n285), .A3(G953), .ZN(new_n337));
  XOR2_X1   g151(.A(new_n335), .B(new_n337), .Z(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n324), .B(new_n338), .C1(new_n332), .C2(new_n333), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n281), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT25), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n340), .A2(KEYINPUT25), .A3(new_n281), .A4(new_n341), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n288), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n340), .A2(new_n341), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n286), .A2(new_n281), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n346), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n284), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n284), .A2(KEYINPUT77), .A3(new_n351), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n292), .B(new_n207), .ZN(new_n356));
  INV_X1    g170(.A(G237), .ZN(new_n357));
  INV_X1    g171(.A(G953), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(G214), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n209), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n242), .A2(G143), .A3(G214), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n362), .A2(KEYINPUT88), .A3(KEYINPUT18), .A4(G131), .ZN(new_n363));
  NAND2_X1  g177(.A1(KEYINPUT18), .A2(G131), .ZN(new_n364));
  INV_X1    g178(.A(new_n362), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT88), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n365), .A2(new_n366), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n356), .B(new_n363), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT19), .B1(new_n292), .B2(KEYINPUT90), .ZN(new_n370));
  INV_X1    g184(.A(G125), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G140), .ZN(new_n372));
  AND4_X1   g186(.A1(KEYINPUT90), .A2(new_n290), .A3(new_n372), .A4(KEYINPUT19), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n207), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT91), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g190(.A(KEYINPUT91), .B(new_n207), .C1(new_n370), .C2(new_n373), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(new_n294), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n360), .A2(new_n195), .A3(new_n361), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n195), .B1(new_n360), .B2(new_n361), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT89), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n381), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT89), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(new_n379), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n369), .B1(new_n378), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(G113), .B(G122), .ZN(new_n388));
  INV_X1    g202(.A(G104), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n388), .B(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT17), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n383), .A2(new_n393), .A3(new_n379), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n394), .B1(new_n393), .B2(new_n383), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n390), .B(new_n369), .C1(new_n302), .C2(new_n395), .ZN(new_n396));
  AOI211_X1 g210(.A(G475), .B(G902), .C1(new_n392), .C2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT20), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT92), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(G475), .B1(new_n392), .B2(new_n396), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n281), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT92), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n402), .A3(KEYINPUT20), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n392), .A2(new_n396), .ZN(new_n404));
  INV_X1    g218(.A(G475), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n404), .A2(new_n398), .A3(new_n405), .A4(new_n281), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT93), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n400), .A2(KEYINPUT93), .A3(new_n398), .A4(new_n281), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n399), .A2(new_n403), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n369), .B1(new_n302), .B2(new_n395), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n411), .A2(new_n391), .ZN(new_n412));
  INV_X1    g226(.A(new_n396), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n281), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G475), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n202), .A2(G143), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n209), .A2(G128), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(KEYINPUT13), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n420), .B(G134), .C1(KEYINPUT13), .C2(new_n419), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(new_n419), .A3(new_n188), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT78), .B(G107), .ZN(new_n423));
  INV_X1    g237(.A(G122), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G116), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n227), .A2(G122), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AND2_X1   g241(.A1(KEYINPUT78), .A2(G107), .ZN(new_n428));
  NOR2_X1   g242(.A1(KEYINPUT78), .A2(G107), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n425), .B(new_n426), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n421), .B(new_n422), .C1(new_n427), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n418), .A2(new_n419), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G134), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n422), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT14), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n425), .A2(new_n426), .A3(new_n436), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n437), .B(G107), .C1(new_n436), .C2(new_n426), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n435), .A2(new_n438), .A3(new_n430), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT94), .ZN(new_n441));
  XOR2_X1   g255(.A(KEYINPUT9), .B(G234), .Z(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(G217), .A3(new_n358), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT94), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n432), .A2(new_n445), .A3(new_n439), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n441), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n444), .B1(new_n441), .B2(new_n446), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n281), .ZN(new_n450));
  INV_X1    g264(.A(G478), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n451), .A2(KEYINPUT15), .ZN(new_n452));
  XOR2_X1   g266(.A(new_n450), .B(new_n452), .Z(new_n453));
  NAND2_X1  g267(.A1(new_n417), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT85), .ZN(new_n455));
  INV_X1    g269(.A(new_n216), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n371), .ZN(new_n457));
  OR2_X1    g271(.A1(new_n205), .A2(new_n371), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n358), .A2(G224), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n459), .B(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT3), .ZN(new_n462));
  INV_X1    g276(.A(G107), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n462), .B1(new_n463), .B2(G104), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n389), .B2(G107), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n462), .B(G104), .C1(new_n428), .C2(new_n429), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G101), .ZN(new_n468));
  INV_X1    g282(.A(G101), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n465), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(KEYINPUT4), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT4), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n467), .A2(new_n472), .A3(G101), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n471), .A2(new_n234), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n226), .A2(KEYINPUT5), .A3(new_n228), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT5), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n316), .A2(new_n476), .A3(G116), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n475), .A2(G113), .A3(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n423), .A2(G104), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n389), .A2(G107), .ZN(new_n480));
  OAI21_X1  g294(.A(G101), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n478), .A2(new_n481), .A3(new_n233), .A4(new_n470), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n474), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(G110), .B(G122), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n485), .B(KEYINPUT81), .Z(new_n486));
  AOI21_X1  g300(.A(new_n486), .B1(new_n474), .B2(new_n482), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n484), .A2(new_n485), .B1(new_n487), .B2(KEYINPUT6), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n487), .A2(KEYINPUT6), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n461), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n485), .B(KEYINPUT8), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n481), .A2(new_n470), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(new_n233), .A3(new_n478), .ZN(new_n494));
  INV_X1    g308(.A(new_n233), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n477), .A2(KEYINPUT83), .A3(G113), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT83), .B1(new_n477), .B2(G113), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n475), .B(KEYINPUT82), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n492), .B(new_n494), .C1(new_n500), .C2(new_n493), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n474), .A2(new_n482), .A3(new_n485), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT84), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n460), .A2(KEYINPUT7), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n457), .B(new_n458), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n504), .B1(new_n458), .B2(new_n503), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n459), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n501), .A2(new_n502), .A3(new_n505), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n281), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n455), .B1(new_n491), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n461), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n487), .A2(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n502), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n511), .B1(new_n513), .B2(new_n489), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n514), .A2(KEYINPUT85), .A3(new_n281), .A4(new_n508), .ZN(new_n515));
  OAI21_X1  g329(.A(G210), .B1(G237), .B2(G902), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(KEYINPUT86), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n510), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT87), .ZN(new_n519));
  INV_X1    g333(.A(new_n517), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n514), .A2(new_n281), .A3(new_n520), .A4(new_n508), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n510), .A2(new_n515), .A3(KEYINPUT87), .A4(new_n517), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n358), .A2(G952), .ZN(new_n524));
  NAND2_X1  g338(.A1(G234), .A2(G237), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  XOR2_X1   g340(.A(new_n526), .B(KEYINPUT95), .Z(new_n527));
  AND3_X1   g341(.A1(new_n525), .A2(G902), .A3(G953), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT21), .B(G898), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(G214), .B1(G237), .B2(G902), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n522), .A2(new_n523), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G469), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT10), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n215), .A2(KEYINPUT79), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT79), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n200), .A2(new_n539), .A3(new_n214), .A4(G128), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(new_n213), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n537), .B1(new_n542), .B2(new_n493), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n481), .A2(new_n470), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(KEYINPUT10), .A3(new_n216), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n197), .A2(new_n199), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n471), .A2(new_n205), .A3(new_n473), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n543), .A2(new_n545), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  XOR2_X1   g362(.A(G110), .B(G140), .Z(new_n549));
  AND2_X1   g363(.A1(new_n358), .A2(G227), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n544), .A2(new_n541), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n493), .A2(new_n456), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n546), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT12), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT80), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n556), .B1(new_n546), .B2(new_n557), .ZN(new_n558));
  OR2_X1    g372(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n555), .A2(new_n558), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n552), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n543), .A2(new_n545), .A3(new_n547), .ZN(new_n562));
  INV_X1    g376(.A(new_n546), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n551), .B1(new_n564), .B2(new_n548), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n536), .B(new_n281), .C1(new_n561), .C2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n564), .A2(new_n548), .A3(new_n551), .ZN(new_n567));
  INV_X1    g381(.A(new_n548), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n559), .B2(new_n560), .ZN(new_n569));
  OAI211_X1 g383(.A(G469), .B(new_n567), .C1(new_n569), .C2(new_n551), .ZN(new_n570));
  NAND2_X1  g384(.A1(G469), .A2(G902), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n566), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n336), .B1(new_n442), .B2(new_n281), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n454), .A2(new_n535), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n354), .A2(new_n355), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(G101), .ZN(G3));
  INV_X1    g392(.A(new_n351), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n259), .A2(new_n281), .A3(new_n267), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G472), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n268), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n579), .A2(new_n582), .A3(new_n575), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n517), .B1(new_n491), .B2(new_n509), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n521), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n532), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT96), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n585), .A2(KEYINPUT96), .A3(new_n532), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(G478), .B1(new_n449), .B2(new_n281), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT97), .B1(new_n447), .B2(new_n448), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT33), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g408(.A(KEYINPUT97), .B(KEYINPUT33), .C1(new_n447), .C2(new_n448), .ZN(new_n595));
  AOI21_X1  g409(.A(G902), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n591), .B1(new_n596), .B2(G478), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n410), .B2(new_n415), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n590), .A2(new_n599), .A3(new_n531), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n583), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT34), .B(G104), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G6));
  NAND3_X1  g417(.A1(new_n399), .A2(new_n403), .A3(new_n406), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n604), .A2(new_n415), .ZN(new_n605));
  INV_X1    g419(.A(new_n453), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n590), .A2(new_n607), .A3(new_n531), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n583), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT35), .B(G107), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G9));
  NAND2_X1  g425(.A1(new_n344), .A2(new_n345), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n287), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n614));
  OR2_X1    g428(.A1(new_n339), .A2(KEYINPUT36), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n334), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n334), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n349), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n613), .A2(new_n614), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT98), .B1(new_n346), .B2(new_n619), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n576), .A2(new_n268), .A3(new_n581), .A4(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT37), .B(G110), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT99), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n624), .B(new_n626), .ZN(G12));
  INV_X1    g441(.A(new_n575), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n588), .A2(new_n628), .A3(new_n589), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n527), .B(KEYINPUT101), .Z(new_n630));
  INV_X1    g444(.A(G900), .ZN(new_n631));
  OR2_X1    g445(.A1(new_n631), .A2(KEYINPUT100), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(KEYINPUT100), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n630), .B1(new_n528), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT102), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n605), .A2(new_n606), .A3(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n623), .A2(new_n629), .A3(new_n284), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G128), .ZN(G30));
  AND2_X1   g453(.A1(new_n522), .A2(new_n523), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n522), .A2(new_n523), .ZN(new_n643));
  INV_X1    g457(.A(new_n641), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n636), .B(KEYINPUT39), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n628), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(KEYINPUT40), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n416), .A2(new_n606), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n648), .A2(KEYINPUT40), .ZN(new_n652));
  AND4_X1   g466(.A1(new_n646), .A2(new_n649), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n621), .A2(new_n622), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n273), .A2(new_n265), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n281), .B1(new_n278), .B2(new_n246), .ZN(new_n656));
  OAI21_X1  g470(.A(G472), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n270), .A2(new_n271), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT104), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n270), .A2(new_n660), .A3(new_n271), .A4(new_n657), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n653), .A2(new_n532), .A3(new_n654), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G143), .ZN(G45));
  INV_X1    g478(.A(new_n597), .ZN(new_n665));
  AND4_X1   g479(.A1(KEYINPUT105), .A2(new_n416), .A3(new_n665), .A4(new_n636), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT105), .B1(new_n598), .B2(new_n636), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n668), .A2(new_n284), .A3(new_n623), .A4(new_n629), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT106), .B(G146), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G48));
  INV_X1    g485(.A(new_n352), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n561), .A2(new_n565), .ZN(new_n673));
  OAI21_X1  g487(.A(G469), .B1(new_n673), .B2(G902), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n566), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n573), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n672), .A2(new_n600), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT41), .B(G113), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G15));
  NAND3_X1  g493(.A1(new_n672), .A2(new_n608), .A3(new_n676), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G116), .ZN(G18));
  AND2_X1   g495(.A1(new_n623), .A2(new_n284), .ZN(new_n682));
  INV_X1    g496(.A(new_n454), .ZN(new_n683));
  INV_X1    g497(.A(new_n531), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n676), .A2(new_n588), .A3(new_n589), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n682), .A2(new_n683), .A3(new_n684), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G119), .ZN(G21));
  OAI211_X1 g502(.A(new_n262), .B(new_n250), .C1(new_n246), .C2(new_n279), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n260), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n581), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n579), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n650), .A2(KEYINPUT107), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n416), .A2(new_n606), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n692), .A2(new_n684), .A3(new_n686), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G122), .ZN(G24));
  NAND4_X1  g512(.A1(new_n621), .A2(new_n622), .A3(new_n581), .A4(new_n690), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n668), .A3(new_n686), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G125), .ZN(G27));
  XNOR2_X1  g516(.A(new_n575), .B(KEYINPUT108), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n284), .A3(new_n351), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n416), .A2(new_n665), .A3(new_n636), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n598), .A2(KEYINPUT105), .A3(new_n636), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n533), .B1(new_n522), .B2(new_n523), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n705), .A2(KEYINPUT42), .A3(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n714), .B1(new_n704), .B2(new_n711), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT109), .B(G131), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G33));
  NAND3_X1  g532(.A1(new_n705), .A2(new_n637), .A3(new_n710), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G134), .ZN(G36));
  OAI21_X1  g534(.A(KEYINPUT43), .B1(new_n416), .B2(new_n597), .ZN(new_n721));
  OR3_X1    g535(.A1(new_n416), .A2(KEYINPUT43), .A3(new_n597), .ZN(new_n722));
  AND4_X1   g536(.A1(new_n582), .A2(new_n623), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n724));
  OR3_X1    g538(.A1(new_n723), .A2(new_n724), .A3(KEYINPUT44), .ZN(new_n725));
  INV_X1    g539(.A(new_n710), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n726), .B1(new_n723), .B2(KEYINPUT44), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n724), .B1(new_n723), .B2(KEYINPUT44), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n725), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT112), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n559), .A2(new_n560), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n551), .B1(new_n732), .B2(new_n548), .ZN(new_n733));
  INV_X1    g547(.A(new_n567), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n731), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI211_X1 g549(.A(KEYINPUT45), .B(new_n567), .C1(new_n569), .C2(new_n551), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(G469), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n571), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n566), .B1(new_n738), .B2(new_n740), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n739), .B1(new_n738), .B2(new_n740), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n573), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n746), .A2(new_n647), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT112), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n725), .A2(new_n748), .A3(new_n727), .A4(new_n728), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n730), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G137), .ZN(G39));
  OR2_X1    g565(.A1(new_n742), .A2(new_n744), .ZN(new_n752));
  OAI211_X1 g566(.A(KEYINPUT47), .B(new_n574), .C1(new_n752), .C2(new_n743), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT47), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n754), .B1(new_n745), .B2(new_n573), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n284), .A2(new_n351), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n712), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G140), .ZN(G42));
  NAND4_X1  g573(.A1(new_n417), .A2(new_n574), .A3(new_n532), .A4(new_n665), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n579), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n646), .B1(new_n761), .B2(KEYINPUT113), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n761), .A2(KEYINPUT113), .ZN(new_n763));
  INV_X1    g577(.A(new_n662), .ZN(new_n764));
  XOR2_X1   g578(.A(new_n675), .B(KEYINPUT49), .Z(new_n765));
  NAND4_X1  g579(.A1(new_n762), .A2(new_n763), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n346), .A2(new_n619), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n628), .A2(new_n636), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n590), .B1(new_n693), .B2(new_n695), .ZN(new_n770));
  AND4_X1   g584(.A1(new_n768), .A2(new_n662), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n669), .A2(new_n701), .A3(new_n638), .ZN(new_n772));
  OAI21_X1  g586(.A(KEYINPUT116), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n638), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n708), .A2(new_n709), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n775), .A2(new_n699), .A3(new_n685), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n662), .A2(new_n770), .A3(new_n768), .A4(new_n769), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n777), .A2(new_n778), .A3(new_n669), .A4(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n773), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT52), .B1(new_n771), .B2(new_n772), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n640), .A2(KEYINPUT114), .A3(new_n534), .A4(new_n598), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n416), .A2(new_n453), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n640), .A2(new_n534), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n788), .B1(new_n535), .B2(new_n599), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n785), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n583), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n577), .A2(new_n791), .A3(new_n624), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT115), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n577), .A2(new_n791), .A3(new_n794), .A4(new_n624), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n687), .A2(new_n680), .A3(new_n677), .A4(new_n697), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n581), .A2(new_n690), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n799), .A2(new_n703), .A3(new_n708), .A4(new_n709), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n284), .A2(new_n769), .A3(new_n453), .A4(new_n605), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n623), .A3(new_n710), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n716), .A2(new_n719), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n796), .A2(new_n798), .A3(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n767), .B1(new_n784), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n773), .A2(new_n780), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT52), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n797), .B1(new_n793), .B2(new_n795), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n808), .A2(new_n782), .A3(new_n809), .A4(new_n804), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n806), .B1(new_n767), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT54), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n767), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n796), .A2(new_n798), .A3(new_n804), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(KEYINPUT53), .A3(new_n782), .A4(new_n783), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT117), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n710), .A2(new_n676), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT120), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT120), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n710), .A2(new_n821), .A3(new_n676), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n579), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n527), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n823), .A2(new_n764), .A3(new_n824), .A4(new_n598), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n825), .A2(new_n524), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n722), .A2(new_n630), .A3(new_n721), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n722), .A2(KEYINPUT118), .A3(new_n630), .A4(new_n721), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(new_n686), .A3(new_n692), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n826), .A2(KEYINPUT123), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT123), .B1(new_n826), .B2(new_n832), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n829), .A2(new_n830), .B1(new_n822), .B2(new_n820), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n672), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n837), .B(KEYINPUT48), .Z(new_n838));
  NAND3_X1  g652(.A1(new_n831), .A2(new_n692), .A3(new_n710), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n674), .A2(new_n573), .A3(new_n566), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n753), .A2(new_n755), .A3(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n831), .A2(KEYINPUT119), .A3(new_n692), .A4(new_n710), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n841), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n533), .A2(new_n642), .A3(new_n645), .A4(new_n676), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n831), .A2(new_n846), .A3(new_n692), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT50), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n831), .A2(new_n846), .A3(KEYINPUT50), .A4(new_n692), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n836), .A2(new_n700), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n845), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n416), .A2(new_n665), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n823), .A2(new_n764), .A3(new_n824), .A4(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT121), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n845), .A2(new_n851), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT51), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g675(.A(KEYINPUT51), .B(new_n859), .C1(new_n853), .C2(new_n856), .ZN(new_n862));
  AOI211_X1 g676(.A(new_n835), .B(new_n838), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n813), .A2(new_n816), .A3(new_n864), .A4(new_n814), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n812), .A2(new_n818), .A3(new_n863), .A4(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(G952), .A2(G953), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n766), .B1(new_n866), .B2(new_n867), .ZN(G75));
  AOI21_X1  g682(.A(new_n281), .B1(new_n813), .B2(new_n816), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n517), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n513), .A2(new_n489), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(new_n511), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT55), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n870), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n874), .B1(new_n870), .B2(new_n871), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n358), .A2(G952), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(G51));
  NAND2_X1  g692(.A1(new_n571), .A2(KEYINPUT57), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n571), .A2(KEYINPUT57), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n773), .A2(new_n781), .A3(new_n780), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n781), .B1(new_n773), .B2(new_n780), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT53), .B1(new_n883), .B2(new_n815), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n784), .A2(new_n805), .A3(new_n767), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT54), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n814), .B1(new_n813), .B2(new_n816), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n879), .B(new_n880), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n673), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n737), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n869), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n877), .B1(new_n890), .B2(new_n892), .ZN(G54));
  AND2_X1   g707(.A1(KEYINPUT58), .A2(G475), .ZN(new_n894));
  OAI211_X1 g708(.A(G902), .B(new_n894), .C1(new_n884), .C2(new_n885), .ZN(new_n895));
  INV_X1    g709(.A(new_n404), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n877), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n813), .A2(new_n816), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n899), .A2(G902), .A3(new_n404), .A4(new_n894), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n897), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n897), .A2(KEYINPUT124), .A3(new_n900), .A4(new_n898), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(G60));
  AND2_X1   g719(.A1(new_n594), .A2(new_n595), .ZN(new_n906));
  NAND2_X1  g720(.A1(G478), .A2(G902), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT59), .Z(new_n908));
  NOR2_X1   g722(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(new_n886), .B2(new_n887), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n898), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n818), .A2(new_n812), .A3(new_n865), .ZN(new_n912));
  INV_X1    g726(.A(new_n908), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n911), .B1(new_n914), .B2(new_n906), .ZN(G63));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n916));
  NAND2_X1  g730(.A1(G217), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT60), .Z(new_n918));
  NAND4_X1  g732(.A1(new_n899), .A2(new_n616), .A3(new_n617), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n898), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n348), .B1(new_n899), .B2(new_n918), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n916), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n921), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n923), .A2(KEYINPUT61), .A3(new_n898), .A4(new_n919), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n922), .A2(new_n924), .ZN(G66));
  INV_X1    g739(.A(G224), .ZN(new_n926));
  OAI21_X1  g740(.A(G953), .B1(new_n529), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(new_n809), .B2(G953), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n872), .B1(G898), .B2(new_n358), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(G69));
  AND2_X1   g744(.A1(new_n223), .A2(new_n235), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n370), .A2(new_n373), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n931), .B(new_n932), .Z(new_n933));
  NAND2_X1  g747(.A1(G900), .A2(G953), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n772), .B(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n747), .A2(new_n672), .A3(new_n770), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n758), .A2(new_n937), .A3(new_n719), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n750), .A2(new_n716), .A3(new_n936), .A4(new_n938), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n933), .B(new_n934), .C1(new_n939), .C2(G953), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n358), .B1(G227), .B2(G900), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n936), .A2(new_n663), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n599), .B1(new_n453), .B2(new_n416), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n726), .A2(new_n648), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n354), .A2(new_n355), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT126), .Z(new_n952));
  NAND4_X1  g766(.A1(new_n948), .A2(new_n750), .A3(new_n758), .A4(new_n952), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n953), .A2(new_n358), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n943), .B(new_n945), .C1(new_n954), .C2(new_n933), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n933), .B1(new_n953), .B2(new_n358), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n944), .B1(new_n956), .B2(new_n942), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n957), .ZN(G72));
  NAND2_X1  g772(.A1(G472), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT63), .Z(new_n960));
  INV_X1    g774(.A(new_n809), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n960), .B1(new_n939), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n274), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n655), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n811), .A2(new_n274), .A3(new_n965), .A4(new_n960), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n964), .A2(new_n898), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n960), .B1(new_n953), .B2(new_n961), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n967), .B1(new_n655), .B2(new_n968), .ZN(G57));
endmodule


