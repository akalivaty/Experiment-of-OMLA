//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1315,
    new_n1316, new_n1317, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT64), .Z(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G226), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G68), .B(G77), .Z(new_n236));
  XNOR2_X1  g0036(.A(G50), .B(G58), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  XNOR2_X1  g0042(.A(KEYINPUT3), .B(G33), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G1698), .ZN(new_n244));
  INV_X1    g0044(.A(KEYINPUT67), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G223), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n250), .A2(G222), .B1(G77), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n247), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n215), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(KEYINPUT65), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT65), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(G33), .A3(G41), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n263), .A2(new_n265), .A3(new_n258), .ZN(new_n266));
  INV_X1    g0066(.A(G41), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  AOI21_X1  g0068(.A(G1), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n266), .A2(G274), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n269), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G226), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n270), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OR2_X1    g0074(.A1(new_n274), .A2(KEYINPUT66), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(KEYINPUT66), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n262), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G200), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n215), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT68), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n283), .B(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n201), .B1(new_n206), .B2(G20), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G150), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT8), .B(G58), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n253), .A2(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n288), .B(new_n290), .C1(new_n291), .C2(new_n293), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n294), .A2(new_n282), .B1(new_n201), .B2(new_n280), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n287), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT9), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n278), .B(new_n297), .C1(new_n298), .C2(new_n277), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT10), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n277), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n302), .B(new_n296), .C1(G179), .C2(new_n277), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(G223), .A2(G1698), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(new_n273), .B2(G1698), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT73), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n253), .ZN(new_n308));
  NAND2_X1  g0108(.A1(KEYINPUT73), .A2(G33), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(KEYINPUT3), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n306), .A2(new_n310), .A3(new_n252), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G87), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT75), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n311), .A2(KEYINPUT75), .A3(new_n312), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(new_n316), .A3(new_n261), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n270), .B1(new_n272), .B2(new_n228), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(G179), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n260), .B1(new_n313), .B2(new_n314), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n318), .B1(new_n321), .B2(new_n316), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n320), .B1(new_n301), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G68), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n202), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(G58), .A2(G68), .ZN(new_n326));
  OAI21_X1  g0126(.A(G20), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n289), .A2(G159), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(G20), .B1(new_n310), .B2(new_n252), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT7), .ZN(new_n332));
  OAI21_X1  g0132(.A(G68), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AOI211_X1 g0133(.A(KEYINPUT7), .B(G20), .C1(new_n310), .C2(new_n252), .ZN(new_n334));
  OAI211_X1 g0134(.A(KEYINPUT16), .B(new_n330), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n332), .A2(G20), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT3), .B1(new_n308), .B2(new_n309), .ZN(new_n338));
  INV_X1    g0138(.A(new_n254), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n332), .B1(new_n243), .B2(G20), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n324), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n336), .B1(new_n342), .B2(new_n329), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n335), .A2(new_n343), .A3(new_n282), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n291), .B1(new_n206), .B2(G20), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n285), .A2(new_n345), .B1(new_n280), .B2(new_n291), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT18), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n323), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n348), .B1(new_n323), .B2(new_n347), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT76), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n323), .A2(new_n347), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT18), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT76), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n323), .A2(new_n347), .A3(new_n348), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n311), .A2(KEYINPUT75), .A3(new_n312), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT75), .B1(new_n311), .B2(new_n312), .ZN(new_n358));
  NOR3_X1   g0158(.A1(new_n357), .A2(new_n358), .A3(new_n260), .ZN(new_n359));
  OAI21_X1  g0159(.A(G200), .B1(new_n359), .B2(new_n318), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n317), .A2(G190), .A3(new_n319), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n360), .A2(new_n344), .A3(new_n346), .A4(new_n361), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT17), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n351), .A2(new_n356), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n289), .A2(G50), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT70), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n365), .B(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G77), .ZN(new_n368));
  OAI22_X1  g0168(.A1(new_n293), .A2(new_n368), .B1(new_n207), .B2(G68), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n282), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT11), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g0172(.A(KEYINPUT11), .B(new_n282), .C1(new_n367), .C2(new_n369), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT12), .B1(new_n279), .B2(G68), .ZN(new_n374));
  OR3_X1    g0174(.A1(new_n279), .A2(KEYINPUT12), .A3(G68), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n324), .B1(new_n206), .B2(G20), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n374), .A2(new_n375), .B1(new_n283), .B2(new_n376), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n372), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n266), .A2(G238), .A3(new_n271), .ZN(new_n379));
  NOR2_X1   g0179(.A1(G226), .A2(G1698), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n380), .B1(new_n228), .B2(G1698), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(new_n243), .B1(G33), .B2(G97), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n270), .B(new_n379), .C1(new_n382), .C2(new_n260), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT13), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n228), .A2(G1698), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(G226), .B2(G1698), .ZN(new_n386));
  INV_X1    g0186(.A(G97), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n386), .A2(new_n255), .B1(new_n253), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n261), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT13), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n389), .A2(new_n390), .A3(new_n270), .A4(new_n379), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n384), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n378), .B1(new_n298), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G200), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n394), .B1(new_n384), .B2(new_n391), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n384), .A2(G179), .A3(new_n391), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n301), .B1(new_n384), .B2(new_n391), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT14), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n392), .A2(new_n399), .A3(G169), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT71), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n398), .A2(KEYINPUT71), .A3(new_n399), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n400), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n378), .A2(KEYINPUT72), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n372), .A2(new_n373), .A3(new_n377), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT72), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n396), .B1(new_n405), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n282), .ZN(new_n412));
  XNOR2_X1  g0212(.A(KEYINPUT15), .B(G87), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(new_n292), .B1(G20), .B2(G77), .ZN(new_n415));
  INV_X1    g0215(.A(new_n291), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n289), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n412), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n280), .A2(new_n368), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT69), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n419), .B(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n368), .B1(new_n206), .B2(G20), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n283), .A2(new_n422), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n418), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n266), .A2(G244), .A3(new_n271), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n425), .A2(new_n270), .ZN(new_n426));
  INV_X1    g0226(.A(G107), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n249), .A2(new_n228), .B1(new_n427), .B2(new_n243), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n428), .B1(new_n246), .B2(G238), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n426), .B1(new_n429), .B2(new_n260), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n424), .B1(new_n430), .B2(new_n301), .ZN(new_n431));
  INV_X1    g0231(.A(G179), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n432), .B(new_n426), .C1(new_n429), .C2(new_n260), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n430), .A2(G200), .ZN(new_n435));
  OAI211_X1 g0235(.A(G190), .B(new_n426), .C1(new_n429), .C2(new_n260), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n436), .A3(new_n424), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NOR4_X1   g0238(.A1(new_n304), .A2(new_n364), .A3(new_n411), .A4(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n268), .A2(G1), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n440), .A2(G250), .ZN(new_n441));
  OR3_X1    g0241(.A1(new_n268), .A2(G1), .A3(G274), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(new_n266), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n252), .ZN(new_n444));
  AND2_X1   g0244(.A1(KEYINPUT73), .A2(G33), .ZN(new_n445));
  NOR2_X1   g0245(.A1(KEYINPUT73), .A2(G33), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n444), .B1(new_n447), .B2(KEYINPUT3), .ZN(new_n448));
  NOR2_X1   g0248(.A1(G238), .A2(G1698), .ZN(new_n449));
  INV_X1    g0249(.A(G244), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n449), .B1(new_n450), .B2(G1698), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n308), .A2(new_n309), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n448), .A2(new_n451), .B1(G116), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n443), .B1(new_n453), .B2(new_n260), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n206), .A2(G33), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n279), .A2(new_n455), .A3(new_n215), .A4(new_n281), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT78), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n454), .A2(G200), .B1(G87), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n207), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT82), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT82), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n459), .A2(new_n462), .A3(new_n207), .ZN(new_n463));
  INV_X1    g0263(.A(G87), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(new_n387), .A3(new_n427), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n461), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n310), .A2(new_n207), .A3(G68), .A4(new_n252), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT19), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(new_n293), .B2(new_n387), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n282), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n414), .A2(new_n279), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT83), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT83), .ZN(new_n475));
  AOI211_X1 g0275(.A(new_n475), .B(new_n472), .C1(new_n470), .C2(new_n282), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n458), .B(KEYINPUT85), .C1(new_n474), .C2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n454), .A2(new_n298), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT85), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n474), .A2(new_n476), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n457), .A2(G87), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n451), .A2(new_n310), .A3(new_n252), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n452), .A2(G116), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n260), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n443), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n483), .B1(new_n488), .B2(new_n394), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n481), .B1(new_n482), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n454), .A2(G169), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n488), .A2(G179), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n457), .A2(new_n414), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(new_n474), .B2(new_n476), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n494), .B1(new_n496), .B2(KEYINPUT84), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT84), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n498), .B(new_n495), .C1(new_n474), .C2(new_n476), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n480), .A2(new_n490), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g0300(.A(G97), .B(G107), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT6), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n502), .A2(new_n387), .A3(G107), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n207), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n289), .A2(G77), .ZN(new_n507));
  XNOR2_X1  g0307(.A(new_n507), .B(KEYINPUT77), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n337), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n251), .B1(new_n445), .B2(new_n446), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n510), .B1(new_n511), .B2(new_n254), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT7), .B1(new_n255), .B2(new_n207), .ZN(new_n513));
  OAI21_X1  g0313(.A(G107), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n412), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n279), .A2(new_n387), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT78), .ZN(new_n518));
  XNOR2_X1  g0318(.A(new_n456), .B(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n517), .B1(new_n519), .B2(G97), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g0321(.A(KEYINPUT5), .B(G41), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n440), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(G257), .A3(new_n266), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n266), .A2(G274), .A3(new_n440), .A4(new_n522), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n243), .A2(G250), .A3(G1698), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G283), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT79), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(KEYINPUT79), .A2(G33), .A3(G283), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT4), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(new_n450), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n534), .A2(new_n248), .A3(new_n252), .A4(new_n254), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n527), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n310), .A2(new_n252), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n450), .A2(G1698), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n533), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n526), .B1(new_n541), .B2(new_n261), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G190), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT80), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n527), .A2(new_n532), .A3(new_n535), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n448), .A2(new_n538), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n545), .B1(new_n533), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n544), .B1(new_n547), .B2(new_n260), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n541), .A2(KEYINPUT80), .A3(new_n261), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n526), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n521), .B(new_n543), .C1(new_n550), .C2(new_n394), .ZN(new_n551));
  OAI21_X1  g0351(.A(KEYINPUT81), .B1(new_n515), .B2(new_n520), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n427), .B1(new_n340), .B2(new_n341), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT77), .ZN(new_n554));
  XNOR2_X1  g0354(.A(new_n507), .B(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n504), .B1(new_n502), .B2(new_n501), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n555), .B1(new_n207), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n282), .B1(new_n553), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT81), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n516), .B1(new_n457), .B2(new_n387), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n552), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n526), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n547), .B2(new_n260), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n301), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT80), .B1(new_n541), .B2(new_n261), .ZN(new_n566));
  AOI211_X1 g0366(.A(new_n544), .B(new_n260), .C1(new_n536), .C2(new_n540), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n432), .B(new_n563), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n562), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n243), .A2(new_n207), .A3(G87), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT22), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT23), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n207), .B2(G107), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n427), .A2(KEYINPUT23), .A3(G20), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n570), .A2(new_n571), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT24), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n207), .A2(G87), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(new_n571), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n310), .A2(new_n578), .A3(new_n252), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n452), .A2(new_n207), .A3(G116), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n575), .A2(new_n576), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n571), .B1(new_n255), .B2(new_n577), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n573), .A2(new_n574), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n579), .A2(new_n582), .A3(new_n583), .A4(new_n580), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT24), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n412), .B1(new_n581), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n279), .A2(G107), .ZN(new_n587));
  XNOR2_X1  g0387(.A(new_n587), .B(KEYINPUT25), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n519), .B2(new_n427), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n523), .A2(G264), .A3(new_n266), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n525), .ZN(new_n592));
  NOR2_X1   g0392(.A1(G250), .A2(G1698), .ZN(new_n593));
  INV_X1    g0393(.A(G257), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n593), .B1(new_n594), .B2(G1698), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(new_n310), .A3(new_n252), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n452), .A2(G294), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n260), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n592), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G190), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n590), .B(new_n600), .C1(new_n394), .C2(new_n599), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n551), .A2(new_n569), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n523), .A2(G270), .A3(new_n266), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n525), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G264), .A2(G1698), .ZN(new_n606));
  INV_X1    g0406(.A(G303), .ZN(new_n607));
  OAI22_X1  g0407(.A1(new_n537), .A2(new_n606), .B1(new_n607), .B2(new_n243), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT86), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n594), .A2(G1698), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n448), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n310), .A2(new_n252), .A3(new_n610), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT86), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n608), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(G190), .B(new_n605), .C1(new_n614), .C2(new_n260), .ZN(new_n615));
  INV_X1    g0415(.A(G116), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n281), .A2(new_n215), .B1(G20), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n532), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n207), .B1(new_n387), .B2(G33), .ZN(new_n619));
  OAI211_X1 g0419(.A(KEYINPUT20), .B(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT20), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n619), .B1(new_n530), .B2(new_n531), .ZN(new_n622));
  INV_X1    g0422(.A(new_n617), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  MUX2_X1   g0425(.A(new_n279), .B(new_n456), .S(G116), .Z(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n611), .A2(new_n613), .ZN(new_n629));
  INV_X1    g0429(.A(new_n608), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n604), .B1(new_n631), .B2(new_n261), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n615), .B(new_n628), .C1(new_n632), .C2(new_n394), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(G179), .A3(new_n627), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n301), .B1(new_n625), .B2(new_n626), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT21), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n260), .B1(new_n629), .B2(new_n630), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n604), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n605), .B1(new_n614), .B2(new_n260), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n636), .B1(new_n640), .B2(new_n635), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n633), .B(new_n634), .C1(new_n639), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n596), .A2(new_n597), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n261), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n644), .A2(G179), .A3(new_n525), .A4(new_n591), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n301), .B2(new_n599), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n586), .B2(new_n589), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n642), .A2(new_n648), .ZN(new_n649));
  AND4_X1   g0449(.A1(new_n439), .A2(new_n500), .A3(new_n602), .A4(new_n649), .ZN(G372));
  OAI21_X1  g0450(.A(new_n483), .B1(new_n474), .B2(new_n476), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT87), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT87), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n653), .B(new_n483), .C1(new_n474), .C2(new_n476), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n478), .B1(G200), .B2(new_n454), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n652), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n496), .A2(new_n493), .ZN(new_n657));
  INV_X1    g0457(.A(new_n521), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n568), .A2(new_n565), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n656), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n490), .A2(new_n479), .A3(new_n477), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n496), .A2(KEYINPUT84), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n664), .A2(new_n499), .A3(new_n493), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n562), .A2(new_n565), .A3(new_n568), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n663), .A2(new_n665), .A3(new_n666), .A4(KEYINPUT26), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n657), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n647), .B(new_n634), .C1(new_n639), .C2(new_n641), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n670), .A2(new_n656), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n669), .B1(new_n671), .B2(new_n602), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n439), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n349), .A2(new_n350), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n405), .A2(new_n410), .ZN(new_n676));
  INV_X1    g0476(.A(new_n434), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n676), .B1(new_n396), .B2(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n344), .A2(new_n346), .ZN(new_n679));
  AOI211_X1 g0479(.A(new_n298), .B(new_n318), .C1(new_n321), .C2(new_n316), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n394), .B1(new_n317), .B2(new_n319), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n679), .A2(new_n682), .A3(KEYINPUT17), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT17), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n361), .B1(new_n394), .B2(new_n322), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n684), .B1(new_n685), .B2(new_n347), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n675), .B1(new_n678), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n300), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n689), .A2(new_n303), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n674), .A2(new_n690), .ZN(G369));
  XNOR2_X1  g0491(.A(KEYINPUT90), .B(G330), .ZN(new_n692));
  INV_X1    g0492(.A(new_n642), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(KEYINPUT88), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(KEYINPUT88), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT27), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT27), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n695), .A2(new_n696), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n698), .A2(new_n700), .A3(G213), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT89), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n698), .A2(new_n700), .A3(KEYINPUT89), .A4(G213), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n703), .A2(G343), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n693), .B1(new_n628), .B2(new_n706), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n639), .A2(new_n641), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n634), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n709), .A2(new_n627), .A3(new_n705), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n692), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n601), .A2(new_n647), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n586), .A2(new_n589), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n705), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT91), .B1(new_n647), .B2(new_n706), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT91), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n714), .A2(new_n717), .A3(new_n646), .A4(new_n705), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n713), .A2(new_n715), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n712), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n713), .A2(new_n715), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n716), .A2(new_n718), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n705), .B1(new_n708), .B2(new_n634), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n724), .A2(new_n725), .B1(new_n648), .B2(new_n706), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n721), .A2(new_n726), .ZN(G399));
  NAND2_X1  g0527(.A1(new_n210), .A2(new_n267), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n465), .A2(G116), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(G1), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n213), .B2(new_n728), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT92), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT28), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT93), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n599), .A2(G179), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n640), .A2(new_n454), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n550), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n564), .A2(new_n637), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n488), .A2(new_n603), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n645), .ZN(new_n740));
  AOI21_X1  g0540(.A(KEYINPUT30), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n734), .B1(new_n737), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n738), .A2(KEYINPUT30), .A3(new_n740), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT30), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n631), .A2(new_n261), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n542), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n599), .A2(new_n488), .A3(G179), .A4(new_n603), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n744), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n748), .B(KEYINPUT93), .C1(new_n550), .C2(new_n736), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n742), .A2(new_n743), .A3(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT31), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n706), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n748), .B(new_n743), .C1(new_n550), .C2(new_n736), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n705), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n750), .A2(new_n752), .B1(new_n754), .B2(new_n751), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n500), .A2(new_n649), .A3(new_n602), .A4(new_n706), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n692), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n673), .A2(new_n706), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT29), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n661), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n656), .A2(KEYINPUT26), .A3(new_n659), .A4(new_n657), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n705), .B1(new_n764), .B2(new_n672), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(KEYINPUT29), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n757), .B1(new_n760), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n733), .B1(new_n767), .B2(G1), .ZN(G364));
  NAND3_X1  g0568(.A1(new_n707), .A2(new_n710), .A3(new_n692), .ZN(new_n769));
  INV_X1    g0569(.A(new_n728), .ZN(new_n770));
  INV_X1    g0570(.A(G13), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n206), .B1(new_n772), .B2(G45), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n712), .B(new_n769), .C1(new_n770), .C2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G13), .A2(G33), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n707), .A2(new_n710), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n770), .A2(new_n774), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n207), .A2(new_n298), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n394), .A2(G179), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G190), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n243), .B1(new_n783), .B2(new_n464), .C1(new_n324), .C2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n432), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n781), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n207), .A2(G190), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(G58), .A2(new_n790), .B1(new_n793), .B2(G77), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n791), .A2(new_n782), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n794), .B1(new_n427), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n784), .A2(new_n298), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n787), .B(new_n796), .C1(G50), .C2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(G179), .A2(G200), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT95), .ZN(new_n800));
  INV_X1    g0600(.A(new_n791), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g0602(.A(KEYINPUT96), .B(G159), .Z(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT32), .Z(new_n806));
  OAI21_X1  g0606(.A(G20), .B1(new_n800), .B2(new_n298), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G97), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n798), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n783), .ZN(new_n810));
  AOI22_X1  g0610(.A1(G303), .A2(new_n810), .B1(new_n790), .B2(G322), .ZN(new_n811));
  INV_X1    g0611(.A(G283), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n812), .B2(new_n795), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(G329), .B2(new_n802), .ZN(new_n814));
  NOR2_X1   g0614(.A1(KEYINPUT33), .A2(G317), .ZN(new_n815));
  AND2_X1   g0615(.A1(KEYINPUT33), .A2(G317), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n785), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G311), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n817), .B(new_n255), .C1(new_n818), .C2(new_n792), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(G326), .B2(new_n797), .ZN(new_n820));
  INV_X1    g0620(.A(G294), .ZN(new_n821));
  INV_X1    g0621(.A(new_n807), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n814), .B(new_n820), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n809), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n215), .B1(G20), .B2(new_n301), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n778), .A2(new_n825), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n210), .A2(new_n537), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n238), .A2(new_n268), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n828), .B(new_n829), .C1(new_n268), .C2(new_n214), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n210), .A2(new_n243), .ZN(new_n831));
  INV_X1    g0631(.A(G355), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n831), .A2(new_n832), .B1(G116), .B2(new_n210), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT94), .Z(new_n834));
  OAI21_X1  g0634(.A(new_n827), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n779), .A2(new_n780), .A3(new_n826), .A4(new_n835), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n775), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(G396));
  NAND3_X1  g0638(.A1(new_n431), .A2(new_n706), .A3(new_n433), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n436), .A2(new_n424), .ZN(new_n840));
  INV_X1    g0640(.A(new_n424), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n840), .A2(new_n435), .B1(new_n841), .B2(new_n705), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n839), .B1(new_n842), .B2(new_n677), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(KEYINPUT99), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n705), .A2(new_n841), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n437), .A2(new_n845), .B1(new_n433), .B2(new_n431), .ZN(new_n846));
  INV_X1    g0646(.A(new_n839), .ZN(new_n847));
  OR3_X1    g0647(.A1(new_n846), .A2(new_n847), .A3(KEYINPUT99), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n758), .A2(new_n844), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n846), .A2(new_n847), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n673), .A2(new_n706), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n755), .A2(new_n756), .ZN(new_n853));
  INV_X1    g0653(.A(new_n692), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n780), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n855), .B2(new_n852), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n825), .A2(new_n776), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT97), .Z(new_n859));
  OAI21_X1  g0659(.A(new_n780), .B1(new_n859), .B2(G77), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n255), .B1(new_n783), .B2(new_n427), .C1(new_n812), .C2(new_n786), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(G303), .B2(new_n797), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n802), .A2(G311), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n795), .A2(new_n464), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n789), .A2(new_n821), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n864), .B(new_n865), .C1(G116), .C2(new_n793), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n862), .A2(new_n808), .A3(new_n863), .A4(new_n866), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n793), .A2(new_n804), .B1(new_n790), .B2(G143), .ZN(new_n868));
  INV_X1    g0668(.A(new_n797), .ZN(new_n869));
  INV_X1    g0669(.A(G137), .ZN(new_n870));
  INV_X1    g0670(.A(G150), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n868), .B1(new_n869), .B2(new_n870), .C1(new_n871), .C2(new_n786), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT34), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n873), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n783), .A2(new_n201), .B1(new_n795), .B2(new_n324), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n807), .B2(G58), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n537), .B1(new_n802), .B2(G132), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT98), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n867), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n860), .B1(new_n881), .B2(new_n825), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n850), .B2(new_n777), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n857), .A2(KEYINPUT100), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT100), .B1(new_n857), .B2(new_n883), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(G384));
  NOR2_X1   g0687(.A1(new_n772), .A2(new_n206), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n406), .A2(new_n409), .A3(new_n705), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n396), .B(new_n889), .C1(new_n405), .C2(new_n410), .ZN(new_n890));
  INV_X1    g0690(.A(new_n410), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n384), .A2(G179), .A3(new_n391), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n392), .A2(G169), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n892), .B1(new_n893), .B2(KEYINPUT14), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n398), .A2(KEYINPUT71), .A3(new_n399), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT71), .B1(new_n398), .B2(new_n399), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n393), .A2(new_n395), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n891), .B(new_n705), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n843), .B1(new_n890), .B2(new_n899), .ZN(new_n900));
  AND4_X1   g0700(.A1(new_n500), .A2(new_n649), .A3(new_n602), .A4(new_n706), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n754), .A2(new_n751), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n753), .A2(KEYINPUT31), .A3(new_n705), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n900), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT40), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n335), .A2(new_n282), .ZN(new_n908));
  INV_X1    g0708(.A(new_n336), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT7), .B1(new_n448), .B2(G20), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n331), .A2(new_n332), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(G68), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n909), .B1(new_n912), .B2(new_n330), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n346), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n703), .A2(new_n704), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n364), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n347), .A2(new_n915), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n352), .A2(new_n919), .A3(new_n362), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n920), .A2(KEYINPUT37), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n323), .A2(new_n914), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(new_n916), .A3(new_n362), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT37), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n918), .A2(KEYINPUT38), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT38), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n920), .B(KEYINPUT37), .Z(new_n928));
  AOI21_X1  g0728(.A(new_n919), .B1(new_n363), .B2(new_n675), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n907), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT103), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n353), .A2(new_n355), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n687), .B1(new_n935), .B2(KEYINPUT76), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n916), .B1(new_n936), .B2(new_n356), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n921), .A2(new_n924), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n927), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n905), .B1(new_n939), .B2(new_n926), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n934), .B1(new_n940), .B2(KEYINPUT40), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n899), .A2(new_n890), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n850), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n902), .A2(new_n903), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n943), .B1(new_n944), .B2(new_n756), .ZN(new_n945));
  AOI221_X4 g0745(.A(new_n927), .B1(new_n921), .B2(new_n924), .C1(new_n364), .C2(new_n917), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT38), .B1(new_n918), .B2(new_n925), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(KEYINPUT103), .A3(new_n906), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n933), .B1(new_n941), .B2(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT104), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n756), .A2(new_n902), .A3(new_n903), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n439), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n692), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n954), .B2(new_n951), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n851), .A2(new_n839), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n942), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n946), .A2(new_n947), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n958), .A2(new_n959), .B1(new_n675), .B2(new_n915), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT101), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n675), .A2(new_n915), .ZN(new_n962));
  INV_X1    g0762(.A(new_n942), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n851), .B2(new_n839), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n939), .A2(new_n926), .ZN(new_n965));
  AOI211_X1 g0765(.A(KEYINPUT101), .B(new_n962), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n676), .A2(new_n706), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT102), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT39), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n931), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n939), .A2(KEYINPUT39), .A3(new_n926), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n961), .B(new_n967), .C1(new_n969), .C2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n439), .A2(new_n760), .A3(new_n766), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n690), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n974), .B(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n888), .B1(new_n956), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n977), .B2(new_n956), .ZN(new_n979));
  INV_X1    g0779(.A(new_n556), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n980), .A2(KEYINPUT35), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(KEYINPUT35), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n981), .A2(G116), .A3(new_n216), .A4(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT36), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n325), .A2(new_n213), .A3(new_n368), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n324), .A2(G50), .ZN(new_n986));
  OAI211_X1 g0786(.A(G1), .B(new_n771), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n979), .A2(new_n984), .A3(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT105), .ZN(G367));
  OAI221_X1 g0789(.A(new_n827), .B1(new_n210), .B2(new_n413), .C1(new_n234), .C2(new_n828), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n780), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n255), .B1(new_n790), .B2(G150), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n786), .B2(new_n803), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G58), .A2(new_n810), .B1(new_n793), .B2(G50), .ZN(new_n994));
  INV_X1    g0794(.A(new_n802), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n994), .B1(new_n368), .B2(new_n795), .C1(new_n995), .C2(new_n870), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n993), .B(new_n996), .C1(G143), .C2(new_n797), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n324), .B2(new_n822), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n537), .B1(new_n786), .B2(new_n821), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n789), .A2(new_n607), .B1(new_n792), .B2(new_n812), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n795), .A2(new_n387), .ZN(new_n1001));
  NOR3_X1   g0801(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(G317), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1002), .B1(new_n1003), .B2(new_n995), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n783), .A2(new_n616), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n1005), .A2(KEYINPUT46), .B1(G311), .B2(new_n797), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(KEYINPUT46), .B2(new_n1005), .C1(new_n822), .C2(new_n427), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n998), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT47), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n991), .B1(new_n1009), .B2(new_n825), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n706), .B1(new_n652), .B2(new_n654), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n669), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n656), .A2(new_n657), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1012), .B1(new_n1013), .B2(new_n1011), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n778), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1010), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT109), .Z(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n724), .A2(new_n725), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n709), .A2(new_n706), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n719), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(new_n711), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n767), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n658), .A2(new_n705), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n551), .A2(new_n569), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(KEYINPUT106), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1026), .A2(KEYINPUT106), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n568), .A2(new_n565), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n1028), .A2(new_n1029), .B1(new_n1030), .B2(new_n1025), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n726), .A2(KEYINPUT45), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT45), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1030), .A2(new_n1025), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1026), .A2(KEYINPUT106), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1034), .B1(new_n1035), .B2(new_n1027), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n648), .A2(new_n706), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n719), .B2(new_n1020), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1033), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1032), .A2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g0840(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n1041));
  NAND3_X1  g0841(.A1(new_n1036), .A2(new_n1038), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1041), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n726), .B2(new_n1031), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1040), .A2(new_n721), .A3(new_n1042), .A4(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1032), .A2(new_n1039), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1044), .A2(new_n1042), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n720), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1024), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT108), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1049), .B(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n767), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n728), .B(KEYINPUT41), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n774), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1036), .A2(new_n1019), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT42), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n569), .B1(new_n1036), .B2(new_n647), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n706), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n1057), .A2(new_n1059), .B1(KEYINPUT43), .B2(new_n1014), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1014), .A2(KEYINPUT43), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1060), .B(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n721), .A2(new_n1036), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1062), .B(new_n1063), .Z(new_n1064));
  OAI21_X1  g0864(.A(new_n1018), .B1(new_n1055), .B2(new_n1064), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT110), .Z(G387));
  OAI21_X1  g0866(.A(KEYINPUT113), .B1(new_n1024), .B2(new_n728), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n767), .A2(new_n1023), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n767), .A2(new_n1023), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT113), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1069), .A2(new_n1070), .A3(new_n770), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1067), .A2(new_n1068), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n719), .A2(new_n778), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n831), .A2(new_n729), .B1(G107), .B2(new_n210), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n231), .A2(new_n268), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n729), .ZN(new_n1076));
  AOI211_X1 g0876(.A(G45), .B(new_n1076), .C1(G68), .C2(G77), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n291), .A2(G50), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT50), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n828), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1074), .B1(new_n1075), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n827), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n780), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n783), .A2(new_n368), .B1(new_n792), .B2(new_n324), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1001), .B(new_n1084), .C1(G50), .C2(new_n790), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n807), .A2(new_n414), .ZN(new_n1086));
  INV_X1    g0886(.A(G159), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n448), .B1(new_n869), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n416), .B2(new_n785), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(KEYINPUT111), .B(G150), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n802), .A2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1085), .A2(new_n1086), .A3(new_n1089), .A4(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G317), .A2(new_n790), .B1(new_n793), .B2(G303), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT112), .B(G322), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1093), .B1(new_n869), .B2(new_n1094), .C1(new_n818), .C2(new_n786), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT48), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n807), .A2(G283), .B1(G294), .B2(new_n810), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT49), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n537), .B1(new_n616), .B2(new_n795), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(G326), .B2(new_n802), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1092), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1083), .B1(new_n1106), .B2(new_n825), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1023), .A2(new_n774), .B1(new_n1073), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1072), .A2(new_n1108), .ZN(G393));
  NAND3_X1  g0909(.A1(new_n1048), .A2(KEYINPUT114), .A3(new_n1045), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT114), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1111), .B(new_n720), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1110), .A2(new_n1069), .A3(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1051), .A2(new_n770), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT115), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1110), .A2(new_n1115), .A3(new_n1112), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1115), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1117));
  NOR3_X1   g0917(.A1(new_n1116), .A2(new_n1117), .A3(new_n773), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n827), .B1(new_n387), .B2(new_n210), .C1(new_n241), .C2(new_n828), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n780), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n255), .B1(new_n795), .B2(new_n427), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n783), .A2(new_n812), .B1(new_n792), .B2(new_n821), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n1121), .B(new_n1122), .C1(G303), .C2(new_n785), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n995), .A2(new_n1094), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n869), .A2(new_n1003), .B1(new_n789), .B2(new_n818), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT52), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n807), .A2(G116), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1123), .A2(new_n1124), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n802), .A2(G143), .B1(G68), .B2(new_n810), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT116), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n869), .A2(new_n871), .B1(new_n789), .B2(new_n1087), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT51), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n807), .A2(G77), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n785), .A2(G50), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n537), .B(new_n864), .C1(new_n416), .C2(new_n793), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1128), .B1(new_n1130), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1120), .B1(new_n1137), .B2(new_n825), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n1031), .B2(new_n1015), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NOR3_X1   g0940(.A1(new_n1118), .A2(KEYINPUT117), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT117), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1117), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1110), .A2(new_n1115), .A3(new_n1112), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1143), .A2(new_n774), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1142), .B1(new_n1145), .B2(new_n1139), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1114), .B1(new_n1141), .B2(new_n1146), .ZN(G390));
  XNOR2_X1  g0947(.A(KEYINPUT54), .B(G143), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n790), .A2(G132), .B1(new_n793), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n795), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n255), .B1(new_n1151), .B2(G50), .ZN(new_n1152));
  INV_X1    g0952(.A(G125), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1150), .B(new_n1152), .C1(new_n995), .C2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n810), .A2(new_n1090), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1155), .A2(KEYINPUT53), .B1(new_n797), .B2(G128), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1156), .B1(KEYINPUT53), .B2(new_n1155), .C1(new_n870), .C2(new_n786), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1154), .B(new_n1157), .C1(G159), .C2(new_n807), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n243), .B1(new_n810), .B2(G87), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1159), .B1(new_n869), .B2(new_n812), .C1(new_n427), .C2(new_n786), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G68), .A2(new_n1151), .B1(new_n793), .B2(G97), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1161), .B1(new_n616), .B2(new_n789), .C1(new_n995), .C2(new_n821), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1160), .B(new_n1162), .C1(G77), .C2(new_n807), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n825), .B1(new_n1158), .B2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1164), .B(new_n780), .C1(new_n416), .C2(new_n859), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n973), .B2(new_n776), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT118), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n958), .A2(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n757), .A2(new_n850), .A3(new_n942), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n764), .A2(new_n672), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n846), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(new_n706), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n963), .B1(new_n1172), .B2(new_n839), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n931), .A2(new_n969), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1169), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1167), .B1(new_n1168), .B2(new_n1175), .ZN(new_n1176));
  NOR3_X1   g0976(.A1(new_n946), .A2(new_n947), .A3(new_n970), .ZN(new_n1177));
  AOI21_X1  g0977(.A(KEYINPUT39), .B1(new_n926), .B2(new_n930), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n969), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n1177), .A2(new_n1178), .B1(new_n964), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1169), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n705), .B(new_n846), .C1(new_n764), .C2(new_n672), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n942), .B1(new_n1182), .B2(new_n847), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1179), .B1(new_n926), .B2(new_n930), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1181), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1180), .A2(new_n1185), .A3(KEYINPUT118), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1180), .A2(new_n1187), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n952), .A2(G330), .A3(new_n900), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1176), .A2(new_n1186), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1166), .B1(new_n1190), .B2(new_n774), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n942), .B1(new_n757), .B2(new_n850), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n957), .B1(new_n1192), .B2(new_n1189), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n848), .A2(new_n844), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n952), .A2(G330), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n963), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n847), .B1(new_n765), .B2(new_n1171), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(new_n1197), .A3(new_n1169), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1193), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n439), .A2(G330), .A3(new_n952), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n975), .A2(new_n1200), .A3(new_n690), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n770), .B1(new_n1190), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1168), .A2(new_n1175), .A3(new_n1167), .ZN(new_n1205));
  AOI21_X1  g1005(.A(KEYINPUT118), .B1(new_n1180), .B2(new_n1185), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1204), .B(new_n1202), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(KEYINPUT119), .B(new_n1191), .C1(new_n1203), .C2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1202), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1213), .A2(new_n770), .A3(new_n1207), .ZN(new_n1214));
  AOI21_X1  g1014(.A(KEYINPUT119), .B1(new_n1214), .B2(new_n1191), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1210), .A2(new_n1215), .ZN(G378));
  NOR3_X1   g1016(.A1(new_n940), .A2(new_n934), .A3(KEYINPUT40), .ZN(new_n1217));
  AOI21_X1  g1017(.A(KEYINPUT103), .B1(new_n948), .B2(new_n906), .ZN(new_n1218));
  OAI211_X1 g1018(.A(G330), .B(new_n932), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n304), .B(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n915), .A2(new_n296), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT122), .Z(new_n1223));
  XOR2_X1   g1023(.A(new_n1221), .B(new_n1223), .Z(new_n1224));
  NOR2_X1   g1024(.A1(new_n1219), .A2(new_n1224), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1221), .B(new_n1223), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n950), .B2(G330), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n974), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1219), .A2(new_n1224), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT101), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n1230), .A2(new_n1231), .B1(new_n973), .B2(new_n969), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(new_n966), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n950), .A2(G330), .A3(new_n1226), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1229), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1201), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1228), .A2(new_n1235), .B1(new_n1236), .B2(new_n1207), .ZN(new_n1237));
  OAI21_X1  g1037(.A(KEYINPUT123), .B1(new_n1237), .B2(KEYINPUT57), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n728), .B1(new_n1237), .B2(KEYINPUT57), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1207), .A2(new_n1236), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1229), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1233), .B1(new_n1234), .B2(new_n1229), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1240), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT123), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT57), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1238), .A2(new_n1239), .A3(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n774), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n780), .B1(new_n859), .B2(G50), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n795), .A2(new_n202), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(G107), .B2(new_n790), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n810), .A2(G77), .B1(new_n793), .B2(new_n414), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n785), .A2(G97), .B1(new_n797), .B2(G116), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  AOI211_X1 g1054(.A(G41), .B(new_n448), .C1(new_n802), .C2(G283), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1254), .B(new_n1256), .C1(G68), .C2(new_n807), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1257), .A2(KEYINPUT58), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(G33), .A2(G41), .ZN(new_n1259));
  AOI211_X1 g1059(.A(G50), .B(new_n1259), .C1(new_n537), .C2(new_n267), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1261), .B(KEYINPUT120), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n869), .A2(new_n1153), .ZN(new_n1263));
  INV_X1    g1063(.A(G128), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n789), .A2(new_n1264), .B1(new_n792), .B2(new_n870), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1263), .B(new_n1265), .C1(G132), .C2(new_n785), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n783), .A2(new_n1148), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(KEYINPUT121), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1266), .B(new_n1268), .C1(new_n871), .C2(new_n822), .ZN(new_n1269));
  OR2_X1    g1069(.A1(new_n1269), .A2(KEYINPUT59), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n802), .A2(G124), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1271), .B(new_n1259), .C1(new_n795), .C2(new_n803), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n1269), .B2(KEYINPUT59), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1270), .A2(new_n1273), .B1(new_n1257), .B2(KEYINPUT58), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1262), .A2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1249), .B1(new_n1275), .B2(new_n825), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n1226), .B2(new_n777), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1248), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1247), .A2(new_n1279), .ZN(G375));
  INV_X1    g1080(.A(KEYINPUT124), .ZN(new_n1281));
  OR3_X1    g1081(.A1(new_n1199), .A2(new_n1281), .A3(new_n773), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n780), .B1(new_n859), .B2(G68), .ZN(new_n1283));
  OAI22_X1  g1083(.A1(new_n783), .A2(new_n1087), .B1(new_n792), .B2(new_n871), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n1250), .B(new_n1284), .C1(G137), .C2(new_n790), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n807), .A2(G50), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n786), .A2(new_n1148), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n537), .B(new_n1287), .C1(G132), .C2(new_n797), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n802), .A2(G128), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1285), .A2(new_n1286), .A3(new_n1288), .A4(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1086), .B1(new_n812), .B2(new_n789), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(KEYINPUT125), .ZN(new_n1292));
  OAI22_X1  g1092(.A1(new_n786), .A2(new_n616), .B1(new_n869), .B2(new_n821), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n255), .B1(new_n795), .B2(new_n368), .ZN(new_n1294));
  OAI22_X1  g1094(.A1(new_n783), .A2(new_n387), .B1(new_n792), .B2(new_n427), .ZN(new_n1295));
  NOR3_X1   g1095(.A1(new_n1293), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n607), .B2(new_n995), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1290), .B1(new_n1292), .B2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1283), .B1(new_n1298), .B2(new_n825), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(new_n942), .B2(new_n777), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1281), .B1(new_n1199), .B2(new_n773), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1282), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1212), .A2(new_n1054), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1305), .ZN(G381));
  NAND2_X1  g1106(.A1(new_n1214), .A2(new_n1191), .ZN(new_n1307));
  OAI21_X1  g1107(.A(KEYINPUT117), .B1(new_n1118), .B2(new_n1140), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1145), .A2(new_n1142), .A3(new_n1139), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(G381), .A2(G384), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1072), .A2(new_n837), .A3(new_n1108), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1310), .A2(new_n1311), .A3(new_n1114), .A4(new_n1312), .ZN(new_n1313));
  OR4_X1    g1113(.A1(G387), .A2(new_n1307), .A3(new_n1313), .A4(G375), .ZN(G407));
  INV_X1    g1114(.A(G343), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(G213), .ZN(new_n1316));
  OR3_X1    g1116(.A1(G375), .A2(new_n1307), .A3(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(G407), .A2(G213), .A3(new_n1317), .ZN(G409));
  INV_X1    g1118(.A(new_n1065), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n837), .B1(new_n1072), .B2(new_n1108), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1312), .A2(new_n1320), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1321), .A2(KEYINPUT110), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(G390), .A2(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1321), .B1(new_n1310), .B2(new_n1114), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1319), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1321), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(G390), .A2(new_n1326), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1310), .B(new_n1114), .C1(KEYINPUT110), .C2(new_n1321), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1327), .A2(new_n1328), .A3(new_n1065), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1325), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT61), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1247), .A2(G378), .A3(new_n1279), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1243), .A2(new_n1053), .ZN(new_n1333));
  OAI211_X1 g1133(.A(new_n1214), .B(new_n1191), .C1(new_n1333), .C2(new_n1278), .ZN(new_n1334));
  AOI22_X1  g1134(.A1(new_n1332), .A2(new_n1334), .B1(G213), .B2(new_n1315), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1315), .A2(G213), .A3(G2897), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(new_n1304), .B(KEYINPUT60), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1202), .A2(new_n728), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(G384), .A2(new_n1339), .A3(new_n1303), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(G384), .B1(new_n1339), .B2(new_n1303), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1336), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1339), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n886), .B1(new_n1344), .B2(new_n1302), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1336), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1345), .A2(new_n1340), .A3(new_n1346), .ZN(new_n1347));
  AND2_X1   g1147(.A1(new_n1343), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1332), .A2(new_n1334), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1349), .A2(new_n1316), .A3(new_n1350), .ZN(new_n1351));
  OAI221_X1 g1151(.A(new_n1331), .B1(new_n1335), .B2(new_n1348), .C1(new_n1351), .C2(KEYINPUT62), .ZN(new_n1352));
  AND2_X1   g1152(.A1(new_n1351), .A2(KEYINPUT62), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1330), .B1(new_n1352), .B2(new_n1353), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1325), .A2(new_n1331), .A3(new_n1329), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1349), .A2(new_n1316), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT126), .ZN(new_n1357));
  AND3_X1   g1157(.A1(new_n1343), .A2(new_n1347), .A3(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1357), .B1(new_n1343), .B2(new_n1347), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1358), .A2(new_n1359), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1355), .B1(new_n1356), .B2(new_n1360), .ZN(new_n1361));
  INV_X1    g1161(.A(KEYINPUT63), .ZN(new_n1362));
  AND3_X1   g1162(.A1(new_n1335), .A2(new_n1362), .A3(new_n1350), .ZN(new_n1363));
  AOI21_X1  g1163(.A(new_n1362), .B1(new_n1335), .B2(new_n1350), .ZN(new_n1364));
  OAI211_X1 g1164(.A(new_n1361), .B(KEYINPUT127), .C1(new_n1363), .C2(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1351), .A2(KEYINPUT63), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1335), .A2(new_n1362), .A3(new_n1350), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1367), .A2(new_n1368), .ZN(new_n1369));
  AOI21_X1  g1169(.A(KEYINPUT127), .B1(new_n1369), .B2(new_n1361), .ZN(new_n1370));
  OAI21_X1  g1170(.A(new_n1354), .B1(new_n1366), .B2(new_n1370), .ZN(G405));
  INV_X1    g1171(.A(G375), .ZN(new_n1372));
  OAI21_X1  g1172(.A(new_n1332), .B1(new_n1372), .B2(new_n1307), .ZN(new_n1373));
  AND2_X1   g1173(.A1(new_n1373), .A2(new_n1350), .ZN(new_n1374));
  NOR2_X1   g1174(.A1(new_n1373), .A2(new_n1350), .ZN(new_n1375));
  NOR2_X1   g1175(.A1(new_n1374), .A2(new_n1375), .ZN(new_n1376));
  INV_X1    g1176(.A(new_n1330), .ZN(new_n1377));
  XNOR2_X1  g1177(.A(new_n1376), .B(new_n1377), .ZN(G402));
endmodule


