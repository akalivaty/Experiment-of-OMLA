//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n572, new_n573,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n635, new_n636, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1225, new_n1226;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(G217));
  NAND4_X1  g028(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NAND4_X1  g031(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT67), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n458), .A2(G567), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n463), .B1(new_n456), .B2(G2106), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(new_n462), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XOR2_X1   g041(.A(new_n466), .B(KEYINPUT69), .Z(G319));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n471), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(new_n472), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2104), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n479), .A2(new_n481), .A3(G125), .ZN(new_n482));
  NAND2_X1  g057(.A1(G113), .A2(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n475), .B1(new_n478), .B2(new_n485), .ZN(G160));
  NAND2_X1  g061(.A1(new_n479), .A2(new_n481), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(new_n472), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT71), .ZN(new_n490));
  INV_X1    g065(.A(G136), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n473), .B2(new_n491), .ZN(new_n492));
  OR2_X1    g067(.A1(G100), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n487), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(KEYINPUT71), .A3(G136), .ZN(new_n496));
  AND4_X1   g071(.A1(new_n489), .A2(new_n492), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  XOR2_X1   g072(.A(new_n497), .B(KEYINPUT72), .Z(G162));
  NAND4_X1  g073(.A1(new_n479), .A2(new_n481), .A3(G138), .A4(new_n472), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n472), .A2(KEYINPUT4), .A3(G138), .ZN(new_n502));
  INV_X1    g077(.A(G126), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(new_n472), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(new_n471), .ZN(new_n505));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT73), .B(G114), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(new_n472), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n501), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(KEYINPUT74), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT74), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(KEYINPUT5), .A3(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(KEYINPUT76), .B1(new_n517), .B2(G62), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT76), .ZN(new_n519));
  INV_X1    g094(.A(G62), .ZN(new_n520));
  AOI211_X1 g095(.A(new_n519), .B(new_n520), .C1(new_n514), .C2(new_n516), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G651), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT75), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT6), .B(G651), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n517), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n526), .B1(new_n517), .B2(new_n527), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n527), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n530), .A2(G88), .B1(G50), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n525), .A2(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  AND3_X1   g110(.A1(new_n515), .A2(KEYINPUT5), .A3(G543), .ZN(new_n536));
  AOI21_X1  g111(.A(G543), .B1(new_n515), .B2(KEYINPUT5), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n527), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT75), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n517), .A2(new_n526), .A3(new_n527), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n539), .A2(G89), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT7), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n532), .A2(G51), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n541), .A2(new_n542), .A3(new_n544), .A4(new_n545), .ZN(G286));
  INV_X1    g121(.A(G286), .ZN(G168));
  AOI22_X1  g122(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G651), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n539), .A2(G90), .A3(new_n540), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n532), .A2(G52), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(G171));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(new_n517), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI211_X1 g131(.A(KEYINPUT77), .B(new_n554), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n556), .B1(new_n514), .B2(new_n516), .ZN(new_n559));
  INV_X1    g134(.A(new_n554), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n557), .A2(G651), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n539), .A2(G81), .A3(new_n540), .ZN(new_n563));
  XNOR2_X1  g138(.A(KEYINPUT78), .B(G43), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n532), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  AND3_X1   g143(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G36), .ZN(new_n570));
  XOR2_X1   g145(.A(new_n570), .B(KEYINPUT79), .Z(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n569), .A2(new_n573), .ZN(G188));
  NAND2_X1  g149(.A1(new_n549), .A2(KEYINPUT6), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT6), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G651), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n575), .A2(new_n577), .A3(G53), .A4(G543), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT80), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT9), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n579), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n578), .A2(new_n579), .A3(KEYINPUT9), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n530), .A2(G91), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT81), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n585), .B1(new_n536), .B2(new_n537), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n514), .A2(KEYINPUT81), .A3(new_n516), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n586), .A2(G65), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(G78), .A2(G543), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g165(.A(KEYINPUT82), .B1(new_n590), .B2(G651), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT82), .ZN(new_n592));
  AOI211_X1 g167(.A(new_n592), .B(new_n549), .C1(new_n588), .C2(new_n589), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n584), .B1(new_n591), .B2(new_n593), .ZN(G299));
  OAI211_X1 g169(.A(new_n551), .B(new_n552), .C1(new_n549), .C2(new_n548), .ZN(G301));
  OAI21_X1  g170(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n532), .A2(G49), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n539), .A2(new_n540), .ZN(new_n598));
  INV_X1    g173(.A(G87), .ZN(new_n599));
  OAI211_X1 g174(.A(new_n596), .B(new_n597), .C1(new_n598), .C2(new_n599), .ZN(G288));
  NAND2_X1  g175(.A1(G73), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G61), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n555), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(G48), .B2(new_n532), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT83), .ZN(new_n605));
  AND3_X1   g180(.A1(new_n530), .A2(new_n605), .A3(G86), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n605), .B1(new_n530), .B2(G86), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n604), .B1(new_n606), .B2(new_n607), .ZN(G305));
  INV_X1    g183(.A(KEYINPUT84), .ZN(new_n609));
  NAND2_X1  g184(.A1(G72), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G60), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n609), .B(new_n610), .C1(new_n555), .C2(new_n611), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n611), .B1(new_n514), .B2(new_n516), .ZN(new_n613));
  INV_X1    g188(.A(new_n610), .ZN(new_n614));
  OAI21_X1  g189(.A(KEYINPUT84), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n612), .A2(G651), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n532), .A2(G47), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n539), .A2(G85), .A3(new_n540), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(G290));
  NAND2_X1  g194(.A1(G301), .A2(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n532), .A2(G54), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n539), .A2(G92), .A3(new_n540), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(KEYINPUT10), .ZN(new_n623));
  AND3_X1   g198(.A1(new_n514), .A2(KEYINPUT81), .A3(new_n516), .ZN(new_n624));
  AOI21_X1  g199(.A(KEYINPUT81), .B1(new_n514), .B2(new_n516), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT85), .B(G66), .ZN(new_n626));
  NOR3_X1   g201(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AND2_X1   g202(.A1(G79), .A2(G543), .ZN(new_n628));
  OAI21_X1  g203(.A(G651), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT10), .ZN(new_n630));
  NAND4_X1  g205(.A1(new_n539), .A2(new_n630), .A3(G92), .A4(new_n540), .ZN(new_n631));
  AND4_X1   g206(.A1(new_n621), .A2(new_n623), .A3(new_n629), .A4(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n620), .B1(new_n632), .B2(G868), .ZN(G284));
  OAI21_X1  g208(.A(new_n620), .B1(new_n632), .B2(G868), .ZN(G321));
  NAND2_X1  g209(.A1(G286), .A2(G868), .ZN(new_n635));
  INV_X1    g210(.A(G299), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(G868), .ZN(G297));
  OAI21_X1  g212(.A(new_n635), .B1(new_n636), .B2(G868), .ZN(G280));
  XNOR2_X1  g213(.A(KEYINPUT86), .B(G559), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n632), .B1(G860), .B2(new_n639), .ZN(G148));
  INV_X1    g215(.A(G868), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n566), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n632), .A2(new_n639), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT87), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n642), .B1(new_n644), .B2(new_n641), .ZN(G323));
  XNOR2_X1  g220(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g221(.A(new_n488), .ZN(new_n647));
  INV_X1    g222(.A(G123), .ZN(new_n648));
  OR3_X1    g223(.A1(new_n647), .A2(KEYINPUT88), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(KEYINPUT88), .B1(new_n647), .B2(new_n648), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n495), .A2(G135), .ZN(new_n651));
  OR2_X1    g226(.A1(G99), .A2(G2105), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n652), .B(G2104), .C1(G111), .C2(new_n472), .ZN(new_n653));
  NAND4_X1  g228(.A1(new_n649), .A2(new_n650), .A3(new_n651), .A4(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(G2096), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n471), .A2(new_n469), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT12), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT13), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2100), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n655), .A2(new_n659), .ZN(G156));
  XNOR2_X1  g235(.A(G2427), .B(G2438), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2430), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT15), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n663), .A2(G2435), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(G2435), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(KEYINPUT14), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2443), .B(G2446), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2451), .B(G2454), .Z(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT89), .B(KEYINPUT16), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1341), .B(G1348), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n672), .B(new_n673), .Z(new_n674));
  AND2_X1   g249(.A1(new_n674), .A2(G14), .ZN(G401));
  XOR2_X1   g250(.A(G2067), .B(G2678), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT90), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT91), .Z(new_n678));
  XOR2_X1   g253(.A(G2072), .B(G2078), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G2084), .B(G2090), .Z(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT92), .B(KEYINPUT17), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n679), .B(new_n683), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n680), .B(new_n682), .C1(new_n684), .C2(new_n678), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n678), .A2(new_n684), .A3(new_n681), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n677), .A2(new_n679), .A3(new_n682), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT18), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n685), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G2096), .B(G2100), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(G227));
  XOR2_X1   g266(.A(G1956), .B(G2474), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT93), .ZN(new_n693));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT94), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1971), .B(G1976), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT19), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n693), .A2(KEYINPUT94), .A3(new_n694), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n697), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT20), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n693), .A2(new_n694), .ZN(new_n704));
  AOI22_X1  g279(.A1(new_n702), .A2(new_n703), .B1(new_n700), .B2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n704), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n706), .A2(new_n699), .A3(new_n695), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n705), .B(new_n707), .C1(new_n703), .C2(new_n702), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1991), .B(G1996), .ZN(new_n711));
  INV_X1    g286(.A(G1981), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1986), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n710), .B(new_n714), .ZN(G229));
  NOR2_X1   g290(.A1(G27), .A2(G29), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G164), .B2(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G2078), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT99), .B(KEYINPUT28), .Z(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G26), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n719), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n488), .A2(G128), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n495), .A2(G140), .ZN(new_n724));
  OR2_X1    g299(.A1(G104), .A2(G2105), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n725), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT97), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n723), .A2(new_n724), .A3(KEYINPUT97), .A4(new_n726), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AND3_X1   g306(.A1(new_n731), .A2(KEYINPUT98), .A3(G29), .ZN(new_n732));
  AOI21_X1  g307(.A(KEYINPUT98), .B1(new_n731), .B2(G29), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n722), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G2067), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n495), .A2(G139), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n469), .A2(G103), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT25), .Z(new_n738));
  AOI22_X1  g313(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT100), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n736), .B(new_n738), .C1(new_n741), .C2(new_n472), .ZN(new_n742));
  MUX2_X1   g317(.A(G33), .B(new_n742), .S(G29), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2072), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n735), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G16), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G19), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n567), .B2(new_n746), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1341), .ZN(new_n749));
  AND2_X1   g324(.A1(KEYINPUT30), .A2(G28), .ZN(new_n750));
  NOR2_X1   g325(.A1(KEYINPUT30), .A2(G28), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n720), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT31), .B(G11), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n752), .B(new_n753), .C1(new_n654), .C2(new_n720), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT102), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n749), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n746), .A2(KEYINPUT23), .A3(G20), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT23), .ZN(new_n758));
  INV_X1    g333(.A(G20), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(G16), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n757), .B(new_n760), .C1(new_n636), .C2(new_n746), .ZN(new_n761));
  INV_X1    g336(.A(G1956), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n746), .A2(G4), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n632), .B2(new_n746), .ZN(new_n765));
  INV_X1    g340(.A(G1348), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n745), .A2(new_n756), .A3(new_n763), .A4(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(G29), .A2(G35), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G162), .B2(G29), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT29), .B(G2090), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(G160), .A2(G29), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT101), .B(KEYINPUT24), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G34), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n773), .B1(G29), .B2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G2084), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G2078), .B2(new_n717), .ZN(new_n779));
  INV_X1    g354(.A(G1961), .ZN(new_n780));
  OAI21_X1  g355(.A(KEYINPUT103), .B1(G5), .B2(G16), .ZN(new_n781));
  OR3_X1    g356(.A1(KEYINPUT103), .A2(G5), .A3(G16), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n781), .B(new_n782), .C1(G301), .C2(new_n746), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n779), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  OAI221_X1 g359(.A(new_n784), .B1(new_n780), .B2(new_n783), .C1(new_n777), .C2(new_n776), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n768), .A2(new_n772), .A3(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT96), .ZN(new_n787));
  INV_X1    g362(.A(G22), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(G16), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(G16), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G303), .B2(G16), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n789), .B1(new_n791), .B2(new_n787), .ZN(new_n792));
  INV_X1    g367(.A(G1971), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G16), .A2(G23), .ZN(new_n795));
  NAND2_X1  g370(.A1(G288), .A2(KEYINPUT95), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n530), .A2(G87), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT95), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n797), .A2(new_n798), .A3(new_n596), .A4(new_n597), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n795), .B1(new_n800), .B2(G16), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT33), .B(G1976), .Z(new_n802));
  XOR2_X1   g377(.A(new_n801), .B(new_n802), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n746), .A2(G6), .ZN(new_n804));
  INV_X1    g379(.A(new_n604), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n530), .A2(G86), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(KEYINPUT83), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n530), .A2(new_n605), .A3(G86), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n804), .B1(new_n809), .B2(new_n746), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT32), .B(G1981), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n794), .A2(new_n803), .A3(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT34), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT36), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n488), .A2(G119), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n495), .A2(G131), .ZN(new_n818));
  OAI21_X1  g393(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n472), .A2(G107), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n817), .B(new_n818), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  MUX2_X1   g396(.A(G25), .B(new_n821), .S(G29), .Z(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT35), .B(G1991), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n822), .B(new_n823), .Z(new_n824));
  INV_X1    g399(.A(G290), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G16), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G16), .B2(G24), .ZN(new_n827));
  INV_X1    g402(.A(G1986), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n824), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n828), .B2(new_n827), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n815), .A2(new_n816), .A3(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n816), .B1(new_n815), .B2(new_n830), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n718), .B(new_n786), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n746), .A2(G21), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(G168), .B2(new_n746), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G1966), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n495), .A2(G141), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n488), .A2(G129), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n469), .A2(G105), .ZN(new_n840));
  NAND3_X1  g415(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT26), .Z(new_n842));
  NAND4_X1  g417(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(G29), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(G29), .B2(G32), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT27), .B(G1996), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n834), .A2(new_n837), .A3(new_n848), .ZN(G311));
  INV_X1    g424(.A(new_n786), .ZN(new_n850));
  INV_X1    g425(.A(new_n833), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n850), .B1(new_n851), .B2(new_n831), .ZN(new_n852));
  INV_X1    g427(.A(new_n837), .ZN(new_n853));
  INV_X1    g428(.A(new_n848), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .A4(new_n718), .ZN(G150));
  INV_X1    g430(.A(G67), .ZN(new_n856));
  INV_X1    g431(.A(G80), .ZN(new_n857));
  OAI22_X1  g432(.A1(new_n555), .A2(new_n856), .B1(new_n857), .B2(new_n512), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(KEYINPUT104), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT104), .ZN(new_n860));
  OAI221_X1 g435(.A(new_n860), .B1(new_n857), .B2(new_n512), .C1(new_n555), .C2(new_n856), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n859), .A2(G651), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n539), .A2(G93), .A3(new_n540), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT105), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n532), .A2(G55), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n864), .B1(new_n863), .B2(new_n865), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n862), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  XOR2_X1   g443(.A(KEYINPUT106), .B(G860), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT37), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n567), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n566), .B(new_n862), .C1(new_n866), .C2(new_n867), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT39), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n632), .A2(G559), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT38), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n875), .B(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n871), .B1(new_n878), .B2(new_n869), .ZN(G145));
  AOI21_X1  g454(.A(new_n731), .B1(new_n742), .B2(KEYINPUT108), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n742), .A2(new_n731), .A3(KEYINPUT108), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n510), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n501), .A2(new_n505), .A3(new_n509), .A4(KEYINPUT107), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n881), .A2(new_n882), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n886), .ZN(new_n888));
  INV_X1    g463(.A(new_n882), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n888), .B1(new_n889), .B2(new_n880), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n843), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n821), .B(new_n657), .Z(new_n893));
  NOR2_X1   g468(.A1(new_n472), .A2(G118), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n894), .B(KEYINPUT109), .Z(new_n895));
  OAI211_X1 g470(.A(new_n895), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n495), .A2(G142), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n488), .A2(G130), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n893), .B(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n887), .A2(new_n890), .A3(new_n844), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n892), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT110), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n892), .A2(new_n901), .ZN(new_n904));
  INV_X1    g479(.A(new_n900), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI211_X1 g481(.A(KEYINPUT110), .B(new_n900), .C1(new_n892), .C2(new_n901), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n902), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  XOR2_X1   g483(.A(G162), .B(G160), .Z(new_n909));
  XOR2_X1   g484(.A(new_n909), .B(new_n654), .Z(new_n910));
  AOI21_X1  g485(.A(G37), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n900), .B1(new_n892), .B2(new_n901), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(new_n903), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n902), .B(KEYINPUT111), .ZN(new_n914));
  INV_X1    g489(.A(new_n910), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g493(.A(KEYINPUT112), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n874), .B(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(new_n644), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT41), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n632), .A2(G299), .ZN(new_n923));
  INV_X1    g498(.A(G65), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n624), .A2(new_n625), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n589), .ZN(new_n926));
  OAI21_X1  g501(.A(G651), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n592), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n590), .A2(KEYINPUT82), .A3(G651), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n623), .A2(new_n629), .A3(new_n621), .A4(new_n631), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n584), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT113), .B1(new_n923), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT113), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n934), .B1(new_n636), .B2(new_n931), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n922), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n923), .A2(new_n932), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT41), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n921), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(new_n937), .B2(new_n921), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n800), .A2(new_n809), .ZN(new_n944));
  NAND3_X1  g519(.A1(G305), .A2(new_n796), .A3(new_n799), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n618), .A2(new_n617), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n525), .A2(new_n947), .A3(new_n533), .A4(new_n616), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n549), .B1(new_n522), .B2(new_n523), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n532), .A2(G50), .ZN(new_n950));
  INV_X1    g525(.A(G88), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n950), .B1(new_n598), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(G290), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT114), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n948), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n954), .B1(new_n948), .B2(new_n953), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n946), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n948), .A2(new_n953), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT114), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n948), .A2(new_n953), .A3(new_n954), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n959), .A2(new_n960), .B1(new_n945), .B2(new_n944), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n957), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g537(.A(new_n962), .B(KEYINPUT42), .Z(new_n963));
  AND2_X1   g538(.A1(new_n943), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n943), .A2(new_n963), .ZN(new_n965));
  OAI21_X1  g540(.A(G868), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n868), .A2(new_n641), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(G295));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n967), .ZN(G331));
  XNOR2_X1  g544(.A(G171), .B(G286), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n863), .A2(new_n865), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT105), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n566), .B1(new_n974), .B2(new_n862), .ZN(new_n975));
  INV_X1    g550(.A(new_n873), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n970), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(G301), .B(G286), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n872), .A2(new_n978), .A3(new_n873), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT41), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n938), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n933), .A2(new_n935), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n982), .B(new_n962), .C1(new_n983), .C2(new_n981), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n936), .A2(new_n939), .A3(new_n980), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n977), .A2(new_n938), .A3(new_n979), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT115), .ZN(new_n988));
  INV_X1    g563(.A(new_n962), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n988), .B1(new_n987), .B2(new_n989), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n984), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT43), .B1(new_n992), .B2(G37), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n985), .A2(new_n962), .A3(new_n986), .ZN(new_n994));
  INV_X1    g569(.A(G37), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(new_n990), .B2(new_n991), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n993), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n999));
  NOR2_X1   g574(.A1(KEYINPUT43), .A2(G37), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n984), .B(new_n1000), .C1(new_n990), .C2(new_n991), .ZN(new_n1001));
  AOI211_X1 g576(.A(KEYINPUT116), .B(KEYINPUT44), .C1(new_n999), .C2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n994), .A2(new_n995), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n987), .A2(new_n989), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT115), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT43), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1001), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1003), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n998), .B1(new_n1002), .B2(new_n1012), .ZN(G397));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n1014));
  AOI22_X1  g589(.A1(new_n495), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT70), .B1(new_n484), .B2(G2105), .ZN(new_n1016));
  AOI211_X1 g591(.A(new_n476), .B(new_n472), .C1(new_n482), .C2(new_n483), .ZN(new_n1017));
  OAI211_X1 g592(.A(G40), .B(new_n1015), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n1020));
  INV_X1    g595(.A(G1384), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1020), .B1(new_n510), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G114), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1024), .A2(KEYINPUT73), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(KEYINPUT73), .ZN(new_n1026));
  OAI21_X1  g601(.A(G2105), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n1027), .A2(new_n507), .B1(new_n504), .B2(new_n471), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1384), .B1(new_n1028), .B2(new_n501), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n1020), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1019), .A2(new_n1023), .A3(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(G2084), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT45), .B1(new_n510), .B2(new_n1021), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1018), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1029), .A2(KEYINPUT45), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1966), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(G8), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  XOR2_X1   g612(.A(KEYINPUT118), .B(G8), .Z(new_n1038));
  NAND2_X1  g613(.A1(G286), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1014), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1014), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1042));
  INV_X1    g617(.A(G1966), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(G2084), .B2(new_n1031), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1041), .B1(new_n1045), .B2(new_n1038), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT125), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1039), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1047), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n510), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1050), .A2(new_n1018), .A3(new_n1022), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1042), .A2(new_n1043), .B1(new_n1051), .B2(new_n777), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1052), .A2(KEYINPUT125), .A3(new_n1039), .ZN(new_n1053));
  OAI22_X1  g628(.A1(new_n1040), .A2(new_n1046), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1054));
  OR2_X1    g629(.A1(new_n1054), .A2(KEYINPUT62), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT49), .ZN(new_n1056));
  NOR2_X1   g631(.A1(G305), .A2(G1981), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n712), .B1(new_n806), .B2(new_n604), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n809), .A2(new_n712), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1058), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(KEYINPUT49), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n510), .A2(new_n1021), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1038), .B1(new_n1018), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT119), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1066), .B(new_n1038), .C1(new_n1018), .C2(new_n1063), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1059), .A2(new_n1062), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1068), .ZN(new_n1071));
  INV_X1    g646(.A(G1976), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1072), .B1(new_n796), .B2(new_n799), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1070), .B(KEYINPUT52), .C1(new_n1071), .C2(new_n1073), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1065), .A2(new_n1067), .B1(new_n800), .B2(G1976), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT120), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(G288), .A2(new_n1072), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1069), .A2(new_n1074), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(G303), .A2(G8), .ZN(new_n1081));
  XOR2_X1   g656(.A(new_n1081), .B(KEYINPUT55), .Z(new_n1082));
  INV_X1    g657(.A(new_n1038), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n886), .A2(KEYINPUT45), .A3(new_n1021), .ZN(new_n1084));
  AOI21_X1  g659(.A(G1971), .B1(new_n1084), .B2(new_n1034), .ZN(new_n1085));
  NOR4_X1   g660(.A1(new_n1050), .A2(new_n1018), .A3(new_n1022), .A4(G2090), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1083), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT121), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1082), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1081), .B(KEYINPUT55), .ZN(new_n1092));
  INV_X1    g667(.A(G8), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1092), .A2(new_n1093), .A3(new_n1087), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1080), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT126), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1042), .B2(G2078), .ZN(new_n1097));
  INV_X1    g672(.A(G2078), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1034), .A2(KEYINPUT126), .A3(new_n1098), .A4(new_n1035), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1097), .A2(KEYINPUT53), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1084), .A2(new_n1034), .A3(new_n1098), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1101), .A2(new_n1102), .B1(new_n780), .B2(new_n1031), .ZN(new_n1103));
  AOI21_X1  g678(.A(G301), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1054), .A2(KEYINPUT62), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1055), .A2(new_n1095), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G288), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1069), .A2(new_n1072), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1071), .B1(new_n1108), .B2(new_n1060), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1084), .A2(new_n1034), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n793), .ZN(new_n1111));
  INV_X1    g686(.A(G2090), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1051), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1111), .A2(new_n1088), .A3(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1114), .A2(new_n1090), .A3(new_n1038), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n1092), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT63), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1052), .A2(G286), .A3(new_n1083), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1094), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AND4_X1   g696(.A1(new_n1069), .A2(new_n1074), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1109), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1087), .A2(new_n1093), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1118), .B1(new_n1082), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT63), .B1(new_n1080), .B2(new_n1125), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1106), .A2(new_n1123), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1122), .A2(new_n1054), .A3(new_n1116), .A4(new_n1120), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT54), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT45), .B1(new_n886), .B2(new_n1021), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT45), .ZN(new_n1132));
  AOI211_X1 g707(.A(new_n1132), .B(G1384), .C1(new_n884), .C2(new_n885), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n477), .A2(new_n472), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1102), .A2(G2078), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1134), .A2(new_n1015), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(G40), .ZN(new_n1139));
  OAI211_X1 g714(.A(G301), .B(new_n1103), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1130), .B1(new_n1141), .B2(new_n1104), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1103), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(G171), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1100), .A2(new_n1103), .A3(G301), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1144), .A2(KEYINPUT54), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1142), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1128), .B1(new_n1129), .B2(new_n1147), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1140), .B1(new_n1149), .B2(G301), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1130), .B1(new_n1143), .B2(G171), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1150), .A2(new_n1130), .B1(new_n1151), .B2(new_n1145), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1152), .A2(new_n1095), .A3(KEYINPUT127), .A4(new_n1054), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1148), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT122), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1031), .A2(new_n762), .ZN(new_n1156));
  XNOR2_X1  g731(.A(KEYINPUT56), .B(G2072), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1084), .A2(new_n1034), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT57), .ZN(new_n1161));
  XNOR2_X1  g736(.A(G299), .B(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1155), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g738(.A(G299), .B(KEYINPUT57), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1164), .A2(KEYINPUT122), .A3(new_n1159), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(G2067), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1018), .A2(new_n1063), .ZN(new_n1168));
  AOI22_X1  g743(.A1(new_n1031), .A2(new_n766), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n1169), .A2(new_n931), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1166), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1164), .A2(new_n1159), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT61), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1175), .B1(new_n1176), .B2(new_n1172), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1169), .B(new_n931), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT60), .ZN(new_n1179));
  XOR2_X1   g754(.A(KEYINPUT123), .B(KEYINPUT58), .Z(new_n1180));
  XNOR2_X1  g755(.A(new_n1180), .B(G1341), .ZN(new_n1181));
  OAI22_X1  g756(.A1(new_n1110), .A2(G1996), .B1(new_n1168), .B2(new_n1181), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1182), .A2(KEYINPUT59), .A3(new_n567), .ZN(new_n1183));
  AOI21_X1  g758(.A(KEYINPUT59), .B1(new_n1182), .B2(new_n567), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT60), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1169), .A2(new_n1186), .A3(new_n632), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1177), .A2(new_n1179), .A3(new_n1185), .A4(new_n1187), .ZN(new_n1188));
  AOI211_X1 g763(.A(new_n1175), .B(new_n1172), .C1(new_n1163), .C2(new_n1165), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1174), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT124), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  OAI211_X1 g767(.A(new_n1174), .B(KEYINPUT124), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1127), .B1(new_n1154), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(KEYINPUT107), .B1(new_n1028), .B2(new_n501), .ZN(new_n1196));
  INV_X1    g771(.A(new_n885), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1021), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1198), .A2(new_n1132), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1199), .A2(new_n1018), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n731), .B(new_n1167), .ZN(new_n1201));
  INV_X1    g776(.A(G1996), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n843), .B(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n821), .B(new_n823), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1200), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(new_n1200), .ZN(new_n1207));
  NOR3_X1   g782(.A1(new_n1207), .A2(G1986), .A3(G290), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n825), .A2(new_n828), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1208), .B1(new_n1200), .B2(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n1210), .B(KEYINPUT117), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1195), .A2(new_n1206), .A3(new_n1211), .ZN(new_n1212));
  OR2_X1    g787(.A1(new_n821), .A2(new_n823), .ZN(new_n1213));
  OAI22_X1  g788(.A1(new_n1204), .A2(new_n1213), .B1(G2067), .B2(new_n731), .ZN(new_n1214));
  AND2_X1   g789(.A1(new_n1214), .A2(new_n1200), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1207), .B1(new_n1201), .B2(new_n844), .ZN(new_n1216));
  AND3_X1   g791(.A1(new_n1200), .A2(KEYINPUT46), .A3(new_n1202), .ZN(new_n1217));
  AOI21_X1  g792(.A(KEYINPUT46), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1218));
  NOR3_X1   g793(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  XNOR2_X1  g794(.A(new_n1219), .B(KEYINPUT47), .ZN(new_n1220));
  XOR2_X1   g795(.A(new_n1208), .B(KEYINPUT48), .Z(new_n1221));
  AOI211_X1 g796(.A(new_n1215), .B(new_n1220), .C1(new_n1206), .C2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1212), .A2(new_n1222), .ZN(G329));
  assign    G231 = 1'b0;
  AOI211_X1 g798(.A(new_n466), .B(G229), .C1(new_n911), .C2(new_n916), .ZN(new_n1225));
  NOR2_X1   g799(.A1(G401), .A2(G227), .ZN(new_n1226));
  AND3_X1   g800(.A1(new_n1225), .A2(new_n1010), .A3(new_n1226), .ZN(G308));
  NAND3_X1  g801(.A1(new_n1225), .A2(new_n1010), .A3(new_n1226), .ZN(G225));
endmodule


