//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n210, new_n211, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1251, new_n1252, new_n1253, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1319, new_n1320, new_n1321;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  NOR2_X1   g0009(.A1(G97), .A2(G107), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G87), .ZN(G355));
  NAND2_X1  g0012(.A1(G1), .A2(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n216), .A2(KEYINPUT0), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n206), .A2(new_n207), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n216), .A2(KEYINPUT0), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n217), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT65), .ZN(new_n225));
  INV_X1    g0025(.A(G226), .ZN(new_n226));
  INV_X1    g0026(.A(G97), .ZN(new_n227));
  INV_X1    g0027(.A(G257), .ZN(new_n228));
  OAI22_X1  g0028(.A1(new_n207), .A2(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(G116), .B2(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT66), .B(G244), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G77), .ZN(new_n232));
  AOI22_X1  g0032(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  AOI22_X1  g0034(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT67), .ZN(new_n236));
  OAI21_X1  g0036(.A(new_n213), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  OR2_X1    g0037(.A1(new_n237), .A2(KEYINPUT1), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n237), .A2(KEYINPUT1), .ZN(new_n239));
  AND3_X1   g0039(.A1(new_n225), .A2(new_n238), .A3(new_n239), .ZN(G361));
  XOR2_X1   g0040(.A(G238), .B(G244), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G232), .ZN(new_n242));
  XOR2_X1   g0042(.A(KEYINPUT2), .B(G226), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G264), .B(G270), .Z(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G358));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT68), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G50), .B(G68), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G58), .B(G77), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  INV_X1    g0056(.A(G169), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT3), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n259), .A2(new_n261), .A3(G223), .A4(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT79), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT3), .B(G33), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n266), .A2(KEYINPUT79), .A3(G223), .A4(new_n262), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(G226), .A3(G1698), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G87), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n265), .A2(new_n267), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  AND2_X1   g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(new_n219), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT81), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  OAI211_X1 g0075(.A(G1), .B(G13), .C1(new_n258), .C2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G1), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n277), .B1(G41), .B2(G45), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(G232), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT80), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n276), .A2(KEYINPUT80), .A3(G232), .A4(new_n278), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT69), .ZN(new_n283));
  OAI21_X1  g0083(.A(G274), .B1(new_n271), .B2(new_n219), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n283), .B1(new_n284), .B2(new_n278), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  AOI21_X1  g0086(.A(G1), .B1(new_n275), .B2(new_n286), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n276), .A2(KEYINPUT69), .A3(new_n287), .A4(G274), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n281), .A2(new_n282), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  AND3_X1   g0089(.A1(new_n273), .A2(new_n274), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n274), .B1(new_n273), .B2(new_n289), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n257), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G58), .A2(G68), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n203), .A2(new_n205), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G20), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G159), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT78), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT7), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(new_n266), .B2(G20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n259), .A2(new_n261), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(KEYINPUT7), .A3(new_n220), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G68), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT78), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n295), .A2(new_n306), .A3(new_n297), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n299), .A2(new_n305), .A3(KEYINPUT16), .A4(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT16), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n202), .B1(new_n301), .B2(new_n303), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n309), .B1(new_n310), .B2(new_n298), .ZN(new_n311));
  NAND3_X1  g0111(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n219), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n308), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(KEYINPUT71), .A2(G58), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT8), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(new_n277), .B2(G20), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n277), .A2(G13), .A3(G20), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT72), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT72), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n321), .A2(new_n277), .A3(G13), .A4(G20), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n313), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n320), .A2(new_n322), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n318), .A2(new_n323), .B1(new_n324), .B2(new_n317), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n314), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n273), .A2(new_n289), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G179), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n292), .A2(new_n326), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT18), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT18), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n292), .A2(new_n326), .A3(new_n333), .A4(new_n330), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT82), .ZN(new_n336));
  INV_X1    g0136(.A(G200), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n290), .B2(new_n291), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n327), .A2(G190), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n326), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n341), .A2(KEYINPUT17), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(KEYINPUT17), .B1(new_n341), .B2(new_n342), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n336), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT17), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n327), .A2(KEYINPUT81), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n273), .A2(new_n274), .A3(new_n289), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n339), .B1(new_n349), .B2(new_n337), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n346), .B1(new_n350), .B2(new_n326), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n341), .A2(KEYINPUT17), .A3(new_n342), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(KEYINPUT82), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n335), .B1(new_n345), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT76), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n258), .A2(G20), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n356), .A2(G77), .B1(G20), .B2(new_n202), .ZN(new_n357));
  INV_X1    g0157(.A(new_n296), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n357), .B1(new_n207), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n359), .A2(KEYINPUT11), .A3(new_n313), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT11), .B1(new_n359), .B2(new_n313), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n355), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n362), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(KEYINPUT76), .A3(new_n360), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n320), .A2(new_n322), .ZN(new_n366));
  OR3_X1    g0166(.A1(new_n366), .A2(KEYINPUT12), .A3(G68), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT12), .B1(new_n366), .B2(G68), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n202), .B1(new_n277), .B2(G20), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n367), .A2(new_n368), .B1(new_n323), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n363), .A2(new_n365), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n371), .B(KEYINPUT77), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT75), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n285), .A2(new_n288), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n266), .A2(G226), .A3(new_n262), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n266), .A2(G232), .A3(G1698), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G33), .A2(G97), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n373), .A2(new_n374), .B1(new_n378), .B2(new_n272), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n285), .A2(KEYINPUT75), .A3(new_n288), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n272), .A2(new_n287), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(G238), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT13), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT13), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n379), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(G179), .A3(new_n387), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n379), .A2(new_n383), .A3(new_n386), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n386), .B1(new_n379), .B2(new_n383), .ZN(new_n390));
  OAI21_X1  g0190(.A(G169), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n388), .B1(new_n391), .B2(KEYINPUT14), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT14), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n385), .A2(new_n387), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n393), .B1(new_n394), .B2(G169), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n372), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n385), .A2(G190), .A3(new_n387), .ZN(new_n397));
  INV_X1    g0197(.A(new_n371), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n337), .B1(new_n385), .B2(new_n387), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n266), .A2(G222), .A3(new_n262), .ZN(new_n403));
  INV_X1    g0203(.A(G77), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n266), .A2(G1698), .ZN(new_n405));
  INV_X1    g0205(.A(G223), .ZN(new_n406));
  OAI221_X1 g0206(.A(new_n403), .B1(new_n404), .B2(new_n266), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n272), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n226), .A2(KEYINPUT70), .ZN(new_n409));
  OR2_X1    g0209(.A1(new_n226), .A2(KEYINPUT70), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n381), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n374), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(G200), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n408), .A2(new_n412), .A3(G190), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n313), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n316), .A2(new_n356), .B1(G150), .B2(new_n296), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n208), .A2(G20), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n207), .B1(new_n277), .B2(G20), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n323), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(G50), .B2(new_n366), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n420), .A2(new_n423), .A3(KEYINPUT9), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT9), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n418), .A2(new_n419), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n313), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n207), .A2(new_n324), .B1(new_n323), .B2(new_n421), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n425), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n416), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n414), .A2(KEYINPUT74), .A3(new_n415), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT10), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n404), .B1(new_n277), .B2(G20), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n404), .A2(new_n324), .B1(new_n323), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g0237(.A(KEYINPUT8), .B(G58), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n438), .A2(new_n358), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n220), .A2(new_n404), .ZN(new_n440));
  INV_X1    g0240(.A(G87), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n441), .A2(KEYINPUT15), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(KEYINPUT15), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT73), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT15), .B(G87), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT73), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  AOI211_X1 g0249(.A(new_n439), .B(new_n440), .C1(new_n449), .C2(new_n356), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n437), .B1(new_n450), .B2(new_n417), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n266), .A2(G232), .A3(new_n262), .ZN(new_n453));
  INV_X1    g0253(.A(G107), .ZN(new_n454));
  INV_X1    g0254(.A(G238), .ZN(new_n455));
  OAI221_X1 g0255(.A(new_n453), .B1(new_n454), .B2(new_n266), .C1(new_n405), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n272), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n285), .A2(new_n288), .B1(new_n381), .B2(new_n231), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G200), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n457), .A2(new_n458), .A3(G190), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n452), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(new_n257), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n457), .A2(new_n458), .A3(new_n329), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n451), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n432), .B(new_n433), .C1(new_n416), .C2(new_n430), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n413), .A2(new_n257), .B1(new_n427), .B2(new_n428), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(G179), .B2(new_n413), .ZN(new_n469));
  AND4_X1   g0269(.A1(new_n435), .A2(new_n466), .A3(new_n467), .A4(new_n469), .ZN(new_n470));
  AND4_X1   g0270(.A1(new_n354), .A2(new_n396), .A3(new_n402), .A4(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT85), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n286), .A2(G1), .ZN(new_n473));
  NAND2_X1  g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(KEYINPUT5), .A2(G41), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(new_n284), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n277), .A2(G45), .ZN(new_n479));
  INV_X1    g0279(.A(new_n476), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n479), .B1(new_n480), .B2(new_n474), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n481), .A2(new_n228), .A3(new_n272), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n259), .A2(new_n261), .A3(G244), .A4(new_n262), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n266), .A2(KEYINPUT4), .A3(G244), .A4(new_n262), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G283), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n266), .A2(G250), .A3(G1698), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n485), .A2(new_n486), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  AOI211_X1 g0289(.A(new_n478), .B(new_n482), .C1(new_n489), .C2(new_n272), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n472), .B1(new_n490), .B2(new_n337), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT83), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n358), .A2(new_n404), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT6), .ZN(new_n495));
  AND2_X1   g0295(.A1(G97), .A2(G107), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(new_n210), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n454), .A2(KEYINPUT6), .A3(G97), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n492), .B(new_n494), .C1(new_n499), .C2(new_n220), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n304), .A2(G107), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n220), .B1(new_n497), .B2(new_n498), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT83), .B1(new_n502), .B2(new_n493), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n500), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT84), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n258), .A2(G1), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n227), .B1(new_n323), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n366), .A2(new_n227), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n505), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  AOI211_X1 g0311(.A(new_n506), .B(new_n313), .C1(new_n320), .C2(new_n322), .ZN(new_n512));
  OAI211_X1 g0312(.A(KEYINPUT84), .B(new_n509), .C1(new_n512), .C2(new_n227), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n504), .A2(new_n313), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n489), .A2(new_n272), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n481), .A2(G274), .A3(new_n276), .ZN(new_n516));
  INV_X1    g0316(.A(new_n482), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(KEYINPUT85), .A3(G200), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n490), .A2(G190), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n491), .A2(new_n514), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n259), .A2(new_n261), .A3(G238), .A4(new_n262), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n259), .A2(new_n261), .A3(G244), .A4(G1698), .ZN(new_n523));
  INV_X1    g0323(.A(G116), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n522), .B(new_n523), .C1(new_n258), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n272), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n276), .A2(G274), .A3(new_n473), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n276), .A2(G250), .A3(new_n479), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT86), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n529), .B1(new_n527), .B2(new_n528), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n526), .B(G190), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT19), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n220), .B1(new_n377), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(G87), .B2(new_n211), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n259), .A2(new_n261), .A3(new_n220), .A4(G68), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n220), .A2(G33), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n533), .B1(new_n537), .B2(new_n227), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n313), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n448), .A2(new_n324), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n323), .A2(G87), .A3(new_n507), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n526), .B1(new_n530), .B2(new_n531), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n543), .B1(G200), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n539), .A2(new_n313), .B1(new_n448), .B2(new_n324), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n449), .A2(new_n512), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n544), .A2(new_n257), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n526), .B(new_n329), .C1(new_n530), .C2(new_n531), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n532), .A2(new_n545), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n504), .A2(new_n313), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n511), .A2(new_n513), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n490), .A2(new_n329), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n518), .A2(new_n257), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n521), .A2(new_n550), .A3(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n366), .A2(G116), .A3(new_n417), .A4(new_n507), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n320), .A2(new_n524), .A3(new_n322), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n312), .A2(new_n219), .B1(G20), .B2(new_n524), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n487), .B(new_n220), .C1(G33), .C2(new_n227), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n561), .A2(KEYINPUT20), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT20), .B1(new_n561), .B2(new_n562), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(KEYINPUT87), .B1(new_n560), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n564), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n561), .A2(KEYINPUT20), .A3(new_n562), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT87), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(new_n558), .A4(new_n559), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n481), .A2(new_n272), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n478), .B1(new_n573), .B2(G270), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n260), .A2(G33), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n576));
  OAI21_X1  g0376(.A(G303), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n259), .A2(new_n261), .A3(G264), .A4(G1698), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n259), .A2(new_n261), .A3(G257), .A4(new_n262), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n272), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n257), .B1(new_n574), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n572), .A2(KEYINPUT21), .A3(new_n582), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n580), .A2(new_n272), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n477), .A2(G270), .A3(new_n276), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n516), .A2(new_n585), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n584), .A2(new_n329), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n572), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT21), .B1(new_n572), .B2(new_n582), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n337), .B1(new_n574), .B2(new_n581), .ZN(new_n591));
  INV_X1    g0391(.A(G190), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n584), .A2(new_n592), .A3(new_n586), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n572), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n589), .A2(new_n590), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT23), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n220), .B2(G107), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n454), .A2(KEYINPUT23), .A3(G20), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n597), .A2(new_n598), .B1(new_n356), .B2(G116), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n259), .A2(new_n261), .A3(new_n220), .A4(G87), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT22), .ZN(new_n601));
  OAI21_X1  g0401(.A(KEYINPUT89), .B1(new_n601), .B2(KEYINPUT88), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT88), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT89), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n604), .A3(KEYINPUT22), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n600), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n600), .A2(new_n606), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n599), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT90), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT24), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n599), .ZN(new_n613));
  AND4_X1   g0413(.A1(new_n220), .A2(new_n259), .A3(new_n261), .A4(G87), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n602), .A2(new_n605), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n600), .A2(new_n606), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n613), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(KEYINPUT24), .B1(new_n618), .B2(KEYINPUT90), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n609), .A2(new_n610), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n313), .B(new_n612), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n366), .A2(G107), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n622), .B(KEYINPUT25), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n512), .A2(G107), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n478), .B1(new_n573), .B2(G264), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n259), .A2(new_n261), .A3(G257), .A4(G1698), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n259), .A2(new_n261), .A3(G250), .A4(new_n262), .ZN(new_n629));
  NAND2_X1  g0429(.A1(G33), .A2(G294), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n272), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n627), .A2(new_n592), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n477), .A2(G264), .A3(new_n276), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n632), .A2(new_n516), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n633), .B1(new_n635), .B2(G200), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n621), .A2(new_n626), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n627), .A2(G179), .A3(new_n632), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n257), .B1(new_n627), .B2(new_n632), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n638), .B1(new_n639), .B2(KEYINPUT91), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT91), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n635), .A2(new_n641), .A3(G179), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n621), .A2(new_n626), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n637), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n471), .A2(new_n557), .A3(new_n595), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g0445(.A(new_n645), .B(KEYINPUT92), .ZN(G372));
  INV_X1    g0446(.A(new_n469), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n345), .A2(new_n353), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT94), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n396), .B(new_n649), .C1(new_n401), .C2(new_n465), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n465), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n402), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n649), .B1(new_n653), .B2(new_n396), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n332), .B(new_n334), .C1(new_n651), .C2(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n435), .A2(new_n467), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n647), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n546), .A2(new_n547), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n527), .A2(new_n528), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(KEYINPUT86), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n660), .A2(new_n661), .B1(new_n272), .B2(new_n525), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n658), .B(new_n549), .C1(new_n662), .C2(G169), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n665), .A2(KEYINPUT26), .A3(new_n550), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n668), .B(new_n532), .C1(new_n662), .C2(new_n337), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n663), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n667), .B1(new_n556), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n664), .B1(new_n666), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n621), .A2(new_n626), .A3(new_n636), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n521), .A2(new_n550), .A3(new_n673), .A4(new_n556), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n574), .A2(G179), .A3(new_n581), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n566), .B2(new_n571), .ZN(new_n677));
  OAI21_X1  g0477(.A(G169), .B1(new_n584), .B2(new_n586), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n571), .B2(new_n566), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n677), .B1(new_n679), .B2(KEYINPUT21), .ZN(new_n680));
  INV_X1    g0480(.A(new_n590), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n611), .B1(new_n609), .B2(new_n610), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n610), .B2(new_n609), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n612), .A2(new_n313), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n625), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n640), .A2(new_n642), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n680), .B(new_n681), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(KEYINPUT93), .B1(new_n675), .B2(new_n687), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n643), .A2(new_n589), .A3(new_n590), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT93), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n689), .A2(new_n674), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n672), .B1(new_n688), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n471), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n657), .A2(new_n693), .ZN(G369));
  NAND2_X1  g0494(.A1(new_n680), .A2(new_n681), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n277), .A2(new_n220), .A3(G13), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G213), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G343), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n572), .A2(new_n701), .ZN(new_n702));
  MUX2_X1   g0502(.A(new_n695), .B(new_n595), .S(new_n702), .Z(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n701), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n644), .B1(new_n685), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n643), .A2(new_n701), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n701), .B1(new_n680), .B2(new_n681), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n644), .ZN(new_n712));
  INV_X1    g0512(.A(new_n643), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(new_n701), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n710), .A2(new_n715), .ZN(G399));
  INV_X1    g0516(.A(new_n214), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(G41), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n211), .A2(G87), .A3(G116), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(G1), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n218), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(new_n719), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT28), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n675), .A2(new_n687), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n701), .B1(new_n725), .B2(new_n672), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT29), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT26), .B1(new_n665), .B2(new_n550), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n556), .A2(new_n670), .A3(new_n667), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n663), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n690), .B1(new_n689), .B2(new_n674), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n557), .A2(new_n687), .A3(KEYINPUT93), .A4(new_n673), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(new_n701), .ZN(new_n734));
  XOR2_X1   g0534(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n735));
  OAI21_X1  g0535(.A(new_n727), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n557), .A2(new_n595), .A3(new_n644), .A4(new_n706), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n482), .B1(new_n489), .B2(new_n272), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n587), .A2(new_n738), .A3(new_n662), .A4(new_n635), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n627), .A2(new_n632), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n544), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n743), .A2(KEYINPUT30), .A3(new_n738), .A4(new_n587), .ZN(new_n744));
  AOI21_X1  g0544(.A(G179), .B1(new_n574), .B2(new_n581), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n518), .A2(new_n544), .A3(new_n745), .A4(new_n742), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n741), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n701), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT31), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n747), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n737), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G330), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n736), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n724), .B1(new_n755), .B2(G1), .ZN(G364));
  NAND2_X1  g0556(.A1(new_n220), .A2(G13), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n277), .B1(new_n758), .B2(G45), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n718), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n705), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(G330), .B2(new_n703), .ZN(new_n763));
  INV_X1    g0563(.A(new_n761), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n219), .B1(G20), .B2(new_n257), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n255), .A2(G45), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT97), .Z(new_n772));
  NOR2_X1   g0572(.A1(new_n717), .A2(new_n266), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n772), .B(new_n773), .C1(G45), .C2(new_n722), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n717), .A2(new_n302), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT96), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n776), .A2(G355), .B1(new_n524), .B2(new_n717), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n770), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n220), .A2(G179), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(new_n592), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n454), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n220), .A2(new_n329), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G190), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n592), .A2(G179), .A3(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n220), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n785), .A2(new_n202), .B1(new_n227), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n783), .A2(new_n592), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n781), .B(new_n788), .C1(G50), .C2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G190), .A2(G200), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n779), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G159), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n794), .A2(KEYINPUT32), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n779), .A2(G190), .A3(G200), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n441), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n794), .B2(KEYINPUT32), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n782), .A2(new_n791), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n266), .B1(new_n799), .B2(new_n404), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n782), .A2(G190), .A3(new_n337), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n800), .B1(G58), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n790), .A2(new_n795), .A3(new_n798), .A4(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G322), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G311), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n302), .B1(new_n799), .B2(new_n807), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n806), .B(new_n808), .C1(G329), .C2(new_n793), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n789), .A2(G326), .ZN(new_n810));
  XNOR2_X1  g0610(.A(KEYINPUT33), .B(G317), .ZN(new_n811));
  INV_X1    g0611(.A(new_n796), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n784), .A2(new_n811), .B1(new_n812), .B2(G303), .ZN(new_n813));
  INV_X1    g0613(.A(new_n787), .ZN(new_n814));
  INV_X1    g0614(.A(new_n780), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n814), .A2(G294), .B1(new_n815), .B2(G283), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n809), .A2(new_n810), .A3(new_n813), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n804), .A2(new_n817), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n764), .B(new_n778), .C1(new_n768), .C2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n767), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n819), .B1(new_n703), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n763), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(G396));
  NOR2_X1   g0623(.A1(new_n465), .A2(new_n701), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n462), .B1(new_n452), .B2(new_n706), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n824), .B1(new_n825), .B2(new_n465), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n734), .B(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n761), .B1(new_n827), .B2(new_n753), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n753), .B2(new_n827), .ZN(new_n829));
  AOI22_X1  g0629(.A1(G97), .A2(new_n814), .B1(new_n789), .B2(G303), .ZN(new_n830));
  INV_X1    g0630(.A(new_n799), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n266), .B1(new_n831), .B2(G116), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n802), .A2(G294), .B1(new_n793), .B2(G311), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n830), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n780), .A2(new_n441), .ZN(new_n835));
  INV_X1    g0635(.A(G283), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n785), .A2(new_n836), .B1(new_n796), .B2(new_n454), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT98), .Z(new_n839));
  AOI22_X1  g0639(.A1(new_n802), .A2(G143), .B1(new_n831), .B2(G159), .ZN(new_n840));
  INV_X1    g0640(.A(new_n789), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  INV_X1    g0642(.A(G150), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n840), .B1(new_n841), .B2(new_n842), .C1(new_n843), .C2(new_n785), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT34), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n302), .B1(new_n793), .B2(G132), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n815), .A2(G68), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n787), .A2(new_n201), .B1(new_n796), .B2(new_n207), .ZN(new_n851));
  NOR4_X1   g0651(.A1(new_n846), .A2(new_n847), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n768), .B1(new_n839), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n768), .A2(new_n765), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n764), .B1(new_n404), .B2(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n853), .B(new_n855), .C1(new_n766), .C2(new_n826), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n829), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G384));
  OAI211_X1 g0658(.A(new_n471), .B(new_n727), .C1(new_n734), .C2(new_n735), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n657), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT99), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n341), .A2(new_n342), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  INV_X1    g0663(.A(new_n699), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n326), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n862), .A2(new_n863), .A3(new_n331), .A4(new_n865), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n305), .A2(new_n307), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT16), .B1(new_n867), .B2(new_n299), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n308), .A2(new_n313), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n325), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n870), .A2(new_n292), .A3(new_n330), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n864), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n862), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n866), .B1(new_n873), .B2(new_n863), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n354), .B2(new_n872), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g0677(.A(KEYINPUT38), .B(new_n874), .C1(new_n354), .C2(new_n872), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n372), .A2(new_n701), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n396), .A2(new_n402), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n391), .A2(KEYINPUT14), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n394), .A2(new_n393), .A3(G169), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(new_n883), .A3(new_n388), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n372), .B(new_n701), .C1(new_n884), .C2(new_n401), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n692), .A2(new_n706), .A3(new_n826), .ZN(new_n887));
  INV_X1    g0687(.A(new_n824), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n879), .A2(new_n889), .B1(new_n335), .B2(new_n699), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n877), .A2(KEYINPUT39), .A3(new_n878), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n351), .A2(new_n352), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n326), .B(new_n864), .C1(new_n892), .C2(new_n335), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n862), .A2(new_n331), .A3(new_n865), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT37), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n866), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n876), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n878), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT39), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n884), .A2(new_n372), .A3(new_n706), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n891), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n890), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n861), .B(new_n905), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n877), .A2(new_n878), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n881), .A2(new_n885), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT40), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n908), .A2(new_n909), .A3(new_n752), .A4(new_n826), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n908), .A2(new_n752), .A3(new_n826), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n878), .B2(new_n898), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n907), .A2(new_n910), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(new_n471), .A3(new_n752), .ZN(new_n914));
  INV_X1    g0714(.A(new_n911), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n909), .B1(new_n899), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n910), .B1(new_n877), .B2(new_n878), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n471), .A2(new_n752), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n914), .A2(G330), .A3(new_n920), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n906), .A2(new_n921), .B1(G1), .B2(new_n757), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n906), .B2(new_n921), .ZN(new_n923));
  INV_X1    g0723(.A(new_n499), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n924), .A2(KEYINPUT35), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(KEYINPUT35), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n925), .A2(G116), .A3(new_n221), .A4(new_n926), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n927), .B(KEYINPUT36), .Z(new_n928));
  NAND3_X1  g0728(.A1(new_n218), .A2(G77), .A3(new_n293), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n207), .A2(G68), .ZN(new_n930));
  AOI211_X1 g0730(.A(new_n277), .B(G13), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n923), .A2(new_n932), .ZN(G367));
  INV_X1    g0733(.A(KEYINPUT44), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n665), .A2(new_n701), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n935), .A2(KEYINPUT100), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(KEYINPUT100), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n521), .A2(new_n556), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n553), .A2(new_n701), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n934), .B1(new_n942), .B2(new_n715), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n936), .A2(new_n937), .B1(new_n939), .B2(new_n940), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(KEYINPUT44), .A3(new_n714), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n942), .A2(new_n715), .A3(KEYINPUT45), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT45), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n944), .B2(new_n714), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n710), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n946), .A2(new_n710), .A3(new_n950), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n711), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n707), .A2(new_n708), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT102), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n958), .A2(new_n712), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n705), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n958), .A2(new_n704), .A3(new_n712), .A4(new_n959), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n755), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(KEYINPUT103), .B1(new_n954), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n754), .B1(new_n961), .B2(new_n962), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT103), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n966), .A2(new_n967), .A3(new_n953), .A4(new_n952), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n754), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n718), .B(KEYINPUT41), .Z(new_n970));
  OAI21_X1  g0770(.A(new_n759), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n944), .A2(new_n712), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n972), .A2(KEYINPUT42), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(KEYINPUT42), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n665), .B1(new_n942), .B2(new_n643), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n973), .A2(new_n974), .B1(new_n701), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n550), .B1(new_n668), .B2(new_n706), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n664), .A2(new_n543), .A3(new_n701), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OR3_X1    g0779(.A1(new_n976), .A2(KEYINPUT43), .A3(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n979), .B(KEYINPUT43), .Z(new_n981));
  NAND2_X1  g0781(.A1(new_n976), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT101), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n976), .A2(KEYINPUT101), .A3(new_n981), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n980), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n710), .A2(new_n944), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n986), .B(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n971), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n773), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n769), .B1(new_n247), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n717), .B2(new_n449), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n801), .A2(new_n843), .B1(new_n792), .B2(new_n842), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n302), .B(new_n993), .C1(G50), .C2(new_n831), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n796), .A2(new_n201), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n787), .A2(new_n202), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n995), .B(new_n996), .C1(G159), .C2(new_n784), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n780), .A2(new_n404), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G143), .B2(new_n789), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n994), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G107), .A2(new_n814), .B1(new_n789), .B2(G311), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n266), .B1(new_n802), .B2(G303), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G283), .A2(new_n831), .B1(new_n793), .B2(G317), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n784), .A2(G294), .B1(new_n815), .B2(G97), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n796), .A2(new_n524), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT46), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1000), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT47), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n764), .B(new_n992), .C1(new_n1009), .C2(new_n768), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n977), .A2(new_n767), .A3(new_n978), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n989), .A2(new_n1012), .ZN(G387));
  NOR2_X1   g0813(.A1(new_n755), .A2(new_n963), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1014), .A2(KEYINPUT106), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(KEYINPUT106), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1015), .A2(new_n718), .A3(new_n964), .A4(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n707), .A2(new_n708), .A3(new_n767), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n776), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n1019), .A2(new_n720), .B1(G107), .B2(new_n214), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n244), .A2(new_n286), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n720), .B(new_n286), .C1(new_n202), .C2(new_n404), .ZN(new_n1022));
  XOR2_X1   g0822(.A(KEYINPUT104), .B(KEYINPUT50), .Z(new_n1023));
  NOR3_X1   g0823(.A1(new_n1023), .A2(G50), .A3(new_n438), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1023), .B1(G50), .B2(new_n438), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n990), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1020), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n761), .B1(new_n1028), .B2(new_n770), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n801), .A2(new_n207), .B1(new_n792), .B2(new_n843), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n302), .B(new_n1030), .C1(G68), .C2(new_n831), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n796), .A2(new_n404), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G97), .B2(new_n815), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G159), .A2(new_n789), .B1(new_n784), .B2(new_n316), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n449), .A2(new_n814), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(G294), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n787), .A2(new_n836), .B1(new_n796), .B2(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n802), .A2(G317), .B1(new_n831), .B2(G303), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n841), .B2(new_n805), .C1(new_n807), .C2(new_n785), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT48), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1038), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n1041), .B2(new_n1040), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT49), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n266), .B1(new_n793), .B2(G326), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n524), .B2(new_n780), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT105), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1036), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1029), .B1(new_n1050), .B2(new_n768), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n963), .A2(new_n760), .B1(new_n1018), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1017), .A2(new_n1052), .ZN(G393));
  AOI22_X1  g0853(.A1(G116), .A2(new_n814), .B1(new_n784), .B2(G303), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1054), .A2(KEYINPUT108), .B1(G294), .B2(new_n831), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(KEYINPUT108), .B2(new_n1054), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT109), .Z(new_n1057));
  AOI22_X1  g0857(.A1(G317), .A2(new_n789), .B1(new_n802), .B2(G311), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT52), .Z(new_n1059));
  OAI21_X1  g0859(.A(new_n302), .B1(new_n792), .B2(new_n805), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n781), .B(new_n1060), .C1(G283), .C2(new_n812), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1057), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n787), .A2(new_n404), .B1(new_n799), .B2(new_n438), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G50), .B2(new_n784), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT107), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G150), .A2(new_n789), .B1(new_n802), .B2(G159), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT51), .Z(new_n1067));
  AOI211_X1 g0867(.A(new_n302), .B(new_n835), .C1(G143), .C2(new_n793), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(new_n202), .C2(new_n796), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1062), .B1(new_n1065), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n768), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n770), .B1(G97), .B2(new_n717), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n251), .A2(new_n773), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n764), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1071), .B(new_n1074), .C1(new_n942), .C2(new_n820), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n954), .B2(new_n759), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT110), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n965), .A2(new_n968), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n719), .B1(new_n954), .B2(new_n964), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1077), .A2(new_n1080), .ZN(G390));
  NAND2_X1  g0881(.A1(new_n891), .A2(new_n901), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n765), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n854), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n761), .B1(new_n1084), .B2(new_n316), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n785), .A2(new_n842), .ZN(new_n1086));
  INV_X1    g0886(.A(G128), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n841), .A2(new_n1087), .B1(new_n780), .B2(new_n207), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1086), .B(new_n1088), .C1(G159), .C2(new_n814), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n796), .A2(new_n843), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1090), .B(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(KEYINPUT54), .B(G143), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n302), .B1(new_n831), .B2(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n802), .A2(G132), .B1(new_n793), .B2(G125), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1089), .A2(new_n1092), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n785), .A2(new_n454), .B1(new_n799), .B2(new_n227), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(KEYINPUT114), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(G77), .A2(new_n814), .B1(new_n789), .B2(G283), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n802), .A2(G116), .B1(new_n793), .B2(G294), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1099), .A2(new_n1100), .A3(new_n849), .A4(new_n1101), .ZN(new_n1102));
  OAI211_X1 g0902(.A(KEYINPUT115), .B(new_n302), .C1(new_n796), .C2(new_n441), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT115), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n797), .B2(new_n266), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1103), .B(new_n1105), .C1(new_n1098), .C2(KEYINPUT114), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1097), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1085), .B1(new_n1107), .B2(new_n768), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT116), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1083), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n826), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n733), .A2(new_n701), .A3(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n908), .B1(new_n1112), .B2(new_n824), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n902), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1082), .A2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n908), .A2(G330), .A3(new_n752), .A4(new_n826), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n825), .A2(new_n465), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n824), .B1(new_n726), .B2(new_n1117), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n1118), .A2(new_n886), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1119), .A2(new_n902), .A3(new_n899), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1115), .A2(new_n1116), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1116), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n891), .A2(new_n901), .B1(new_n1113), .B2(new_n902), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1120), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1126));
  AND4_X1   g0926(.A1(new_n557), .A2(new_n595), .A3(new_n644), .A4(new_n706), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n750), .A2(new_n751), .ZN(new_n1128));
  OAI211_X1 g0928(.A(G330), .B(new_n826), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n886), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n1130), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1116), .A2(new_n1130), .B1(new_n887), .B2(new_n888), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT111), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1130), .A2(new_n1116), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n824), .B2(new_n1112), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(KEYINPUT111), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n753), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n471), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n657), .A2(new_n859), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(KEYINPUT112), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1141), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT112), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1144), .A2(new_n1126), .A3(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1121), .A2(new_n1125), .A3(new_n1145), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n718), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1110), .B1(new_n759), .B2(new_n1126), .C1(new_n1148), .C2(new_n1150), .ZN(G378));
  NOR2_X1   g0951(.A1(new_n266), .A2(G41), .ZN(new_n1152));
  AOI211_X1 g0952(.A(G50), .B(new_n1152), .C1(new_n258), .C2(new_n275), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1152), .B1(new_n836), .B2(new_n792), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n996), .B(new_n1154), .C1(new_n449), .C2(new_n831), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1032), .B1(G116), .B2(new_n789), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n784), .A2(G97), .B1(new_n815), .B2(G58), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n802), .A2(G107), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT117), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .A4(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT58), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1153), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n812), .A2(new_n1094), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT118), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n801), .A2(new_n1087), .B1(new_n799), .B2(new_n842), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G125), .B2(new_n789), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(G150), .A2(new_n814), .B1(new_n784), .B2(G132), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1164), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n815), .A2(G159), .ZN(new_n1170));
  AOI211_X1 g0970(.A(G33), .B(G41), .C1(new_n793), .C2(G124), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1162), .B1(new_n1161), .B2(new_n1160), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n768), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1175), .B(new_n761), .C1(G50), .C2(new_n1084), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n656), .A2(new_n469), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n864), .B1(new_n420), .B2(new_n423), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT55), .Z(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1179), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n656), .A2(new_n469), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  XOR2_X1   g0983(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1180), .A2(new_n1184), .A3(new_n1182), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1176), .B1(new_n1188), .B2(new_n765), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT121), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT120), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1188), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n913), .B2(G330), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1192), .B(G330), .C1(new_n916), .C2(new_n917), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1193), .A2(new_n1195), .A3(new_n905), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n890), .A2(new_n904), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1192), .ZN(new_n1198));
  INV_X1    g0998(.A(G330), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1198), .B1(new_n918), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1197), .B1(new_n1200), .B2(new_n1194), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1190), .B1(new_n1196), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n905), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1200), .A2(new_n1197), .A3(new_n1194), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1203), .A2(KEYINPUT121), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1202), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1189), .B1(new_n1206), .B2(new_n760), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1149), .A2(new_n1142), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT122), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1149), .A2(KEYINPUT122), .A3(new_n1142), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(KEYINPUT57), .B1(new_n1212), .B2(new_n1206), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT57), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1149), .A2(KEYINPUT122), .A3(new_n1142), .ZN(new_n1216));
  AOI21_X1  g1016(.A(KEYINPUT122), .B1(new_n1149), .B2(new_n1142), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1215), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n718), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1207), .B1(new_n1213), .B2(new_n1219), .ZN(G375));
  NAND2_X1  g1020(.A1(new_n886), .A2(new_n765), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n761), .B1(new_n1084), .B2(G68), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n801), .A2(new_n836), .B1(new_n799), .B2(new_n454), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n266), .B(new_n1223), .C1(G303), .C2(new_n793), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n998), .B1(G97), .B2(new_n812), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(G116), .A2(new_n784), .B1(new_n789), .B2(G294), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1224), .A2(new_n1035), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n266), .B1(new_n780), .B2(new_n201), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT123), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n799), .A2(new_n843), .B1(new_n792), .B2(new_n1087), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(G137), .B2(new_n802), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(G132), .A2(new_n789), .B1(new_n784), .B2(new_n1094), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n814), .A2(G50), .B1(new_n812), .B2(G159), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1227), .B1(new_n1229), .B2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1222), .B1(new_n1235), .B2(new_n768), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1138), .A2(new_n760), .B1(new_n1221), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1240), .A2(new_n970), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1238), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(G381));
  INV_X1    g1043(.A(G375), .ZN(new_n1244));
  INV_X1    g1044(.A(G378), .ZN(new_n1245));
  INV_X1    g1045(.A(G390), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(G393), .A2(G396), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1246), .A2(new_n857), .A3(new_n1247), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(new_n1248), .A2(G387), .A3(G381), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1244), .A2(new_n1245), .A3(new_n1249), .ZN(G407));
  NAND2_X1  g1050(.A1(new_n700), .A2(G213), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT124), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1244), .A2(new_n1245), .A3(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(G407), .A2(new_n1253), .A3(G213), .ZN(G409));
  OAI211_X1 g1054(.A(G378), .B(new_n1207), .C1(new_n1213), .C2(new_n1219), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1189), .B1(new_n1256), .B2(new_n760), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1203), .A2(KEYINPUT121), .A3(new_n1204), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT121), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n1258), .A2(new_n1259), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1257), .B1(new_n1260), .B2(new_n970), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1245), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1255), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1240), .A2(KEYINPUT60), .A3(new_n1143), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n718), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1240), .B1(KEYINPUT60), .B2(new_n1143), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n857), .B1(new_n1267), .B2(new_n1238), .ZN(new_n1268));
  OAI211_X1 g1068(.A(G384), .B(new_n1237), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1263), .A2(new_n1271), .A3(new_n1251), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1252), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1268), .A2(KEYINPUT62), .A3(new_n1269), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1263), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT127), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1263), .A2(KEYINPUT127), .A3(new_n1276), .A4(new_n1275), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1274), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1263), .A2(new_n1275), .ZN(new_n1282));
  INV_X1    g1082(.A(G2897), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1251), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1271), .A2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1270), .B1(new_n1283), .B2(new_n1275), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT61), .B1(new_n1282), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1281), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n989), .A2(new_n1012), .A3(G390), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(G390), .B1(new_n989), .B2(new_n1012), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n822), .B1(new_n1017), .B2(new_n1052), .ZN(new_n1293));
  OAI22_X1  g1093(.A1(new_n1291), .A2(new_n1292), .B1(new_n1247), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1292), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1247), .A2(new_n1293), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1295), .A2(new_n1296), .A3(new_n1290), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1294), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1289), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT125), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT63), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1270), .A2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1263), .A2(new_n1275), .A3(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT61), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1294), .A2(new_n1297), .A3(new_n1304), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1251), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(new_n1255), .B2(new_n1262), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1303), .B(new_n1305), .C1(new_n1306), .C2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT63), .B1(new_n1308), .B2(new_n1271), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1300), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1294), .A2(new_n1297), .A3(new_n1304), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1263), .A2(new_n1251), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1312), .B1(new_n1313), .B2(new_n1287), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1272), .A2(new_n1301), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1314), .A2(new_n1315), .A3(KEYINPUT125), .A4(new_n1303), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1311), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1299), .A2(new_n1317), .ZN(G405));
  NAND2_X1  g1118(.A1(G375), .A2(new_n1245), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1255), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(new_n1320), .B(new_n1270), .ZN(new_n1321));
  XOR2_X1   g1121(.A(new_n1321), .B(new_n1298), .Z(G402));
endmodule


