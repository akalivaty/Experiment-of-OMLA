//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n972, new_n973,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1023, new_n1024;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n202));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n205), .A2(KEYINPUT26), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(KEYINPUT26), .ZN(new_n207));
  AOI22_X1  g006(.A1(new_n206), .A2(new_n207), .B1(G169gat), .B2(G176gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT27), .B(G183gat), .ZN(new_n209));
  INV_X1    g008(.A(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT28), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n209), .A2(KEYINPUT28), .A3(new_n210), .ZN(new_n214));
  AOI211_X1 g013(.A(new_n204), .B(new_n208), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n203), .A2(KEYINPUT24), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n203), .A2(KEYINPUT24), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(G169gat), .B2(G176gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT66), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n205), .A2(KEYINPUT23), .ZN(new_n227));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n222), .A2(new_n226), .A3(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n219), .B1(new_n216), .B2(new_n217), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT25), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n235), .B1(new_n228), .B2(KEYINPUT67), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n236), .B(new_n227), .C1(KEYINPUT67), .C2(new_n228), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n231), .A2(new_n233), .B1(new_n238), .B2(new_n226), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n215), .B1(new_n239), .B2(KEYINPUT68), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n224), .B(KEYINPUT66), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(new_n229), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n232), .B1(new_n243), .B2(new_n222), .ZN(new_n244));
  NOR3_X1   g043(.A1(new_n242), .A2(new_n234), .A3(new_n237), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n241), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT29), .B1(new_n240), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G226gat), .A2(G233gat), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n202), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n231), .A2(new_n233), .ZN(new_n251));
  INV_X1    g050(.A(new_n245), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT68), .ZN(new_n253));
  INV_X1    g052(.A(new_n215), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n246), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT29), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n257), .A2(KEYINPUT75), .A3(new_n248), .ZN(new_n258));
  OR2_X1    g057(.A1(new_n239), .A2(new_n215), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(new_n249), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n250), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G197gat), .B(G204gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT73), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT22), .ZN(new_n264));
  INV_X1    g063(.A(G211gat), .ZN(new_n265));
  INV_X1    g064(.A(G218gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G211gat), .B(G218gat), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n263), .A2(new_n269), .A3(new_n267), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT74), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT74), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n271), .A2(new_n275), .A3(new_n272), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n273), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n259), .A2(new_n256), .A3(new_n248), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n240), .A2(new_n249), .A3(new_n246), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G8gat), .B(G36gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(G64gat), .B(G92gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n279), .A2(KEYINPUT30), .A3(new_n284), .A4(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n249), .B1(new_n255), .B2(new_n256), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n290), .A2(KEYINPUT75), .B1(new_n249), .B2(new_n259), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n277), .B1(new_n291), .B2(new_n250), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n287), .B1(new_n292), .B2(new_n283), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(G1gat), .B(G29gat), .Z(new_n295));
  XNOR2_X1  g094(.A(G57gat), .B(G85gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n298));
  XOR2_X1   g097(.A(new_n297), .B(new_n298), .Z(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G225gat), .A2(G233gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303));
  INV_X1    g102(.A(G155gat), .ZN(new_n304));
  INV_X1    g103(.A(G162gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n303), .B1(new_n306), .B2(KEYINPUT2), .ZN(new_n307));
  INV_X1    g106(.A(G141gat), .ZN(new_n308));
  INV_X1    g107(.A(G148gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G141gat), .A2(G148gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(KEYINPUT77), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT77), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n314), .B1(new_n310), .B2(new_n311), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n307), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n306), .A2(new_n303), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT2), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n310), .A2(new_n318), .A3(new_n311), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G113gat), .B(G120gat), .ZN(new_n322));
  OR2_X1    g121(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G127gat), .B(G134gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n325), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n327), .B1(new_n322), .B2(new_n323), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n321), .A2(new_n329), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n316), .A2(new_n320), .B1(new_n328), .B2(new_n326), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n302), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT5), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n312), .B(KEYINPUT77), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n334), .A2(new_n307), .B1(new_n319), .B2(new_n317), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT78), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT3), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT78), .B1(new_n321), .B2(KEYINPUT3), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n321), .A2(KEYINPUT3), .B1(new_n328), .B2(new_n326), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n302), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n321), .A2(KEYINPUT4), .A3(new_n329), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n329), .A2(KEYINPUT70), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT70), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n326), .A2(new_n328), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n335), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n343), .B1(new_n347), .B2(KEYINPUT4), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n333), .B1(new_n342), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n336), .B1(new_n335), .B2(new_n337), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n321), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n341), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT4), .B1(new_n321), .B2(new_n329), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(new_n347), .B2(KEYINPUT4), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n302), .A2(KEYINPUT5), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n353), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n300), .B1(new_n350), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT6), .ZN(new_n360));
  OR2_X1    g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n333), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n353), .A2(new_n301), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n362), .B1(new_n363), .B2(new_n348), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(new_n299), .A3(new_n357), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n359), .A2(new_n365), .A3(new_n360), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  AOI211_X1 g166(.A(new_n283), .B(new_n287), .C1(new_n261), .C2(new_n278), .ZN(new_n368));
  NOR3_X1   g167(.A1(new_n368), .A2(KEYINPUT76), .A3(KEYINPUT30), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT76), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n279), .A2(new_n284), .A3(new_n288), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT30), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n294), .B(new_n367), .C1(new_n369), .C2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT29), .B1(new_n271), .B2(new_n272), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n321), .B1(new_n375), .B2(KEYINPUT3), .ZN(new_n376));
  INV_X1    g175(.A(G228gat), .ZN(new_n377));
  INV_X1    g176(.A(G233gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT29), .B1(new_n338), .B2(new_n339), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n376), .B(new_n379), .C1(new_n277), .C2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n256), .B1(new_n351), .B2(new_n352), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n280), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n379), .B1(new_n384), .B2(new_n376), .ZN(new_n385));
  OAI21_X1  g184(.A(G22gat), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n376), .ZN(new_n387));
  INV_X1    g186(.A(new_n379), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(G22gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n390), .A3(new_n381), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G78gat), .B(G106gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT31), .B(G50gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n397));
  INV_X1    g196(.A(new_n272), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n269), .B1(new_n263), .B2(new_n267), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n256), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n337), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n388), .B1(new_n401), .B2(new_n321), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n383), .A2(new_n274), .A3(new_n276), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n387), .A2(new_n388), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n397), .B1(new_n404), .B2(new_n390), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n392), .A2(new_n396), .A3(new_n405), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n386), .B(new_n391), .C1(new_n397), .C2(new_n395), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n344), .A2(new_n346), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n255), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(G227gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n412), .A2(new_n378), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n240), .A2(new_n409), .A3(new_n246), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n411), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT32), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT33), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  XOR2_X1   g217(.A(G15gat), .B(G43gat), .Z(new_n419));
  XNOR2_X1  g218(.A(G71gat), .B(G99gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT71), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n416), .B1(new_n421), .B2(KEYINPUT33), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n415), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n423), .B1(new_n415), .B2(new_n424), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n422), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n413), .B1(new_n411), .B2(new_n414), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT34), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI211_X1 g229(.A(KEYINPUT34), .B(new_n413), .C1(new_n411), .C2(new_n414), .ZN(new_n431));
  OR2_X1    g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n415), .A2(new_n424), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT71), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n415), .A2(new_n423), .A3(new_n424), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n430), .A2(new_n431), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n422), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n408), .A2(new_n433), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT35), .B1(new_n374), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT83), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT83), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n443), .B(KEYINPUT35), .C1(new_n374), .C2(new_n440), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n433), .A2(new_n439), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT82), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT82), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n433), .A2(new_n439), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n366), .A2(KEYINPUT81), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n450), .A2(new_n361), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT81), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n359), .A2(new_n365), .A3(new_n452), .A4(new_n360), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT35), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n289), .A2(new_n293), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT76), .B1(new_n368), .B2(KEYINPUT30), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n371), .A2(new_n370), .A3(new_n372), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n449), .A2(new_n454), .A3(new_n458), .A4(new_n408), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n442), .A2(new_n444), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT72), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT36), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n445), .A2(KEYINPUT72), .A3(KEYINPUT36), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n406), .A2(new_n407), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n294), .B1(new_n369), .B2(new_n373), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n301), .B1(new_n353), .B2(new_n355), .ZN(new_n469));
  OR2_X1    g268(.A1(new_n330), .A2(new_n331), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT39), .B1(new_n470), .B2(new_n302), .ZN(new_n471));
  OR2_X1    g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT39), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n472), .A2(new_n299), .A3(new_n474), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n475), .A2(KEYINPUT40), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(KEYINPUT40), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(new_n359), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n468), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT37), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n279), .A2(new_n481), .A3(new_n284), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n287), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n279), .B2(new_n284), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT38), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND4_X1   g284(.A1(new_n361), .A2(new_n450), .A3(new_n371), .A4(new_n453), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n281), .A2(new_n280), .A3(new_n282), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(new_n261), .B2(new_n278), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT38), .B1(new_n488), .B2(KEYINPUT37), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n489), .A2(new_n287), .A3(new_n482), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n485), .A2(new_n486), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n467), .B1(new_n480), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n374), .A2(new_n408), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n466), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n460), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G15gat), .B(G22gat), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n496), .A2(G1gat), .ZN(new_n497));
  INV_X1    g296(.A(G8gat), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT85), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT16), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n499), .B1(new_n500), .B2(G1gat), .ZN(new_n501));
  INV_X1    g300(.A(G1gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n502), .A2(KEYINPUT85), .A3(KEYINPUT16), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n496), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n497), .A2(new_n498), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT87), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT86), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n497), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n504), .A2(new_n508), .ZN(new_n511));
  OAI21_X1  g310(.A(G8gat), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(G71gat), .A2(G78gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT9), .ZN(new_n515));
  NAND2_X1  g314(.A1(G71gat), .A2(G78gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(G57gat), .ZN(new_n518));
  INV_X1    g317(.A(G64gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G57gat), .A2(G64gat), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n520), .A2(KEYINPUT91), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT91), .B1(new_n520), .B2(new_n521), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n517), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n516), .B1(new_n514), .B2(KEYINPUT90), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n520), .A2(new_n521), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n527));
  OAI221_X1 g326(.A(new_n525), .B1(KEYINPUT90), .B2(new_n516), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT93), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n513), .B1(KEYINPUT21), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT21), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G231gat), .A2(G233gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n534), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n533), .B(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n536), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G127gat), .B(G155gat), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n542), .B(KEYINPUT20), .Z(new_n543));
  NAND3_X1  g342(.A1(new_n537), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n543), .B1(new_n537), .B2(new_n541), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n531), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n537), .A2(new_n541), .ZN(new_n548));
  INV_X1    g347(.A(new_n543), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n531), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(new_n551), .A3(new_n544), .ZN(new_n552));
  XOR2_X1   g351(.A(G183gat), .B(G211gat), .Z(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n547), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n554), .B1(new_n547), .B2(new_n552), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G134gat), .B(G162gat), .Z(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT84), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g362(.A(KEYINPUT84), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR3_X1   g364(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(G29gat), .ZN(new_n569));
  INV_X1    g368(.A(G36gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n568), .A2(KEYINPUT15), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT15), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n566), .B1(new_n563), .B2(new_n564), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n574), .B1(new_n575), .B2(new_n571), .ZN(new_n576));
  XOR2_X1   g375(.A(G43gat), .B(G50gat), .Z(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n573), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n568), .A2(KEYINPUT15), .A3(new_n572), .A4(new_n577), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(KEYINPUT17), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT88), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n579), .A2(KEYINPUT88), .A3(KEYINPUT17), .A4(new_n580), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OR2_X1    g384(.A1(KEYINPUT95), .A2(G92gat), .ZN(new_n586));
  INV_X1    g385(.A(G85gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(KEYINPUT95), .A2(G92gat), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT7), .ZN(new_n590));
  NAND2_X1  g389(.A1(G85gat), .A2(G92gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(G99gat), .A2(G106gat), .ZN(new_n592));
  AOI22_X1  g391(.A1(new_n590), .A2(new_n591), .B1(new_n592), .B2(KEYINPUT8), .ZN(new_n593));
  NAND3_X1  g392(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n589), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G99gat), .B(G106gat), .Z(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n596), .A2(new_n589), .A3(new_n593), .A4(new_n594), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n579), .A2(new_n580), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT17), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n585), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n579), .A2(new_n580), .ZN(new_n606));
  OAI211_X1 g405(.A(KEYINPUT96), .B(new_n605), .C1(new_n606), .C2(new_n600), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT96), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n600), .B1(new_n579), .B2(new_n580), .ZN(new_n609));
  INV_X1    g408(.A(new_n605), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G190gat), .B(G218gat), .Z(new_n613));
  NAND3_X1  g412(.A1(new_n604), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n613), .B1(new_n604), .B2(new_n612), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT97), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g416(.A1(new_n583), .A2(new_n584), .B1(new_n602), .B2(new_n601), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n618), .A2(new_n600), .B1(new_n607), .B2(new_n611), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n619), .A2(KEYINPUT97), .A3(new_n613), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n560), .B1(new_n617), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(KEYINPUT97), .B1(new_n619), .B2(new_n613), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n615), .A2(new_n616), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n622), .A2(new_n623), .A3(new_n614), .A4(new_n559), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT94), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n621), .A2(new_n627), .A3(new_n624), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n558), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G113gat), .B(G141gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT11), .ZN(new_n633));
  INV_X1    g432(.A(G169gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(G197gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  INV_X1    g437(.A(new_n513), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n618), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G229gat), .A2(G233gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n513), .A2(new_n601), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n640), .A2(KEYINPUT18), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n641), .B(KEYINPUT13), .Z(new_n644));
  AOI22_X1  g443(.A1(new_n507), .A2(new_n512), .B1(new_n580), .B2(new_n579), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n606), .A2(new_n512), .A3(new_n507), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT89), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n642), .A2(KEYINPUT89), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n644), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n645), .B1(new_n618), .B2(new_n639), .ZN(new_n652));
  AOI21_X1  g451(.A(KEYINPUT18), .B1(new_n652), .B2(new_n641), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n638), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT18), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n642), .ZN(new_n656));
  INV_X1    g455(.A(new_n641), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n638), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n658), .A2(new_n643), .A3(new_n650), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(G120gat), .B(G148gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT100), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n598), .A2(new_n599), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n530), .A2(KEYINPUT10), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT98), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n595), .A2(new_n668), .A3(new_n596), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n596), .B1(new_n595), .B2(new_n668), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n528), .B(new_n524), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n666), .A2(new_n529), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT10), .ZN(new_n675));
  AOI21_X1  g474(.A(KEYINPUT99), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT99), .ZN(new_n677));
  AOI211_X1 g476(.A(new_n677), .B(KEYINPUT10), .C1(new_n672), .C2(new_n673), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n667), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(G230gat), .A2(G233gat), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n680), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n672), .A2(new_n673), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n665), .B1(new_n685), .B2(KEYINPUT101), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT101), .ZN(new_n687));
  INV_X1    g486(.A(new_n665), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n684), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n631), .A2(new_n661), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n495), .A2(KEYINPUT102), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT102), .B1(new_n495), .B2(new_n692), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n367), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(new_n502), .ZN(G1324gat));
  INV_X1    g496(.A(new_n695), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT16), .B(G8gat), .Z(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(new_n468), .A3(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n698), .A2(new_n468), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n704), .A2(KEYINPUT103), .A3(G8gat), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT103), .B1(new_n704), .B2(G8gat), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n702), .B(new_n703), .C1(new_n705), .C2(new_n706), .ZN(G1325gat));
  INV_X1    g506(.A(new_n449), .ZN(new_n708));
  OR3_X1    g507(.A1(new_n695), .A2(G15gat), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(G15gat), .B1(new_n695), .B2(new_n466), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(G1326gat));
  OR3_X1    g510(.A1(new_n695), .A2(KEYINPUT104), .A3(new_n408), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT104), .B1(new_n695), .B2(new_n408), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT43), .B(G22gat), .Z(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1327gat));
  NAND2_X1  g515(.A1(new_n629), .A2(new_n630), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n717), .B1(new_n460), .B2(new_n494), .ZN(new_n718));
  INV_X1    g517(.A(new_n690), .ZN(new_n719));
  INV_X1    g518(.A(new_n661), .ZN(new_n720));
  INV_X1    g519(.A(new_n557), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n555), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n367), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(new_n569), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT45), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n444), .A2(new_n459), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n467), .A2(new_n445), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n730), .A2(new_n458), .A3(new_n367), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n443), .B1(new_n731), .B2(KEYINPUT35), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n485), .A2(new_n486), .A3(new_n490), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n456), .A2(new_n457), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n478), .B1(new_n735), .B2(new_n294), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n408), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n493), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n465), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n728), .B1(new_n733), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n460), .A2(new_n494), .A3(KEYINPUT105), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n717), .A2(KEYINPUT44), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n717), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n733), .B2(new_n739), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(KEYINPUT44), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n747), .A2(new_n723), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n748), .A2(new_n725), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n727), .B1(new_n749), .B2(new_n569), .ZN(G1328gat));
  NAND3_X1  g549(.A1(new_n724), .A2(new_n570), .A3(new_n468), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT106), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT46), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n748), .A2(new_n468), .ZN(new_n756));
  OAI22_X1  g555(.A1(new_n754), .A2(new_n755), .B1(new_n570), .B2(new_n756), .ZN(G1329gat));
  AOI21_X1  g556(.A(G43gat), .B1(new_n724), .B2(new_n449), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n465), .A2(G43gat), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n758), .B1(new_n748), .B2(new_n759), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g560(.A(G50gat), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n762), .B1(new_n748), .B2(new_n467), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT48), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n408), .A2(G50gat), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT107), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n724), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  OR3_X1    g567(.A1(new_n763), .A2(new_n764), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n764), .B1(new_n763), .B2(new_n768), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1331gat));
  AND2_X1   g570(.A1(new_n740), .A2(new_n741), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n621), .A2(new_n627), .A3(new_n624), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n627), .B1(new_n621), .B2(new_n624), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n722), .B(new_n720), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(new_n690), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n777), .A2(new_n367), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(new_n518), .ZN(G1332gat));
  INV_X1    g578(.A(new_n777), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n458), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n784));
  AND2_X1   g583(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(new_n784), .B2(new_n783), .ZN(G1333gat));
  NAND3_X1  g586(.A1(new_n780), .A2(G71gat), .A3(new_n465), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n777), .A2(new_n708), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(G71gat), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g589(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n790), .B(new_n791), .ZN(G1334gat));
  NAND2_X1  g591(.A1(new_n780), .A2(new_n467), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g593(.A1(new_n722), .A2(new_n661), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n744), .B(new_n795), .C1(new_n733), .C2(new_n739), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n718), .A2(KEYINPUT51), .A3(new_n795), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(new_n690), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(new_n587), .A3(new_n725), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n795), .A2(new_n719), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n747), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(G85gat), .B1(new_n806), .B2(new_n367), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n803), .A2(new_n807), .ZN(G1336gat));
  NAND2_X1  g607(.A1(new_n586), .A2(new_n588), .ZN(new_n809));
  INV_X1    g608(.A(new_n782), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n809), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n810), .A2(G92gat), .A3(new_n690), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT110), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n811), .B(new_n812), .C1(new_n801), .C2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n814), .B1(new_n798), .B2(new_n799), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n804), .B1(new_n743), .B2(new_n746), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n468), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n816), .B1(new_n818), .B2(new_n809), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n819), .A2(new_n820), .A3(new_n812), .ZN(new_n821));
  AOI211_X1 g620(.A(new_n458), .B(new_n804), .C1(new_n743), .C2(new_n746), .ZN(new_n822));
  INV_X1    g621(.A(new_n809), .ZN(new_n823));
  OAI22_X1  g622(.A1(new_n822), .A2(new_n823), .B1(new_n801), .B2(new_n814), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT111), .B1(new_n824), .B2(KEYINPUT52), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n815), .B1(new_n821), .B2(new_n825), .ZN(G1337gat));
  INV_X1    g625(.A(G99gat), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n802), .A2(new_n827), .A3(new_n449), .ZN(new_n828));
  OAI21_X1  g627(.A(G99gat), .B1(new_n806), .B2(new_n466), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(G1338gat));
  INV_X1    g629(.A(KEYINPUT112), .ZN(new_n831));
  AOI211_X1 g630(.A(new_n408), .B(new_n804), .C1(new_n743), .C2(new_n746), .ZN(new_n832));
  INV_X1    g631(.A(G106gat), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n719), .A2(new_n467), .A3(new_n833), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT113), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT114), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT115), .B1(new_n800), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840));
  AOI211_X1 g639(.A(new_n840), .B(new_n837), .C1(new_n798), .C2(new_n799), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g641(.A(KEYINPUT112), .B(G106gat), .C1(new_n806), .C2(new_n408), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n834), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(KEYINPUT53), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n833), .B1(new_n817), .B2(new_n467), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n796), .A2(new_n797), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT51), .B1(new_n718), .B2(new_n795), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n836), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n846), .B1(new_n847), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT53), .B1(new_n800), .B2(new_n836), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n854), .B(KEYINPUT116), .C1(new_n832), .C2(new_n833), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n845), .A2(new_n856), .ZN(G1339gat));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n858));
  OAI21_X1  g657(.A(KEYINPUT117), .B1(new_n775), .B2(new_n719), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n631), .A2(new_n860), .A3(new_n720), .A4(new_n690), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n648), .A2(new_n649), .ZN(new_n864));
  OAI22_X1  g663(.A1(new_n864), .A2(new_n644), .B1(new_n641), .B2(new_n652), .ZN(new_n865));
  INV_X1    g664(.A(new_n637), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n867), .A2(new_n660), .ZN(new_n868));
  INV_X1    g667(.A(new_n673), .ZN(new_n869));
  INV_X1    g668(.A(new_n671), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n529), .B1(new_n870), .B2(new_n669), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n675), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n677), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n674), .A2(KEYINPUT99), .A3(new_n675), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n682), .B1(new_n875), .B2(new_n667), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n688), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n875), .A2(new_n667), .A3(new_n682), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n681), .A2(new_n879), .A3(KEYINPUT54), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT55), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n878), .A2(new_n880), .A3(KEYINPUT55), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n685), .A2(new_n688), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n868), .A2(new_n883), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n717), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n661), .A2(new_n883), .A3(new_n884), .A4(new_n885), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n686), .A2(new_n867), .A3(new_n660), .A4(new_n689), .ZN(new_n889));
  AOI22_X1  g688(.A1(new_n888), .A2(new_n889), .B1(new_n629), .B2(new_n630), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n558), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n862), .A2(new_n863), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n863), .B1(new_n862), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n782), .A2(new_n367), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(new_n730), .A3(new_n895), .ZN(new_n896));
  XOR2_X1   g695(.A(new_n896), .B(KEYINPUT119), .Z(new_n897));
  INV_X1    g696(.A(G113gat), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n661), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n894), .A2(new_n895), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n408), .A3(new_n449), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(new_n720), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n903), .A2(new_n898), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n858), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  OAI221_X1 g704(.A(KEYINPUT120), .B1(new_n903), .B2(new_n898), .C1(new_n897), .C2(new_n899), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1340gat));
  OAI21_X1  g706(.A(G120gat), .B1(new_n902), .B2(new_n690), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n690), .A2(G120gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n897), .B2(new_n909), .ZN(G1341gat));
  OAI21_X1  g709(.A(G127gat), .B1(new_n902), .B2(new_n558), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n558), .A2(G127gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n896), .B2(new_n912), .ZN(G1342gat));
  NAND2_X1  g712(.A1(new_n862), .A2(new_n891), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT118), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n862), .A2(new_n891), .A3(new_n863), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR4_X1   g716(.A1(new_n917), .A2(new_n367), .A3(new_n468), .A4(new_n717), .ZN(new_n918));
  INV_X1    g717(.A(G134gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n918), .A2(new_n919), .A3(new_n730), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT56), .Z(new_n921));
  OAI21_X1  g720(.A(G134gat), .B1(new_n902), .B2(new_n717), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1343gat));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT58), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n888), .A2(KEYINPUT121), .A3(new_n889), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT121), .B1(new_n888), .B2(new_n889), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n717), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n887), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n722), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n862), .ZN(new_n931));
  OAI211_X1 g730(.A(KEYINPUT57), .B(new_n467), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n892), .A2(new_n893), .A3(new_n408), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(KEYINPUT57), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n895), .A2(new_n466), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n934), .A2(new_n661), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(G141gat), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n465), .A2(new_n408), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n720), .A2(G141gat), .ZN(new_n940));
  AND4_X1   g739(.A1(new_n894), .A2(new_n895), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n925), .B1(new_n938), .B2(new_n942), .ZN(new_n943));
  AOI211_X1 g742(.A(KEYINPUT58), .B(new_n941), .C1(new_n937), .C2(G141gat), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n924), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n915), .A2(new_n467), .A3(new_n916), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT57), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n935), .B1(new_n948), .B2(new_n932), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n308), .B1(new_n949), .B2(new_n661), .ZN(new_n950));
  OAI21_X1  g749(.A(KEYINPUT58), .B1(new_n950), .B2(new_n941), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n938), .A2(new_n925), .A3(new_n942), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n951), .A2(new_n952), .A3(KEYINPUT122), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n945), .A2(new_n953), .ZN(G1344gat));
  AND2_X1   g753(.A1(new_n901), .A2(new_n939), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n955), .A2(new_n309), .A3(new_n719), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT123), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT59), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n775), .A2(new_n719), .ZN(new_n961));
  OR2_X1    g760(.A1(new_n930), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n408), .A2(KEYINPUT57), .ZN(new_n963));
  AOI22_X1  g762(.A1(new_n946), .A2(KEYINPUT57), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n964), .A2(new_n719), .A3(new_n936), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n960), .B1(new_n965), .B2(G148gat), .ZN(new_n966));
  AOI211_X1 g765(.A(KEYINPUT59), .B(new_n309), .C1(new_n949), .C2(new_n719), .ZN(new_n967));
  OAI22_X1  g766(.A1(new_n958), .A2(new_n959), .B1(new_n966), .B2(new_n967), .ZN(G1345gat));
  NAND3_X1  g767(.A1(new_n955), .A2(new_n304), .A3(new_n722), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n949), .A2(new_n722), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n969), .B1(new_n970), .B2(new_n304), .ZN(G1346gat));
  NAND3_X1  g770(.A1(new_n918), .A2(new_n305), .A3(new_n939), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n949), .A2(new_n744), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n972), .B1(new_n973), .B2(new_n305), .ZN(G1347gat));
  NAND2_X1  g773(.A1(new_n468), .A2(new_n367), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n708), .A2(new_n975), .A3(new_n467), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n894), .A2(new_n976), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n977), .A2(new_n634), .A3(new_n720), .ZN(new_n978));
  NOR3_X1   g777(.A1(new_n917), .A2(new_n725), .A3(new_n810), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(new_n730), .ZN(new_n980));
  XOR2_X1   g779(.A(new_n980), .B(KEYINPUT124), .Z(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(new_n661), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n978), .B1(new_n982), .B2(new_n634), .ZN(G1348gat));
  INV_X1    g782(.A(G176gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n981), .A2(new_n984), .A3(new_n719), .ZN(new_n985));
  OAI21_X1  g784(.A(G176gat), .B1(new_n977), .B2(new_n690), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(G1349gat));
  OAI21_X1  g786(.A(G183gat), .B1(new_n977), .B2(new_n558), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n722), .A2(new_n209), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n988), .B1(new_n980), .B2(new_n989), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n990), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g790(.A1(new_n894), .A2(new_n744), .A3(new_n976), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n992), .A2(G190gat), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT61), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT125), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n992), .A2(new_n994), .A3(G190gat), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n998), .B1(new_n996), .B2(new_n997), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n981), .A2(new_n210), .A3(new_n744), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(G1351gat));
  NAND2_X1  g800(.A1(new_n979), .A2(new_n939), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n661), .A2(new_n636), .ZN(new_n1003));
  OAI21_X1  g802(.A(KEYINPUT126), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  OR3_X1    g803(.A1(new_n1002), .A2(KEYINPUT126), .A3(new_n1003), .ZN(new_n1005));
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n1006));
  NOR2_X1   g805(.A1(new_n465), .A2(new_n975), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n964), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1006), .B1(new_n1008), .B2(new_n720), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1009), .A2(G197gat), .ZN(new_n1010));
  NOR3_X1   g809(.A1(new_n1008), .A2(new_n1006), .A3(new_n720), .ZN(new_n1011));
  OAI211_X1 g810(.A(new_n1004), .B(new_n1005), .C1(new_n1010), .C2(new_n1011), .ZN(G1352gat));
  NOR3_X1   g811(.A1(new_n1002), .A2(G204gat), .A3(new_n690), .ZN(new_n1013));
  XNOR2_X1  g812(.A(new_n1013), .B(KEYINPUT62), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n964), .A2(new_n719), .A3(new_n1007), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1015), .A2(G204gat), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1014), .A2(new_n1016), .ZN(G1353gat));
  NAND3_X1  g816(.A1(new_n964), .A2(new_n722), .A3(new_n1007), .ZN(new_n1018));
  AND3_X1   g817(.A1(new_n1018), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1019));
  AOI21_X1  g818(.A(KEYINPUT63), .B1(new_n1018), .B2(G211gat), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n722), .A2(new_n265), .ZN(new_n1021));
  OAI22_X1  g820(.A1(new_n1019), .A2(new_n1020), .B1(new_n1002), .B2(new_n1021), .ZN(G1354gat));
  OAI21_X1  g821(.A(G218gat), .B1(new_n1008), .B2(new_n717), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n744), .A2(new_n266), .ZN(new_n1024));
  OAI21_X1  g823(.A(new_n1023), .B1(new_n1002), .B2(new_n1024), .ZN(G1355gat));
endmodule


