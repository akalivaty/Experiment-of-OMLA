//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 0 0 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n587, new_n588,
    new_n589, new_n590, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n631, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT65), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT66), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(new_n452), .B2(G2106), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT3), .B1(new_n461), .B2(KEYINPUT69), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(new_n471), .A3(G2104), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n468), .A2(G137), .A3(new_n469), .A4(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(G125), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n468), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n463), .B(new_n473), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  AOI211_X1 g055(.A(KEYINPUT68), .B(new_n468), .C1(new_n476), .C2(new_n477), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n480), .A2(new_n481), .ZN(G160));
  NAND2_X1  g057(.A1(new_n469), .A2(new_n472), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT70), .ZN(new_n486));
  OAI221_X1 g061(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n468), .C2(G112), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n483), .A2(new_n468), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G124), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n492), .B(KEYINPUT71), .ZN(G162));
  NAND4_X1  g068(.A1(new_n468), .A2(G138), .A3(new_n469), .A4(new_n472), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT73), .ZN(new_n496));
  OR2_X1    g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(new_n475), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n497), .A2(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n502), .B1(new_n466), .B2(new_n467), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n495), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n469), .A2(new_n472), .A3(G126), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT72), .A2(G114), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT72), .A2(G114), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(G2104), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G2105), .B1(G102), .B2(new_n462), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT74), .A2(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n517), .A2(KEYINPUT74), .A3(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G62), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n514), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G651), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT75), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g099(.A(KEYINPUT75), .B1(new_n521), .B2(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT6), .B(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n526), .A2(new_n516), .A3(new_n518), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G50), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n527), .A2(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR3_X1   g106(.A1(new_n524), .A2(new_n525), .A3(new_n531), .ZN(G166));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT76), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT76), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n535), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n534), .A2(KEYINPUT7), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(KEYINPUT7), .B1(new_n534), .B2(new_n536), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n526), .A2(G51), .A3(G543), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n516), .A2(new_n518), .A3(G63), .A4(G651), .ZN(new_n541));
  INV_X1    g116(.A(G89), .ZN(new_n542));
  OAI211_X1 g117(.A(new_n540), .B(new_n541), .C1(new_n527), .C2(new_n542), .ZN(new_n543));
  OAI21_X1  g118(.A(KEYINPUT77), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n540), .A2(new_n541), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n526), .A2(new_n516), .A3(new_n518), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G89), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n537), .A2(new_n538), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT77), .ZN(new_n549));
  NAND4_X1  g124(.A1(new_n545), .A2(new_n547), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n544), .A2(new_n550), .ZN(G168));
  NAND2_X1  g126(.A1(G77), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G64), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n519), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G651), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(KEYINPUT78), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(KEYINPUT78), .ZN(new_n557));
  AND2_X1   g132(.A1(new_n526), .A2(G543), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n546), .A2(G90), .B1(new_n558), .B2(G52), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(G301));
  INV_X1    g135(.A(G301), .ZN(G171));
  INV_X1    g136(.A(G651), .ZN(new_n562));
  AND2_X1   g137(.A1(new_n516), .A2(new_n518), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G56), .ZN(new_n564));
  NAND2_X1  g139(.A1(G68), .A2(G543), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(G81), .ZN(new_n567));
  INV_X1    g142(.A(G43), .ZN(new_n568));
  OAI22_X1  g143(.A1(new_n527), .A2(new_n567), .B1(new_n529), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G860), .ZN(G153));
  AND3_X1   g146(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G36), .ZN(G176));
  NAND2_X1  g148(.A1(G1), .A2(G3), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT8), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n572), .A2(new_n575), .ZN(G188));
  INV_X1    g151(.A(G53), .ZN(new_n577));
  OR3_X1    g152(.A1(new_n529), .A2(KEYINPUT9), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(KEYINPUT9), .B1(new_n529), .B2(new_n577), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n563), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G91), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n527), .A2(new_n582), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n583), .A2(KEYINPUT79), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n583), .A2(KEYINPUT79), .ZN(new_n585));
  OAI221_X1 g160(.A(new_n580), .B1(new_n562), .B2(new_n581), .C1(new_n584), .C2(new_n585), .ZN(G299));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n587));
  NAND2_X1  g162(.A1(G168), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n544), .A2(KEYINPUT80), .A3(new_n550), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G286));
  OR3_X1    g166(.A1(new_n524), .A2(new_n525), .A3(new_n531), .ZN(G303));
  OAI21_X1  g167(.A(G651), .B1(new_n563), .B2(G74), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n594), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n546), .A2(G87), .B1(new_n558), .B2(G49), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G288));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G61), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n519), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(new_n558), .B2(G48), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n546), .A2(G86), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G305));
  AOI22_X1  g179(.A1(new_n563), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n605), .A2(new_n562), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n526), .A2(G47), .A3(G543), .ZN(new_n607));
  INV_X1    g182(.A(G85), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n527), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(KEYINPUT82), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT82), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n563), .A2(G85), .A3(new_n526), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(new_n607), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n610), .B2(new_n613), .ZN(G290));
  NAND2_X1  g189(.A1(G301), .A2(G868), .ZN(new_n615));
  INV_X1    g190(.A(G92), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n527), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT10), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n519), .B2(new_n620), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n621), .A2(G651), .B1(new_n558), .B2(G54), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n615), .B1(new_n624), .B2(G868), .ZN(G284));
  OAI21_X1  g200(.A(new_n615), .B1(new_n624), .B2(G868), .ZN(G321));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(G299), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(new_n590), .B2(new_n627), .ZN(G297));
  OAI21_X1  g204(.A(new_n628), .B1(new_n590), .B2(new_n627), .ZN(G280));
  XOR2_X1   g205(.A(KEYINPUT83), .B(G559), .Z(new_n631));
  OAI21_X1  g206(.A(new_n624), .B1(G860), .B2(new_n631), .ZN(G148));
  NAND2_X1  g207(.A1(new_n624), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G868), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(G868), .B2(new_n570), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n499), .A2(new_n500), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(new_n462), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2100), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n488), .A2(G123), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n484), .A2(G135), .ZN(new_n643));
  OAI221_X1 g218(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n468), .C2(G111), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2096), .Z(new_n646));
  NAND2_X1  g221(.A1(new_n641), .A2(new_n646), .ZN(G156));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2435), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2438), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(KEYINPUT14), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT16), .B(G1341), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n656), .B(new_n658), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(G14), .B1(new_n653), .B2(new_n659), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT84), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT85), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  AND3_X1   g244(.A1(new_n667), .A2(KEYINPUT17), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n669), .B1(new_n667), .B2(KEYINPUT17), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n664), .A2(new_n666), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n669), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT18), .ZN(new_n675));
  OR3_X1    g250(.A1(new_n673), .A2(new_n675), .A3(G2100), .ZN(new_n676));
  OAI21_X1  g251(.A(G2100), .B1(new_n673), .B2(new_n675), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT86), .B(G2096), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n676), .A2(new_n677), .A3(new_n679), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G227));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  XOR2_X1   g260(.A(G1961), .B(G1966), .Z(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1971), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n685), .A2(new_n686), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n688), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT20), .ZN(new_n695));
  OAI221_X1 g270(.A(new_n692), .B1(new_n690), .B2(new_n688), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n695), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT87), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n697), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1991), .B(G1996), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT88), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n700), .B(new_n704), .Z(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(G229));
  NOR2_X1   g281(.A1(G16), .A2(G23), .ZN(new_n707));
  INV_X1    g282(.A(G288), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(G16), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT33), .B(G1976), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(G16), .A2(G22), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G166), .B2(G16), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT92), .B(G1971), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G6), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n601), .A2(G651), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n558), .A2(G48), .ZN(new_n720));
  AND3_X1   g295(.A1(new_n719), .A2(new_n603), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n718), .B1(new_n721), .B2(new_n717), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT32), .B(G1981), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n716), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT34), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n716), .A2(new_n726), .A3(KEYINPUT34), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G25), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n488), .A2(G119), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT89), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n484), .A2(G131), .ZN(new_n736));
  OAI221_X1 g311(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n468), .C2(G107), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n733), .B1(new_n740), .B2(new_n732), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT35), .B(G1991), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n741), .B(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n717), .A2(G24), .ZN(new_n745));
  INV_X1    g320(.A(G290), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(new_n717), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G1986), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(G1986), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n744), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n731), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT36), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n732), .A2(G33), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT25), .Z(new_n756));
  AND2_X1   g331(.A1(new_n637), .A2(G127), .ZN(new_n757));
  NAND2_X1  g332(.A1(G115), .A2(G2104), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n466), .B(new_n467), .C1(new_n757), .C2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G139), .ZN(new_n761));
  INV_X1    g336(.A(new_n484), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n756), .B(new_n760), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n754), .B1(new_n764), .B2(new_n732), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2072), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n570), .A2(G16), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G16), .B2(G19), .ZN(new_n768));
  INV_X1    g343(.A(G1341), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT30), .B(G28), .ZN(new_n771));
  OR2_X1    g346(.A1(KEYINPUT31), .A2(G11), .ZN(new_n772));
  NAND2_X1  g347(.A1(KEYINPUT31), .A2(G11), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n771), .A2(new_n732), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n645), .B2(new_n732), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT97), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n768), .A2(new_n769), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n770), .A2(new_n777), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT24), .ZN(new_n781));
  INV_X1    g356(.A(G34), .ZN(new_n782));
  AOI21_X1  g357(.A(G29), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n781), .B2(new_n782), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G160), .B2(new_n732), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n785), .A2(G2084), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n766), .A2(new_n780), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G16), .A2(G21), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G168), .B2(G16), .ZN(new_n789));
  INV_X1    g364(.A(G1966), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G29), .A2(G32), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n484), .A2(G141), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT95), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n462), .A2(G105), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT96), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n488), .A2(G129), .ZN(new_n797));
  NAND3_X1  g372(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT26), .Z(new_n799));
  NAND3_X1  g374(.A1(new_n796), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n794), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n792), .B1(new_n801), .B2(G29), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT27), .B(G1996), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G2084), .B2(new_n785), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n787), .A2(new_n791), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n732), .A2(G26), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n484), .A2(G140), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT94), .ZN(new_n809));
  OAI221_X1 g384(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n468), .C2(G116), .ZN(new_n810));
  INV_X1    g385(.A(G128), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n489), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n807), .B1(new_n813), .B2(new_n732), .ZN(new_n814));
  MUX2_X1   g389(.A(new_n807), .B(new_n814), .S(KEYINPUT28), .Z(new_n815));
  INV_X1    g390(.A(G2067), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n717), .A2(G4), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n624), .B2(new_n717), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT93), .B(G1348), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(G27), .A2(G29), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G164), .B2(G29), .ZN(new_n823));
  INV_X1    g398(.A(G2078), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(G5), .A2(G16), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(G171), .B2(G16), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(G1961), .Z(new_n828));
  NAND4_X1  g403(.A1(new_n817), .A2(new_n821), .A3(new_n825), .A4(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(G2090), .ZN(new_n830));
  NOR2_X1   g405(.A1(G29), .A2(G35), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(G162), .B2(G29), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n832), .B(new_n834), .ZN(new_n835));
  AOI211_X1 g410(.A(new_n806), .B(new_n829), .C1(new_n830), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n717), .A2(G20), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT100), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT23), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(G299), .B2(G16), .ZN(new_n840));
  INV_X1    g415(.A(G1956), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT99), .ZN(new_n843));
  OR3_X1    g418(.A1(new_n835), .A2(new_n843), .A3(new_n830), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n843), .B1(new_n835), .B2(new_n830), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT101), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI211_X1 g423(.A(KEYINPUT101), .B(new_n842), .C1(new_n844), .C2(new_n845), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n753), .B(new_n836), .C1(new_n848), .C2(new_n849), .ZN(G150));
  INV_X1    g425(.A(G150), .ZN(G311));
  NAND2_X1  g426(.A1(G80), .A2(G543), .ZN(new_n852));
  INV_X1    g427(.A(G67), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n519), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(G651), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n526), .A2(G93), .A3(new_n516), .A4(new_n518), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT103), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n526), .A2(G55), .A3(G543), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n857), .B1(new_n856), .B2(new_n858), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n855), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(G860), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(KEYINPUT37), .Z(new_n863));
  NAND2_X1  g438(.A1(new_n624), .A2(G559), .ZN(new_n864));
  XNOR2_X1  g439(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT104), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n570), .B1(new_n861), .B2(new_n867), .ZN(new_n868));
  OAI211_X1 g443(.A(KEYINPUT104), .B(new_n855), .C1(new_n859), .C2(new_n860), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n861), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n871), .A2(KEYINPUT104), .A3(new_n570), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n866), .B(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT105), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(G860), .B1(new_n874), .B2(new_n875), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR3_X1   g453(.A1(new_n874), .A2(KEYINPUT105), .A3(new_n875), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n863), .B1(new_n878), .B2(new_n879), .ZN(G145));
  XNOR2_X1  g455(.A(new_n813), .B(new_n512), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n881), .A2(new_n801), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n801), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n764), .A2(KEYINPUT106), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n763), .B(KEYINPUT106), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n887), .B1(new_n882), .B2(new_n883), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n739), .B(new_n639), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n488), .A2(G130), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n484), .A2(G142), .ZN(new_n891));
  OAI221_X1 g466(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n468), .C2(G118), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n889), .B(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n886), .A2(new_n888), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(G162), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n897), .A2(new_n645), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n645), .ZN(new_n899));
  OAI22_X1  g474(.A1(new_n898), .A2(new_n899), .B1(new_n481), .B2(new_n480), .ZN(new_n900));
  XNOR2_X1  g475(.A(G162), .B(new_n645), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(G160), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n896), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n886), .A2(new_n888), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n894), .ZN(new_n906));
  AOI21_X1  g481(.A(G37), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n905), .B1(new_n908), .B2(new_n895), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n886), .A2(KEYINPUT107), .A3(new_n888), .A4(new_n894), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n909), .A2(new_n910), .A3(new_n902), .A4(new_n900), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g488(.A1(new_n861), .A2(new_n627), .ZN(new_n914));
  XNOR2_X1  g489(.A(G299), .B(new_n623), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n915), .B(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n870), .A2(new_n872), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(new_n633), .ZN(new_n919));
  MUX2_X1   g494(.A(new_n917), .B(new_n915), .S(new_n919), .Z(new_n920));
  NOR2_X1   g495(.A1(G290), .A2(G305), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n609), .A2(KEYINPUT82), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n612), .A2(new_n611), .A3(new_n607), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n721), .B1(new_n924), .B2(new_n606), .ZN(new_n925));
  NOR3_X1   g500(.A1(new_n921), .A2(new_n925), .A3(G166), .ZN(new_n926));
  NAND2_X1  g501(.A1(G290), .A2(G305), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(new_n721), .A3(new_n606), .ZN(new_n928));
  AOI21_X1  g503(.A(G303), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(G288), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(G166), .B1(new_n921), .B2(new_n925), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n927), .A2(G303), .A3(new_n928), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n708), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT42), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n926), .A2(new_n929), .A3(G288), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n708), .B1(new_n931), .B2(new_n932), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n930), .A2(KEYINPUT108), .A3(new_n933), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n934), .B1(new_n940), .B2(KEYINPUT42), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n920), .B(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n914), .B1(new_n942), .B2(new_n627), .ZN(G295));
  OAI21_X1  g518(.A(new_n914), .B1(new_n942), .B2(new_n627), .ZN(G331));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n588), .A2(G171), .A3(new_n589), .ZN(new_n947));
  NAND2_X1  g522(.A1(G301), .A2(G168), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n873), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n918), .A2(new_n947), .A3(new_n948), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n915), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(new_n949), .B2(new_n873), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n950), .A2(new_n951), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n956), .B1(new_n957), .B2(new_n955), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n940), .B(new_n954), .C1(new_n958), .C2(new_n917), .ZN(new_n959));
  INV_X1    g534(.A(G37), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n958), .A2(new_n953), .ZN(new_n962));
  OR2_X1    g537(.A1(new_n952), .A2(new_n917), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n940), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n946), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n940), .ZN(new_n966));
  AOI211_X1 g541(.A(new_n915), .B(new_n956), .C1(new_n957), .C2(new_n955), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n952), .A2(new_n917), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n969), .A2(KEYINPUT111), .A3(new_n960), .A4(new_n959), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n945), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n954), .B1(new_n958), .B2(new_n917), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n972), .A2(new_n966), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n961), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT43), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT44), .B1(new_n971), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT43), .B1(new_n973), .B2(new_n961), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n969), .A2(new_n945), .A3(new_n960), .A4(new_n959), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(KEYINPUT110), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n975), .A2(new_n982), .A3(new_n945), .A4(new_n969), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n980), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n977), .A2(new_n984), .ZN(G397));
  INV_X1    g560(.A(G1384), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n510), .A2(G2105), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n462), .A2(G102), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n494), .A2(KEYINPUT4), .B1(new_n501), .B2(new_n503), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n986), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G40), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n480), .A2(new_n995), .A3(new_n481), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n813), .B(G2067), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n801), .B(G1996), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n739), .B(new_n742), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(G290), .B(G1986), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n998), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(G1384), .B1(new_n505), .B2(new_n511), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n996), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI211_X1 g584(.A(KEYINPUT50), .B(G1384), .C1(new_n505), .C2(new_n511), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OR2_X1    g586(.A1(new_n1011), .A2(G1348), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n996), .A2(new_n1007), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n816), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(KEYINPUT45), .B(new_n986), .C1(new_n989), .C2(new_n990), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n993), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n991), .A2(new_n1017), .A3(new_n992), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT56), .B(G2072), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1019), .A2(new_n1020), .A3(new_n996), .A4(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT57), .ZN(new_n1023));
  XNOR2_X1  g598(.A(G299), .B(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n991), .A2(KEYINPUT50), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n1026), .A3(new_n996), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n841), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1022), .A2(new_n1024), .A3(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1015), .A2(new_n1029), .A3(new_n624), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1022), .A2(new_n1028), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1024), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT60), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n624), .B1(new_n1015), .B2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1012), .A2(KEYINPUT60), .A3(new_n623), .A4(new_n1014), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1036), .A2(new_n1037), .B1(new_n1035), .B2(new_n1015), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT61), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1022), .A2(new_n1024), .A3(new_n1028), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1024), .B1(new_n1022), .B2(new_n1028), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1019), .A2(new_n996), .A3(new_n1020), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT58), .B(G1341), .ZN(new_n1044));
  OAI22_X1  g619(.A1(new_n1043), .A2(G1996), .B1(new_n1013), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n570), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT59), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1033), .A2(KEYINPUT61), .A3(new_n1029), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1045), .A2(KEYINPUT59), .A3(new_n570), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1042), .A2(new_n1048), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT121), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1038), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1054), .A2(KEYINPUT121), .A3(new_n1049), .A4(new_n1042), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1034), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1019), .A2(new_n1020), .A3(new_n824), .A4(new_n996), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT123), .B(G1961), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1058), .A2(new_n1059), .B1(new_n1027), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1016), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n512), .A2(KEYINPUT120), .A3(KEYINPUT45), .A4(new_n986), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1063), .A2(new_n993), .A3(new_n996), .A4(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n1066));
  OR3_X1    g641(.A1(new_n1065), .A2(new_n1066), .A3(G2078), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1061), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1057), .B1(new_n1068), .B2(G301), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1027), .A2(new_n1060), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n473), .A2(new_n463), .ZN(new_n1072));
  NOR4_X1   g647(.A1(new_n478), .A2(new_n1066), .A3(new_n995), .A4(G2078), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n993), .A2(new_n1072), .A3(new_n1016), .A4(new_n1073), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1070), .A2(new_n1071), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT126), .ZN(new_n1076));
  OAI21_X1  g651(.A(G171), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1061), .A2(new_n1074), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(KEYINPUT126), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1069), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT125), .B1(new_n1078), .B2(G171), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT125), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1061), .A2(new_n1082), .A3(G301), .A4(new_n1074), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1068), .A2(G171), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1081), .A2(new_n1057), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT49), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT116), .B(G86), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n546), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n719), .A2(new_n1090), .A3(new_n720), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G1981), .ZN(new_n1092));
  INV_X1    g667(.A(G1981), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n602), .A2(new_n1093), .A3(new_n603), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1088), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1093), .B1(new_n602), .B2(new_n1090), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1096), .A2(KEYINPUT117), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1087), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n602), .A2(new_n1093), .A3(new_n603), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT117), .B1(new_n1099), .B2(new_n1096), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1092), .A2(new_n1088), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1100), .A2(KEYINPUT49), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G8), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1013), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1098), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT118), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1098), .A2(new_n1102), .A3(new_n1104), .A4(new_n1107), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT114), .B(G1976), .Z(new_n1109));
  NOR2_X1   g684(.A1(new_n708), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT52), .B1(new_n1104), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n708), .B2(G1976), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1104), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1104), .B(new_n1113), .C1(KEYINPUT52), .C2(new_n1110), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1106), .A2(new_n1108), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(G303), .A2(G8), .ZN(new_n1118));
  NAND2_X1  g693(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1121), .B1(new_n1118), .B2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1027), .A2(G2090), .ZN(new_n1126));
  INV_X1    g701(.A(G1971), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1126), .B1(new_n1127), .B2(new_n1043), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1125), .B1(new_n1128), .B2(new_n1103), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1125), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1043), .A2(new_n1127), .ZN(new_n1131));
  OAI211_X1 g706(.A(G8), .B(new_n1130), .C1(new_n1131), .C2(new_n1126), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1117), .A2(new_n1129), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1065), .A2(new_n790), .ZN(new_n1134));
  INV_X1    g709(.A(G2084), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1025), .A2(new_n1026), .A3(new_n1135), .A4(new_n996), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(G168), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1137), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT122), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1137), .A2(new_n1140), .A3(KEYINPUT51), .A4(G8), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n790), .A2(new_n1065), .B1(new_n1011), .B2(new_n1135), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1103), .B1(new_n1142), .B2(G168), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1139), .B(new_n1141), .C1(KEYINPUT51), .C2(new_n1143), .ZN(new_n1144));
  OR3_X1    g719(.A1(new_n1142), .A2(new_n1103), .A3(G168), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1133), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1086), .A2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1056), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1141), .B1(new_n1143), .B2(KEYINPUT51), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1140), .B1(new_n1143), .B2(KEYINPUT51), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1145), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT62), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT62), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1144), .A2(new_n1153), .A3(new_n1145), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1133), .A2(new_n1084), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1152), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1142), .A2(new_n1103), .A3(G286), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1117), .A2(new_n1129), .A3(new_n1132), .A4(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT63), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1158), .B(new_n1159), .ZN(new_n1160));
  OR2_X1    g735(.A1(G288), .A2(G1976), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1161), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1104), .B1(new_n1162), .B2(new_n1099), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT119), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1128), .A2(new_n1103), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .A4(new_n1130), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n1163), .A2(new_n1164), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1164), .B1(new_n1163), .B2(new_n1168), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1156), .A2(new_n1160), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1006), .B1(new_n1148), .B2(new_n1172), .ZN(new_n1173));
  NOR3_X1   g748(.A1(new_n997), .A2(G1986), .A3(G290), .ZN(new_n1174));
  OAI22_X1  g749(.A1(new_n1003), .A2(new_n997), .B1(KEYINPUT48), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1175), .B1(KEYINPUT48), .B2(new_n1174), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n997), .B1(new_n999), .B2(new_n801), .ZN(new_n1177));
  INV_X1    g752(.A(G1996), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT46), .B1(new_n998), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT46), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n997), .A2(new_n1180), .A3(G1996), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1177), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT47), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n813), .A2(new_n816), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n740), .A2(new_n743), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1184), .B1(new_n1001), .B2(new_n1185), .ZN(new_n1186));
  AOI211_X1 g761(.A(new_n1176), .B(new_n1183), .C1(new_n998), .C2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1173), .A2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g763(.A(G319), .B1(new_n660), .B2(new_n661), .ZN(new_n1190));
  INV_X1    g764(.A(new_n1190), .ZN(new_n1191));
  AOI21_X1  g765(.A(KEYINPUT127), .B1(new_n683), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n1193));
  AOI211_X1 g767(.A(new_n1193), .B(new_n1190), .C1(new_n681), .C2(new_n682), .ZN(new_n1194));
  OAI21_X1  g768(.A(new_n705), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g769(.A(new_n1195), .B1(new_n907), .B2(new_n911), .ZN(new_n1196));
  NAND3_X1  g770(.A1(new_n1196), .A2(new_n980), .A3(new_n983), .ZN(G225));
  INV_X1    g771(.A(G225), .ZN(G308));
endmodule


