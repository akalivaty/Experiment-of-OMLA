//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 1 1 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  OR4_X1    g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n462), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n474), .A2(KEYINPUT69), .A3(G137), .A4(new_n462), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n464), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n477), .B1(new_n472), .B2(new_n473), .ZN(new_n478));
  AND2_X1   g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  OAI21_X1  g054(.A(G2105), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n462), .B1(new_n472), .B2(new_n473), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT70), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n474), .A2(new_n462), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI211_X1 g065(.A(new_n485), .B(new_n488), .C1(G136), .C2(new_n490), .ZN(G162));
  OAI211_X1 g066(.A(G138), .B(new_n462), .C1(new_n465), .C2(new_n466), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n474), .A2(new_n494), .A3(G138), .A4(new_n462), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n462), .A2(G114), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OR2_X1    g075(.A1(G102), .A2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n501), .A2(new_n503), .A3(KEYINPUT71), .A4(G2104), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n500), .A2(new_n504), .B1(new_n486), .B2(G126), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n496), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT72), .B1(new_n508), .B2(KEYINPUT6), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n510), .A2(new_n511), .A3(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT73), .B(G88), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n513), .A2(new_n514), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n513), .A2(G543), .A3(new_n514), .ZN(new_n520));
  OAI221_X1 g095(.A(new_n517), .B1(new_n518), .B2(new_n508), .C1(new_n519), .C2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  AOI22_X1  g097(.A1(new_n509), .A2(new_n512), .B1(KEYINPUT6), .B2(new_n508), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n523), .A2(G89), .A3(new_n515), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(G51), .A3(G543), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n528));
  AND2_X1   g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n527), .A2(new_n528), .B1(new_n515), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n524), .A2(new_n525), .A3(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  XOR2_X1   g107(.A(KEYINPUT74), .B(G52), .Z(new_n533));
  NAND3_X1  g108(.A1(new_n523), .A2(G543), .A3(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n537));
  OAI221_X1 g112(.A(new_n534), .B1(new_n535), .B2(new_n508), .C1(new_n536), .C2(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  INV_X1    g114(.A(new_n520), .ZN(new_n540));
  AND3_X1   g115(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n540), .A2(G43), .B1(new_n541), .B2(G81), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n508), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR3_X1   g121(.A1(new_n543), .A2(KEYINPUT75), .A3(new_n508), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n542), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NOR2_X1   g129(.A1(KEYINPUT78), .A2(G65), .ZN(new_n555));
  AND2_X1   g130(.A1(KEYINPUT78), .A2(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n515), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT77), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n508), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(G91), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT76), .B1(new_n537), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n523), .A2(new_n563), .A3(G91), .A4(new_n515), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n560), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n513), .A2(G53), .A3(G543), .A4(new_n514), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT79), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n565), .A2(new_n567), .A3(KEYINPUT79), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G299));
  NAND4_X1  g148(.A1(new_n513), .A2(G49), .A3(G543), .A4(new_n514), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n513), .A2(G87), .A3(new_n514), .A4(new_n515), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  AND2_X1   g152(.A1(KEYINPUT5), .A2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(KEYINPUT5), .A2(G543), .ZN(new_n579));
  OAI21_X1  g154(.A(G61), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n508), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT80), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n582), .B(new_n583), .ZN(new_n584));
  AND2_X1   g159(.A1(G48), .A2(G543), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n513), .A2(new_n514), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(KEYINPUT81), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT81), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n523), .A2(new_n588), .A3(new_n585), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n587), .A2(new_n589), .B1(new_n541), .B2(G86), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n584), .A2(new_n590), .ZN(G305));
  NAND2_X1  g166(.A1(new_n540), .A2(G47), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n541), .A2(G85), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n592), .B(new_n593), .C1(new_n508), .C2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  INV_X1    g171(.A(G54), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n597), .B1(new_n520), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(new_n598), .B2(new_n520), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n513), .A2(G92), .A3(new_n514), .A4(new_n515), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n601), .B(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n604), .A2(new_n508), .ZN(new_n605));
  AND3_X1   g180(.A1(new_n600), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n596), .B1(new_n606), .B2(G868), .ZN(G284));
  OAI21_X1  g182(.A(new_n596), .B1(new_n606), .B2(G868), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(new_n572), .B2(G868), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(new_n572), .B2(G868), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n606), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n606), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g192(.A1(new_n465), .A2(new_n466), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n462), .A2(G2104), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n487), .A2(G123), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n490), .A2(G135), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n462), .A2(G111), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n624), .B(new_n625), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n623), .A2(G2100), .B1(G2096), .B2(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(G2096), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n629), .B(new_n630), .C1(G2100), .C2(new_n623), .ZN(G156));
  INV_X1    g206(.A(KEYINPUT14), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n635), .B2(new_n634), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n637), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  AND3_X1   g220(.A1(new_n644), .A2(G14), .A3(new_n645), .ZN(G401));
  INV_X1    g221(.A(KEYINPUT18), .ZN(new_n647));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(KEYINPUT17), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n648), .A2(new_n649), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n647), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2100), .ZN(new_n654));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n650), .B2(KEYINPUT18), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2096), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n654), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1971), .B(G1976), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  XOR2_X1   g235(.A(G1956), .B(G2474), .Z(new_n661));
  XOR2_X1   g236(.A(G1961), .B(G1966), .Z(new_n662));
  AND2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT20), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n661), .A2(new_n662), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n660), .A2(new_n663), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n660), .B2(new_n666), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1991), .B(G1996), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1981), .B(G1986), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G229));
  NAND3_X1  g250(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT25), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(G139), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(new_n679), .B2(new_n489), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n680), .A2(KEYINPUT90), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(KEYINPUT90), .ZN(new_n682));
  NAND2_X1  g257(.A1(G115), .A2(G2104), .ZN(new_n683));
  INV_X1    g258(.A(G127), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(new_n618), .B2(new_n684), .ZN(new_n685));
  AOI22_X1  g260(.A1(new_n681), .A2(new_n682), .B1(G2105), .B2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n687), .B2(G33), .ZN(new_n689));
  INV_X1    g264(.A(G2072), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT91), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n687), .A2(G32), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n487), .A2(G129), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT93), .Z(new_n695));
  NAND3_X1  g270(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT26), .Z(new_n697));
  INV_X1    g272(.A(G105), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(new_n619), .ZN(new_n699));
  INV_X1    g274(.A(G141), .ZN(new_n700));
  OAI21_X1  g275(.A(KEYINPUT92), .B1(new_n489), .B2(new_n700), .ZN(new_n701));
  OR3_X1    g276(.A1(new_n489), .A2(KEYINPUT92), .A3(new_n700), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n695), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n693), .B1(new_n704), .B2(G29), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT27), .B(G1996), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n689), .A2(new_n690), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n687), .A2(G27), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G164), .B2(new_n687), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G2078), .ZN(new_n711));
  NOR3_X1   g286(.A1(new_n707), .A2(new_n708), .A3(new_n711), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n705), .A2(new_n706), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n687), .B1(KEYINPUT24), .B2(G34), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(KEYINPUT24), .B2(G34), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n481), .B2(G29), .ZN(new_n716));
  INV_X1    g291(.A(G2084), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NOR2_X1   g295(.A1(G171), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G5), .B2(new_n720), .ZN(new_n722));
  INV_X1    g297(.A(G1961), .ZN(new_n723));
  AOI211_X1 g298(.A(new_n718), .B(new_n719), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n692), .A2(new_n712), .A3(new_n713), .A4(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n720), .A2(G21), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G168), .B2(new_n720), .ZN(new_n727));
  OAI22_X1  g302(.A1(new_n722), .A2(new_n723), .B1(G1966), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(G1966), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT30), .B(G28), .ZN(new_n730));
  OR2_X1    g305(.A1(KEYINPUT31), .A2(G11), .ZN(new_n731));
  NAND2_X1  g306(.A1(KEYINPUT31), .A2(G11), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n730), .A2(new_n687), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n729), .B(new_n733), .C1(new_n687), .C2(new_n628), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n728), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT94), .Z(new_n736));
  INV_X1    g311(.A(KEYINPUT95), .ZN(new_n737));
  OR3_X1    g312(.A1(new_n725), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n720), .A2(G22), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G166), .B2(new_n720), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(G1971), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(G1971), .ZN(new_n742));
  OR2_X1    g317(.A1(G6), .A2(G16), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G305), .B2(new_n720), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT32), .B(G1981), .Z(new_n745));
  OAI211_X1 g320(.A(new_n741), .B(new_n742), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(G288), .A2(KEYINPUT86), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT86), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n574), .A2(new_n575), .A3(new_n748), .A4(new_n576), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  MUX2_X1   g325(.A(G23), .B(new_n750), .S(G16), .Z(new_n751));
  XOR2_X1   g326(.A(KEYINPUT33), .B(G1976), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n746), .B(new_n753), .C1(new_n744), .C2(new_n745), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT34), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT36), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(KEYINPUT87), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n754), .A2(new_n755), .ZN(new_n759));
  MUX2_X1   g334(.A(G24), .B(G290), .S(G16), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT85), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1986), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n687), .A2(G25), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n487), .A2(G119), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT84), .ZN(new_n765));
  OAI21_X1  g340(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n766));
  INV_X1    g341(.A(G107), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(G2105), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n490), .B2(G131), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n763), .B1(new_n771), .B2(new_n687), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT35), .B(G1991), .Z(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n772), .B(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n757), .A2(KEYINPUT87), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n762), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n756), .A2(new_n758), .A3(new_n759), .A4(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G4), .A2(G16), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n606), .B2(G16), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT88), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT89), .B(G1348), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n781), .B(new_n782), .Z(new_n783));
  XOR2_X1   g358(.A(KEYINPUT96), .B(KEYINPUT23), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n720), .A2(G20), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n572), .B2(new_n720), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1956), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n687), .A2(G35), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G162), .B2(new_n687), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT29), .B(G2090), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n687), .A2(G26), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT28), .Z(new_n794));
  NAND2_X1  g369(.A1(new_n487), .A2(G128), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n490), .A2(G140), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n462), .A2(G116), .ZN(new_n797));
  OAI21_X1  g372(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n795), .B(new_n796), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n794), .B1(new_n799), .B2(G29), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G2067), .ZN(new_n801));
  NOR2_X1   g376(.A1(G16), .A2(G19), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n549), .B2(G16), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(G1341), .Z(new_n804));
  NAND3_X1  g379(.A1(new_n792), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n783), .A2(new_n788), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n737), .B1(new_n725), .B2(new_n736), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n738), .A2(new_n778), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n756), .A2(new_n759), .A3(new_n777), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n809), .A2(KEYINPUT87), .A3(new_n757), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n808), .A2(new_n811), .ZN(G311));
  INV_X1    g387(.A(G311), .ZN(G150));
  NAND2_X1  g388(.A1(new_n606), .A2(G559), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT38), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n515), .A2(G67), .ZN(new_n816));
  AND2_X1   g391(.A1(G80), .A2(G543), .ZN(new_n817));
  OAI21_X1  g392(.A(G651), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n523), .A2(G55), .A3(G543), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n513), .A2(G93), .A3(new_n514), .A4(new_n515), .ZN(new_n820));
  AND3_X1   g395(.A1(new_n819), .A2(new_n820), .A3(KEYINPUT97), .ZN(new_n821));
  AOI21_X1  g396(.A(KEYINPUT97), .B1(new_n819), .B2(new_n820), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n818), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(new_n549), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n548), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n815), .B(new_n827), .Z(new_n828));
  AND2_X1   g403(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n829), .A2(new_n830), .A3(G860), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n823), .A2(G860), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT37), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n831), .A2(new_n833), .ZN(G145));
  XOR2_X1   g409(.A(KEYINPUT98), .B(G37), .Z(new_n835));
  NAND2_X1  g410(.A1(new_n487), .A2(G130), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n490), .A2(G142), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n462), .A2(G118), .ZN(new_n838));
  OAI21_X1  g413(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n839));
  OAI211_X1 g414(.A(new_n836), .B(new_n837), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n770), .B(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n686), .B1(new_n695), .B2(new_n703), .ZN(new_n842));
  AND3_X1   g417(.A1(new_n695), .A2(new_n703), .A3(new_n686), .ZN(new_n843));
  OR3_X1    g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n799), .B(new_n506), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n622), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n628), .B(new_n481), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G162), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n844), .A2(new_n845), .A3(new_n848), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n850), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n853), .B1(new_n850), .B2(new_n854), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n835), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g433(.A(new_n827), .B(new_n614), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n570), .A2(new_n571), .A3(new_n606), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT99), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n570), .A2(new_n606), .A3(KEYINPUT99), .A4(new_n571), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n606), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n572), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n859), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT41), .B1(new_n866), .B2(new_n860), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n606), .B1(new_n570), .B2(new_n571), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT41), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n869), .B1(new_n864), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n868), .B1(new_n873), .B2(new_n859), .ZN(new_n874));
  XNOR2_X1  g449(.A(G305), .B(G166), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n750), .B(G290), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n875), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT42), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n874), .B(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(G868), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(G868), .B2(new_n824), .ZN(G295));
  OAI21_X1  g456(.A(new_n880), .B1(G868), .B2(new_n824), .ZN(G331));
  INV_X1    g457(.A(KEYINPUT44), .ZN(new_n883));
  INV_X1    g458(.A(new_n877), .ZN(new_n884));
  XNOR2_X1  g459(.A(G301), .B(G286), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n823), .A2(new_n548), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n823), .A2(new_n548), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(G301), .B(G168), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n825), .A2(new_n889), .A3(new_n826), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT101), .B1(new_n867), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n870), .B1(new_n862), .B2(new_n863), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n895));
  NOR3_X1   g470(.A1(new_n894), .A2(new_n895), .A3(new_n891), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n872), .A2(new_n860), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(new_n894), .B2(KEYINPUT41), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT100), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n825), .A2(new_n889), .A3(new_n900), .A4(new_n826), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n888), .A2(new_n890), .A3(KEYINPUT100), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n884), .B1(new_n897), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n901), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n867), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n906), .B(new_n884), .C1(new_n873), .C2(new_n892), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n835), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT43), .B1(new_n904), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n883), .B1(new_n909), .B2(KEYINPUT103), .ZN(new_n910));
  INV_X1    g485(.A(G37), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n864), .A2(new_n872), .ZN(new_n915));
  INV_X1    g490(.A(new_n860), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n871), .B1(new_n916), .B2(new_n870), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n892), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n894), .B1(new_n901), .B2(new_n902), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n877), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n912), .A2(new_n913), .A3(new_n914), .A4(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(new_n907), .A3(new_n911), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT102), .B1(new_n922), .B2(KEYINPUT43), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n925), .B(KEYINPUT43), .C1(new_n904), .C2(new_n908), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n910), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n897), .A2(new_n903), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n877), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n929), .A2(new_n914), .A3(new_n835), .A4(new_n907), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n883), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n927), .A2(new_n933), .ZN(G397));
  INV_X1    g509(.A(G1384), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT45), .B1(new_n506), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT45), .ZN(new_n937));
  AOI211_X1 g512(.A(new_n937), .B(G1384), .C1(new_n496), .C2(new_n505), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n469), .A2(new_n475), .ZN(new_n940));
  AND4_X1   g515(.A1(G40), .A2(new_n940), .A3(new_n480), .A4(new_n463), .ZN(new_n941));
  AOI21_X1  g516(.A(G1966), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n506), .A2(new_n935), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n941), .ZN(new_n945));
  AOI21_X1  g520(.A(G1384), .B1(new_n496), .B2(new_n505), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT50), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n945), .A2(G2084), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(G286), .B1(new_n942), .B2(new_n949), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n940), .A2(G40), .A3(new_n480), .A4(new_n463), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n951), .B1(new_n946), .B2(new_n943), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n506), .A2(new_n935), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT50), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(new_n954), .A3(new_n717), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n936), .A2(new_n938), .A3(new_n951), .ZN(new_n956));
  OAI211_X1 g531(.A(G168), .B(new_n955), .C1(new_n956), .C2(G1966), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n950), .A2(KEYINPUT51), .A3(G8), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(G8), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT51), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT120), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT120), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n958), .A2(new_n961), .A3(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n963), .A2(KEYINPUT62), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT127), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT62), .ZN(new_n969));
  INV_X1    g544(.A(new_n965), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n964), .B1(new_n958), .B2(new_n961), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G8), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n973), .B1(new_n941), .B2(new_n946), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n586), .A2(KEYINPUT81), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n588), .B1(new_n523), .B2(new_n585), .ZN(new_n976));
  INV_X1    g551(.A(G86), .ZN(new_n977));
  OAI22_X1  g552(.A1(new_n975), .A2(new_n976), .B1(new_n977), .B2(new_n537), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n580), .A2(new_n581), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n583), .B1(new_n979), .B2(G651), .ZN(new_n980));
  AOI211_X1 g555(.A(KEYINPUT80), .B(new_n508), .C1(new_n580), .C2(new_n581), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(G1981), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1981), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n584), .A2(new_n590), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT111), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT49), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n974), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI211_X1 g563(.A(KEYINPUT111), .B(KEYINPUT49), .C1(new_n983), .C2(new_n985), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n747), .A2(G1976), .A3(new_n749), .ZN(new_n990));
  INV_X1    g565(.A(G40), .ZN(new_n991));
  AOI211_X1 g566(.A(new_n991), .B(new_n464), .C1(new_n469), .C2(new_n475), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n946), .A2(new_n992), .A3(new_n480), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n990), .A2(new_n993), .A3(G8), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n994), .A2(KEYINPUT109), .A3(KEYINPUT52), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT109), .B1(new_n994), .B2(KEYINPUT52), .ZN(new_n996));
  OAI22_X1  g571(.A1(new_n988), .A2(new_n989), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1976), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT52), .B1(G288), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n974), .A2(new_n990), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT110), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n974), .A2(new_n1002), .A3(new_n990), .A4(new_n999), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n997), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(KEYINPUT108), .B(KEYINPUT55), .ZN(new_n1007));
  AND3_X1   g582(.A1(G303), .A2(G8), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1007), .B1(G303), .B2(G8), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n953), .A2(new_n937), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n946), .A2(KEYINPUT45), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(new_n941), .A3(new_n1012), .ZN(new_n1013));
  XOR2_X1   g588(.A(KEYINPUT105), .B(G1971), .Z(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g591(.A(KEYINPUT107), .B(G2090), .Z(new_n1017));
  NAND3_X1  g592(.A1(new_n952), .A2(new_n954), .A3(new_n1017), .ZN(new_n1018));
  AOI211_X1 g593(.A(new_n973), .B(new_n1010), .C1(new_n1016), .C2(new_n1018), .ZN(new_n1019));
  OR2_X1    g594(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n946), .A2(new_n943), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n946), .A2(new_n947), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1021), .A2(new_n941), .A3(new_n1022), .A4(new_n1017), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n956), .B2(new_n1014), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1020), .B1(new_n1024), .B2(G8), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1019), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT125), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1006), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n974), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT111), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n978), .A2(new_n982), .A3(G1981), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n984), .B1(new_n584), .B2(new_n590), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1029), .B1(new_n1033), .B2(KEYINPUT49), .ZN(new_n1034));
  INV_X1    g609(.A(new_n989), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n994), .A2(KEYINPUT52), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT109), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n994), .A2(KEYINPUT109), .A3(KEYINPUT52), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1036), .A2(new_n1004), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1014), .B1(new_n939), .B2(new_n941), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n952), .A2(new_n954), .A3(new_n1017), .ZN(new_n1044));
  OAI211_X1 g619(.A(G8), .B(new_n1020), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n973), .B1(new_n1016), .B2(new_n1023), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1045), .B1(new_n1046), .B2(new_n1020), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT125), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(new_n945), .B2(new_n948), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n952), .A2(new_n954), .A3(KEYINPUT115), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n723), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G2078), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT53), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n956), .A2(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n1013), .B2(G2078), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1052), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G171), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1028), .A2(new_n1048), .A3(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n963), .A2(KEYINPUT127), .A3(KEYINPUT62), .A4(new_n965), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n968), .A2(new_n972), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1042), .A2(KEYINPUT112), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1034), .A2(new_n1035), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT112), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(new_n1067), .A3(new_n1004), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n942), .A2(new_n949), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1070), .A2(new_n973), .A3(G286), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1071), .A2(KEYINPUT63), .A3(new_n1045), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1020), .B1(new_n1073), .B2(G8), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1006), .A2(new_n1026), .A3(new_n1071), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT63), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1069), .A2(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1067), .B1(new_n1066), .B2(new_n1004), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n997), .A2(new_n1005), .A3(KEYINPUT112), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1019), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI211_X1 g656(.A(G1976), .B(G288), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n974), .B1(new_n1082), .B2(new_n1031), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1078), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT114), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT56), .B(G2072), .Z(new_n1087));
  NOR2_X1   g662(.A1(new_n1013), .A2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1022), .B(new_n941), .C1(new_n946), .C2(new_n943), .ZN(new_n1089));
  INV_X1    g664(.A(G1956), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT113), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT113), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1089), .A2(new_n1093), .A3(new_n1090), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1088), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n568), .B(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1086), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  OR2_X1    g673(.A1(new_n1013), .A2(new_n1087), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1089), .A2(new_n1093), .A3(new_n1090), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1093), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1097), .B(new_n1099), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1102), .A2(KEYINPUT114), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1098), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1050), .A2(new_n782), .A3(new_n1051), .ZN(new_n1105));
  INV_X1    g680(.A(new_n993), .ZN(new_n1106));
  INV_X1    g681(.A(G2067), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1109), .A2(KEYINPUT116), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT116), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1111), .A2(new_n606), .A3(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1097), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1104), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(KEYINPUT61), .A3(new_n1102), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT58), .B(G1341), .ZN(new_n1121));
  OAI22_X1  g696(.A1(new_n1013), .A2(G1996), .B1(new_n1106), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n548), .B1(KEYINPUT117), .B2(KEYINPUT59), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OR2_X1    g699(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1124), .B(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1120), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT118), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1116), .A2(new_n1129), .A3(new_n1117), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1128), .B(new_n1130), .C1(new_n1098), .C2(new_n1103), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1127), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT60), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT119), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1134), .B1(new_n606), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1137), .A2(KEYINPUT119), .A3(new_n865), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1111), .A2(new_n1134), .A3(new_n1114), .ZN(new_n1139));
  OAI221_X1 g714(.A(new_n1136), .B1(new_n1135), .B2(new_n606), .C1(new_n1110), .C2(new_n1113), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1119), .B1(new_n1133), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n1143));
  OR3_X1    g718(.A1(new_n478), .A2(new_n1143), .A3(new_n479), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1143), .B1(new_n478), .B2(new_n479), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1144), .A2(G2105), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n992), .A2(new_n1146), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n1147), .A2(KEYINPUT123), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(KEYINPUT123), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1148), .A2(new_n939), .A3(new_n1055), .A4(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1052), .A2(new_n1150), .A3(new_n1058), .A4(G301), .ZN(new_n1151));
  AOI21_X1  g726(.A(KEYINPUT54), .B1(new_n1060), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI211_X1 g729(.A(KEYINPUT124), .B(KEYINPUT54), .C1(new_n1060), .C2(new_n1151), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1052), .A2(new_n1058), .A3(new_n1150), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(G171), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1052), .A2(G301), .A3(new_n1058), .A4(new_n1056), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1158), .A2(KEYINPUT54), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(KEYINPUT126), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT126), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1158), .A2(new_n1162), .A3(KEYINPUT54), .A4(new_n1159), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1027), .B1(new_n1006), .B2(new_n1026), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1042), .A2(new_n1047), .A3(KEYINPUT125), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n970), .A2(new_n971), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1156), .A2(new_n1164), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1064), .B(new_n1085), .C1(new_n1142), .C2(new_n1169), .ZN(new_n1170));
  OR3_X1    g745(.A1(new_n1011), .A2(G1996), .A3(new_n951), .ZN(new_n1171));
  XOR2_X1   g746(.A(new_n1171), .B(KEYINPUT104), .Z(new_n1172));
  NOR2_X1   g747(.A1(new_n1011), .A2(new_n951), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n704), .A2(G1996), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n799), .B(new_n1107), .ZN(new_n1176));
  AND2_X1   g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  OAI22_X1  g752(.A1(new_n1172), .A2(new_n704), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n770), .B(new_n773), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1178), .B1(new_n1173), .B2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g756(.A(G290), .B(G1986), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n1173), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1170), .A2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1172), .B(KEYINPUT46), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1176), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1173), .B1(new_n1187), .B2(new_n704), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT47), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n1178), .A2(new_n774), .A3(new_n770), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n799), .A2(G2067), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1173), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NOR3_X1   g768(.A1(new_n1174), .A2(G1986), .A3(G290), .ZN(new_n1194));
  XOR2_X1   g769(.A(new_n1194), .B(KEYINPUT48), .Z(new_n1195));
  NAND2_X1  g770(.A1(new_n1181), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1190), .A2(new_n1193), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1185), .A2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g774(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1201));
  NAND3_X1  g775(.A1(new_n932), .A2(new_n1201), .A3(new_n857), .ZN(G225));
  INV_X1    g776(.A(G225), .ZN(G308));
endmodule


