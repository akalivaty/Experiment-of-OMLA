//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n448, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n560, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n639,
    new_n640, new_n642, new_n643, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1231, new_n1232, new_n1233;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n456), .A2(G2106), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n458), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  XNOR2_X1  g039(.A(KEYINPUT67), .B(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT67), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n469), .A2(new_n471), .A3(KEYINPUT3), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n472), .A2(G137), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n467), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n479), .B1(new_n481), .B2(G125), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n475), .A2(new_n480), .ZN(new_n483));
  INV_X1    g058(.A(G125), .ZN(new_n484));
  NOR3_X1   g059(.A1(new_n483), .A2(KEYINPUT66), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n478), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n477), .B1(new_n486), .B2(G2105), .ZN(G160));
  NOR2_X1   g062(.A1(new_n473), .A2(G112), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n472), .A2(new_n475), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G136), .ZN(new_n493));
  XOR2_X1   g068(.A(new_n493), .B(KEYINPUT68), .Z(new_n494));
  NOR2_X1   g069(.A1(new_n491), .A2(new_n473), .ZN(new_n495));
  AOI211_X1 g070(.A(new_n490), .B(new_n494), .C1(G124), .C2(new_n495), .ZN(G162));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  AND4_X1   g073(.A1(new_n473), .A2(new_n498), .A3(new_n475), .A4(new_n480), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n472), .A2(G138), .A3(new_n473), .A4(new_n475), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(KEYINPUT4), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n472), .A2(G126), .A3(G2105), .A4(new_n475), .ZN(new_n502));
  OR2_X1    g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n503), .B(G2104), .C1(G114), .C2(new_n473), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n501), .A2(new_n505), .ZN(G164));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  OR2_X1    g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n513), .A2(new_n514), .B1(new_n507), .B2(new_n508), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n519), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n516), .A2(new_n522), .ZN(G166));
  OAI211_X1 g098(.A(G51), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n524));
  OAI211_X1 g099(.A(G63), .B(G651), .C1(new_n514), .C2(new_n513), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT69), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT70), .B(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  OR2_X1    g106(.A1(KEYINPUT70), .A2(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(KEYINPUT70), .A2(KEYINPUT7), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n532), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n509), .A2(G89), .A3(new_n519), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n527), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n526), .B1(new_n524), .B2(new_n525), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(G168));
  AOI22_X1  g114(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n521), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n514), .A2(new_n513), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n507), .A2(new_n508), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  XOR2_X1   g121(.A(KEYINPUT71), .B(G52), .Z(new_n547));
  AOI22_X1  g122(.A1(G90), .A2(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n541), .A2(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  OAI211_X1 g125(.A(G43), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n515), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g128(.A(G56), .B1(new_n514), .B2(new_n513), .ZN(new_n554));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n521), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT72), .ZN(G153));
  AND3_X1   g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G36), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n542), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(G651), .A2(new_n567), .B1(new_n544), .B2(G91), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(KEYINPUT73), .ZN(new_n570));
  INV_X1    g145(.A(G53), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n510), .B2(new_n571), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n546), .B(G53), .C1(KEYINPUT73), .C2(new_n569), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n572), .A2(new_n573), .A3(KEYINPUT74), .ZN(new_n574));
  AOI21_X1  g149(.A(KEYINPUT74), .B1(new_n572), .B2(new_n573), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n568), .B1(new_n574), .B2(new_n575), .ZN(G299));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n577), .B1(new_n537), .B2(new_n538), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n544), .A2(G89), .B1(new_n531), .B2(new_n534), .ZN(new_n579));
  INV_X1    g154(.A(new_n538), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT75), .A4(new_n527), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G286));
  INV_X1    g158(.A(G166), .ZN(G303));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n585));
  INV_X1    g160(.A(G49), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n510), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n546), .A2(KEYINPUT76), .A3(G49), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n519), .A2(G74), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(new_n544), .B2(G87), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(G288));
  NAND2_X1  g167(.A1(new_n544), .A2(G86), .ZN(new_n593));
  XOR2_X1   g168(.A(new_n593), .B(KEYINPUT78), .Z(new_n594));
  INV_X1    g169(.A(KEYINPUT77), .ZN(new_n595));
  INV_X1    g170(.A(G61), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n542), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n519), .A2(KEYINPUT77), .A3(G61), .ZN(new_n598));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G651), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n546), .A2(G48), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n594), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(KEYINPUT79), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT79), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n594), .A2(new_n607), .A3(new_n604), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(G305));
  INV_X1    g185(.A(G47), .ZN(new_n611));
  INV_X1    g186(.A(G85), .ZN(new_n612));
  OAI22_X1  g187(.A1(new_n510), .A2(new_n611), .B1(new_n612), .B2(new_n515), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n614), .A2(new_n521), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n613), .A2(new_n615), .ZN(G290));
  NAND2_X1  g191(.A1(G301), .A2(G868), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT80), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(G66), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(G66), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n519), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G79), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n545), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n621), .B(KEYINPUT81), .C1(new_n622), .C2(new_n545), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(G651), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n544), .A2(KEYINPUT10), .A3(G92), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT10), .ZN(new_n629));
  INV_X1    g204(.A(G92), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n515), .B2(new_n630), .ZN(new_n631));
  AOI22_X1  g206(.A1(new_n628), .A2(new_n631), .B1(G54), .B2(new_n546), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n617), .B1(new_n634), .B2(G868), .ZN(G284));
  OAI21_X1  g210(.A(new_n617), .B1(new_n634), .B2(G868), .ZN(G321));
  MUX2_X1   g211(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g212(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g213(.A(G559), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n634), .B1(new_n639), .B2(G860), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT82), .ZN(G148));
  NAND2_X1  g216(.A1(new_n634), .A2(new_n639), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(G868), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g219(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR3_X1   g220(.A1(new_n483), .A2(new_n465), .A3(G2105), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT12), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT13), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2100), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n492), .A2(G135), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n495), .A2(G123), .ZN(new_n651));
  OR2_X1    g226(.A1(G99), .A2(G2105), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n652), .B(G2104), .C1(G111), .C2(new_n473), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n650), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(G2096), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n649), .A2(new_n655), .ZN(G156));
  XNOR2_X1  g231(.A(G2427), .B(G2438), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2430), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT15), .B(G2435), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(KEYINPUT14), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n668));
  XNOR2_X1  g243(.A(G2451), .B(G2454), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(G14), .B1(new_n667), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n671), .B2(new_n667), .ZN(G401));
  XOR2_X1   g248(.A(G2067), .B(G2678), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT84), .ZN(new_n675));
  XOR2_X1   g250(.A(G2084), .B(G2090), .Z(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2072), .B(G2078), .Z(new_n678));
  NOR3_X1   g253(.A1(new_n675), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT18), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(KEYINPUT17), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n681), .A2(new_n675), .A3(new_n676), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n676), .B1(new_n675), .B2(new_n678), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT85), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(new_n675), .B2(new_n681), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n680), .B(new_n682), .C1(new_n685), .C2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G2096), .B(G2100), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G227));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT19), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G1956), .B(G2474), .Z(new_n695));
  XOR2_X1   g270(.A(G1961), .B(G1966), .Z(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n695), .A2(new_n696), .ZN(new_n699));
  NOR3_X1   g274(.A1(new_n694), .A2(new_n699), .A3(new_n697), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n694), .A2(new_n699), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n702));
  AOI211_X1 g277(.A(new_n698), .B(new_n700), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(new_n701), .B2(new_n702), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1991), .B(G1996), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT87), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n706), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1981), .B(G1986), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n709), .A2(new_n711), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(G229));
  XOR2_X1   g289(.A(KEYINPUT88), .B(G29), .Z(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n716), .A2(G35), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G162), .B2(new_n716), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT29), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G2090), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n715), .A2(G26), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT28), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n495), .A2(G128), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n492), .A2(G140), .ZN(new_n724));
  OR2_X1    g299(.A1(G104), .A2(G2105), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n725), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT93), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n723), .A2(new_n724), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G29), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n722), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G2067), .ZN(new_n732));
  INV_X1    g307(.A(G16), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G5), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G171), .B2(new_n733), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1961), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n557), .A2(new_n733), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n733), .B2(G19), .ZN(new_n738));
  INV_X1    g313(.A(G1341), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT31), .B(G11), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT96), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n743));
  AND3_X1   g318(.A1(new_n743), .A2(KEYINPUT97), .A3(G28), .ZN(new_n744));
  AOI21_X1  g319(.A(KEYINPUT97), .B1(new_n743), .B2(G28), .ZN(new_n745));
  OAI221_X1 g320(.A(new_n730), .B1(new_n743), .B2(G28), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n740), .A2(new_n742), .A3(new_n746), .ZN(new_n747));
  OAI22_X1  g322(.A1(new_n738), .A2(new_n739), .B1(new_n654), .B2(new_n715), .ZN(new_n748));
  NOR3_X1   g323(.A1(new_n736), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(G4), .A2(G16), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n634), .B2(G16), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G1348), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n492), .A2(G141), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n495), .A2(G129), .ZN(new_n755));
  NAND3_X1  g330(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT26), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n466), .A2(G105), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n754), .A2(new_n755), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(new_n730), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n730), .B2(G32), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT27), .B(G1996), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n752), .A2(new_n753), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n749), .A2(new_n766), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n730), .A2(G33), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n492), .A2(G139), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT25), .Z(new_n771));
  AOI22_X1  g346(.A1(new_n481), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n769), .B(new_n771), .C1(new_n473), .C2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT94), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n768), .B1(new_n774), .B2(G29), .ZN(new_n775));
  AOI211_X1 g350(.A(new_n732), .B(new_n767), .C1(new_n442), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n733), .A2(G21), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G168), .B2(new_n733), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1966), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n715), .A2(G27), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G164), .B2(new_n715), .ZN(new_n781));
  OAI22_X1  g356(.A1(new_n775), .A2(new_n442), .B1(G2078), .B2(new_n781), .ZN(new_n782));
  AOI211_X1 g357(.A(new_n779), .B(new_n782), .C1(G2078), .C2(new_n781), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n776), .A2(new_n783), .ZN(new_n784));
  OAI22_X1  g359(.A1(new_n752), .A2(new_n753), .B1(new_n764), .B2(new_n765), .ZN(new_n785));
  NAND2_X1  g360(.A1(G160), .A2(G29), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT24), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(G34), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(G34), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n715), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(G2084), .B1(new_n786), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n785), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n786), .A2(G2084), .A3(new_n790), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT95), .Z(new_n794));
  NAND2_X1  g369(.A1(new_n733), .A2(G20), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT23), .ZN(new_n796));
  INV_X1    g371(.A(G299), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n733), .ZN(new_n798));
  INV_X1    g373(.A(G1956), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n792), .A2(new_n794), .A3(new_n800), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n720), .A2(new_n784), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT92), .B(KEYINPUT36), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n492), .A2(G131), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT89), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n473), .A2(G107), .ZN(new_n807));
  OAI21_X1  g382(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n495), .A2(G119), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(new_n716), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G25), .B2(new_n716), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT35), .B(G1991), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n814), .A2(new_n815), .ZN(new_n818));
  MUX2_X1   g393(.A(G24), .B(G290), .S(G16), .Z(new_n819));
  INV_X1    g394(.A(G1986), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NOR3_X1   g397(.A1(new_n817), .A2(new_n818), .A3(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n609), .A2(G16), .ZN(new_n825));
  OR2_X1    g400(.A1(G6), .A2(G16), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(KEYINPUT90), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT90), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n825), .A2(new_n829), .A3(new_n826), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT32), .B(G1981), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n828), .A2(new_n832), .A3(new_n830), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n733), .A2(G23), .ZN(new_n836));
  INV_X1    g411(.A(G288), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n837), .B2(new_n733), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT33), .B(G1976), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n733), .A2(G22), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(G166), .B2(new_n733), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G1971), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n834), .A2(new_n835), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(KEYINPUT91), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT91), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n834), .A2(new_n847), .A3(new_n835), .A4(new_n844), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT34), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n824), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n846), .A2(KEYINPUT34), .A3(new_n848), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n804), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n851), .A2(new_n852), .A3(new_n804), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n803), .B1(new_n854), .B2(new_n855), .ZN(G311));
  INV_X1    g431(.A(new_n855), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n802), .B1(new_n857), .B2(new_n853), .ZN(G150));
  NAND2_X1  g433(.A1(new_n634), .A2(G559), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT38), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n861));
  INV_X1    g436(.A(G67), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(new_n517), .B2(new_n518), .ZN(new_n863));
  NAND2_X1  g438(.A1(G80), .A2(G543), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n861), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  OAI211_X1 g441(.A(KEYINPUT98), .B(new_n864), .C1(new_n542), .C2(new_n862), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(G651), .A3(new_n867), .ZN(new_n868));
  AOI22_X1  g443(.A1(G93), .A2(new_n544), .B1(new_n546), .B2(G55), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n557), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n557), .B1(new_n868), .B2(new_n869), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n860), .B(new_n872), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n873), .A2(KEYINPUT39), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(KEYINPUT39), .ZN(new_n875));
  NOR3_X1   g450(.A1(new_n874), .A2(new_n875), .A3(G860), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n868), .A2(new_n869), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(G860), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT37), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n876), .A2(new_n879), .ZN(G145));
  XNOR2_X1  g455(.A(G160), .B(new_n654), .ZN(new_n881));
  XNOR2_X1  g456(.A(G162), .B(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n774), .B(new_n761), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n811), .B(new_n647), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n505), .ZN(new_n886));
  AOI211_X1 g461(.A(KEYINPUT99), .B(new_n499), .C1(new_n500), .C2(KEYINPUT4), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT99), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n889));
  INV_X1    g464(.A(new_n499), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n886), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n729), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n492), .A2(G142), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n894), .B(KEYINPUT100), .Z(new_n895));
  NAND2_X1  g470(.A1(new_n495), .A2(G130), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n473), .A2(G118), .ZN(new_n897));
  OAI21_X1  g472(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n895), .B(new_n896), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n893), .B(new_n899), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n885), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n885), .A2(new_n900), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n882), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n885), .A2(new_n900), .ZN(new_n904));
  INV_X1    g479(.A(new_n882), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n885), .A2(new_n900), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g483(.A(KEYINPUT101), .B(G37), .Z(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g486(.A1(new_n870), .A2(new_n871), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n642), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n572), .A2(new_n573), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT74), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n572), .A2(new_n573), .A3(KEYINPUT74), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n918), .A2(new_n568), .A3(new_n627), .A4(new_n632), .ZN(new_n919));
  NAND2_X1  g494(.A1(G299), .A2(new_n633), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n913), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(KEYINPUT41), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT41), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n919), .A2(new_n920), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n922), .B1(new_n913), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT42), .ZN(new_n928));
  XNOR2_X1  g503(.A(G290), .B(KEYINPUT102), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n609), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n929), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(new_n606), .A3(new_n608), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(G303), .B(G288), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n930), .A2(new_n932), .A3(new_n934), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n928), .B(new_n938), .ZN(new_n939));
  MUX2_X1   g514(.A(new_n877), .B(new_n939), .S(G868), .Z(G295));
  MUX2_X1   g515(.A(new_n877), .B(new_n939), .S(G868), .Z(G331));
  XNOR2_X1  g516(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n527), .A2(new_n535), .A3(new_n536), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n944), .A2(new_n580), .B1(new_n541), .B2(new_n548), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n945), .B1(new_n582), .B2(G171), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT104), .B1(new_n946), .B2(new_n872), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n948));
  AOI21_X1  g523(.A(G301), .B1(new_n578), .B2(new_n581), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n912), .B(new_n948), .C1(new_n949), .C2(new_n945), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n582), .A2(G171), .ZN(new_n952));
  INV_X1    g527(.A(new_n945), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(new_n872), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT105), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT105), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n946), .A2(new_n956), .A3(new_n872), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n926), .B1(new_n951), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT106), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n926), .B(new_n961), .C1(new_n951), .C2(new_n958), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n946), .B(new_n872), .ZN(new_n963));
  OR2_X1    g538(.A1(new_n963), .A2(new_n921), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n960), .A2(new_n938), .A3(new_n962), .A4(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G37), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n962), .A2(new_n964), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n938), .B1(new_n968), .B2(new_n960), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n943), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT107), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n972), .B(new_n943), .C1(new_n967), .C2(new_n969), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n923), .A2(KEYINPUT108), .A3(new_n925), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n974), .B(new_n963), .C1(KEYINPUT108), .C2(new_n923), .ZN(new_n975));
  INV_X1    g550(.A(new_n958), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n947), .A2(new_n950), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n975), .B1(new_n921), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n938), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n981), .A2(new_n909), .A3(new_n965), .A4(new_n942), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n971), .A2(new_n973), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n960), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n962), .A2(new_n964), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n980), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n986), .A2(new_n966), .A3(new_n965), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n987), .A2(new_n943), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n981), .A2(new_n909), .A3(new_n965), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n988), .B1(KEYINPUT43), .B2(new_n989), .ZN(new_n990));
  MUX2_X1   g565(.A(new_n983), .B(new_n990), .S(KEYINPUT44), .Z(G397));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n889), .A2(new_n890), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT99), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n501), .A2(new_n888), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n505), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n992), .B1(new_n996), .B2(G1384), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n467), .A2(G40), .A3(new_n476), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n481), .A2(new_n479), .A3(G125), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT66), .B1(new_n483), .B2(new_n484), .ZN(new_n1001));
  AOI22_X1  g576(.A1(new_n1000), .A2(new_n1001), .B1(G113), .B2(G2104), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n999), .B1(new_n473), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n997), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(G290), .A2(G1986), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1004), .A2(KEYINPUT48), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G2067), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n728), .B(new_n1007), .ZN(new_n1008));
  OR2_X1    g583(.A1(new_n812), .A2(new_n815), .ZN(new_n1009));
  INV_X1    g584(.A(G1996), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n761), .B(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n812), .A2(new_n815), .ZN(new_n1012));
  AND4_X1   g587(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1004), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1006), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT48), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1008), .A2(new_n762), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT126), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n1004), .A2(new_n1018), .B1(new_n1019), .B2(KEYINPUT46), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(KEYINPUT46), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n1004), .A2(new_n1010), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1021), .B1(new_n1004), .B2(new_n1010), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g599(.A(new_n1024), .B(KEYINPUT47), .Z(new_n1025));
  NAND2_X1  g600(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1026));
  OAI22_X1  g601(.A1(new_n1012), .A2(new_n1026), .B1(G2067), .B2(new_n728), .ZN(new_n1027));
  AOI211_X1 g602(.A(new_n1017), .B(new_n1025), .C1(new_n1004), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1384), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n998), .B1(G2105), .B2(new_n486), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n892), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G8), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1981), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n594), .A2(new_n604), .A3(new_n1035), .ZN(new_n1036));
  XOR2_X1   g611(.A(KEYINPUT111), .B(G86), .Z(new_n1037));
  AOI21_X1  g612(.A(new_n603), .B1(new_n544), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1036), .B1(new_n1038), .B2(new_n1035), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT49), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1036), .B(KEYINPUT49), .C1(new_n1038), .C2(new_n1035), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(new_n1034), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1976), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1043), .A2(new_n1044), .A3(new_n837), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1036), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1034), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1031), .A2(G8), .A3(new_n1044), .A4(G288), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT110), .B1(new_n837), .B2(G1976), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1031), .A2(new_n1049), .A3(G8), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n1048), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1050), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1043), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(G166), .A2(new_n1033), .ZN(new_n1055));
  XNOR2_X1  g630(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1055), .B(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1029), .B1(new_n501), .B2(new_n505), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1003), .B1(KEYINPUT50), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n892), .A2(new_n1060), .A3(new_n1029), .ZN(new_n1061));
  INV_X1    g636(.A(G2090), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1003), .B1(new_n992), .B2(new_n1058), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n892), .A2(KEYINPUT45), .A3(new_n1029), .ZN(new_n1065));
  AOI21_X1  g640(.A(G1971), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g641(.A(G8), .B(new_n1057), .C1(new_n1063), .C2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1047), .B1(new_n1054), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1030), .B1(new_n1058), .B2(KEYINPUT50), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n994), .A2(new_n995), .ZN(new_n1071));
  AOI21_X1  g646(.A(G1384), .B1(new_n1071), .B2(new_n886), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1070), .B(KEYINPUT112), .C1(new_n1072), .C2(new_n1060), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT112), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1060), .B1(new_n892), .B2(new_n1029), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1074), .B1(new_n1075), .B2(new_n1069), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(new_n1076), .A3(new_n1062), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1066), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1057), .B1(new_n1079), .B2(G8), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1067), .B(new_n1043), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n997), .A2(new_n1084), .A3(new_n1030), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT45), .B1(new_n892), .B2(new_n1029), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT113), .B1(new_n1086), .B2(new_n1003), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1058), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT45), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1085), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G1966), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(G2084), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(G286), .A2(new_n1033), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1083), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1094), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1097), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1099), .A2(KEYINPUT114), .A3(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1082), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT63), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1105), .A2(new_n1033), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT63), .B1(new_n1106), .B2(new_n1057), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1107), .A2(new_n1081), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n1101), .B2(new_n1098), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1068), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1092), .A2(G168), .A3(new_n1095), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(G8), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1099), .A2(G168), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT51), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AOI211_X1 g689(.A(KEYINPUT51), .B(new_n1033), .C1(new_n1099), .C2(G168), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT51), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1033), .B1(new_n1099), .B2(G168), .ZN(new_n1120));
  INV_X1    g695(.A(G168), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1089), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n997), .A2(new_n1030), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1122), .B1(new_n1123), .B2(KEYINPUT113), .ZN(new_n1124));
  AOI21_X1  g699(.A(G1966), .B1(new_n1124), .B2(new_n1085), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1121), .B1(new_n1125), .B2(new_n1094), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1119), .B1(new_n1120), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT62), .B1(new_n1127), .B2(new_n1115), .ZN(new_n1128));
  AOI21_X1  g703(.A(G1961), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n443), .A2(KEYINPUT53), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1130), .B1(new_n1090), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1064), .A2(new_n1065), .A3(new_n443), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(G171), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1137), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1118), .A2(new_n1128), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1110), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1136), .A2(G171), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT121), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n473), .B1(new_n1002), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(new_n1143), .B2(new_n1002), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n997), .A2(new_n1142), .A3(new_n999), .A4(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n999), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT122), .B1(new_n1086), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1131), .B1(new_n1072), .B2(KEYINPUT45), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1146), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT123), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1146), .A2(new_n1148), .A3(new_n1152), .A4(new_n1149), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1141), .A2(new_n1151), .A3(new_n1153), .A4(new_n1130), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1154), .A2(KEYINPUT124), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(KEYINPUT124), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1155), .A2(new_n1156), .A3(new_n1137), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT54), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1157), .A2(KEYINPUT125), .A3(new_n1158), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1141), .B(new_n1130), .C1(new_n1131), .C2(new_n1090), .ZN(new_n1164));
  AND4_X1   g739(.A1(new_n1153), .A2(new_n1151), .A3(new_n1130), .A4(new_n1135), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1164), .B(KEYINPUT54), .C1(new_n1165), .C2(G301), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1166), .B(new_n1082), .C1(new_n1127), .C2(new_n1115), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT119), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n799), .B1(new_n1075), .B2(new_n1069), .ZN(new_n1169));
  XNOR2_X1  g744(.A(KEYINPUT56), .B(G2072), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1064), .A2(new_n1065), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT117), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT57), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n914), .A2(new_n1174), .A3(new_n568), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1175), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT117), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1169), .A2(new_n1178), .A3(new_n1171), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1173), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1169), .A2(new_n1176), .A3(new_n1171), .ZN(new_n1181));
  AND2_X1   g756(.A1(new_n1181), .A2(KEYINPUT61), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1184));
  OAI21_X1  g759(.A(KEYINPUT118), .B1(new_n1184), .B2(G1996), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT118), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1064), .A2(new_n1065), .A3(new_n1186), .A4(new_n1010), .ZN(new_n1187));
  XOR2_X1   g762(.A(KEYINPUT58), .B(G1341), .Z(new_n1188));
  NAND2_X1  g763(.A1(new_n1031), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1185), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT59), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1190), .A2(new_n1191), .A3(new_n557), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1192), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1191), .B1(new_n1190), .B2(new_n557), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1183), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1181), .A2(KEYINPUT115), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT115), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1169), .A2(new_n1197), .A3(new_n1171), .A4(new_n1176), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1172), .A2(new_n1177), .ZN(new_n1200));
  AOI21_X1  g775(.A(KEYINPUT61), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1168), .B1(new_n1195), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1201), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1194), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1192), .ZN(new_n1205));
  NAND4_X1  g780(.A1(new_n1203), .A2(new_n1205), .A3(KEYINPUT119), .A4(new_n1183), .ZN(new_n1206));
  AOI22_X1  g781(.A1(new_n1093), .A2(new_n753), .B1(new_n1032), .B2(new_n1007), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1207), .A2(KEYINPUT60), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1208), .B(new_n634), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1209), .B1(KEYINPUT60), .B2(new_n1207), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1202), .A2(new_n1206), .A3(new_n1210), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1207), .A2(new_n633), .ZN(new_n1212));
  XNOR2_X1  g787(.A(new_n1212), .B(KEYINPUT116), .ZN(new_n1213));
  INV_X1    g788(.A(new_n1180), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1199), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1167), .B1(new_n1211), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1140), .B1(new_n1163), .B2(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g792(.A(G290), .B(new_n820), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1014), .B1(new_n1013), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1028), .B1(new_n1217), .B2(new_n1219), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g795(.A1(G227), .A2(G401), .A3(new_n463), .ZN(new_n1222));
  NAND3_X1  g796(.A1(new_n712), .A2(new_n713), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g797(.A(new_n1223), .B1(new_n908), .B2(new_n909), .ZN(new_n1224));
  NAND2_X1  g798(.A1(new_n973), .A2(new_n982), .ZN(new_n1225));
  AOI21_X1  g799(.A(new_n972), .B1(new_n987), .B2(new_n943), .ZN(new_n1226));
  OAI211_X1 g800(.A(new_n1224), .B(KEYINPUT127), .C1(new_n1225), .C2(new_n1226), .ZN(new_n1227));
  INV_X1    g801(.A(new_n1227), .ZN(new_n1228));
  AOI21_X1  g802(.A(KEYINPUT127), .B1(new_n983), .B2(new_n1224), .ZN(new_n1229));
  NOR2_X1   g803(.A1(new_n1228), .A2(new_n1229), .ZN(G308));
  OAI21_X1  g804(.A(new_n1224), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1231));
  INV_X1    g805(.A(KEYINPUT127), .ZN(new_n1232));
  NAND2_X1  g806(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g807(.A1(new_n1233), .A2(new_n1227), .ZN(G225));
endmodule


