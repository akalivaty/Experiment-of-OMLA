//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n806,
    new_n807, new_n809, new_n810, new_n811, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932;
  INV_X1    g000(.A(KEYINPUT6), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(G120gat), .ZN(new_n205));
  INV_X1    g004(.A(G120gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(G113gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n203), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(G113gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n204), .A2(G120gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT69), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n208), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  AND2_X1   g012(.A1(G127gat), .A2(G134gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(G127gat), .A2(G134gat), .ZN(new_n215));
  NOR3_X1   g014(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT68), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n217));
  OR2_X1    g016(.A1(G127gat), .A2(G134gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(G127gat), .A2(G134gat), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n213), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n209), .B1(new_n214), .B2(new_n215), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G113gat), .B(G120gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT70), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT70), .B1(new_n205), .B2(new_n207), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n222), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G155gat), .ZN(new_n231));
  INV_X1    g030(.A(G162gat), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT2), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G141gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n234), .A2(G148gat), .ZN(new_n235));
  INV_X1    g034(.A(G148gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n236), .A2(G141gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n233), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT75), .B1(new_n235), .B2(new_n237), .ZN(new_n239));
  XNOR2_X1  g038(.A(G155gat), .B(G162gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n238), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(G141gat), .B(G148gat), .Z(new_n243));
  OAI211_X1 g042(.A(new_n243), .B(new_n233), .C1(KEYINPUT75), .C2(new_n240), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(KEYINPUT4), .B1(new_n230), .B2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n223), .B1(new_n226), .B2(new_n225), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n213), .A2(new_n221), .B1(new_n247), .B2(new_n228), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT4), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n242), .A2(new_n244), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT5), .ZN(new_n253));
  NAND2_X1  g052(.A1(G225gat), .A2(G233gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n245), .A2(KEYINPUT3), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n242), .A2(new_n244), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n230), .A3(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n252), .A2(new_n253), .A3(new_n254), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT77), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n250), .A2(new_n256), .B1(new_n229), .B2(new_n222), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n246), .A2(new_n251), .B1(new_n261), .B2(new_n255), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT77), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n262), .A2(new_n263), .A3(new_n253), .A4(new_n254), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n254), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n230), .A2(new_n245), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n250), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n254), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n253), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n260), .A2(new_n264), .B1(new_n265), .B2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(G57gat), .B(G85gat), .Z(new_n272));
  XNOR2_X1  g071(.A(G1gat), .B(G29gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n274), .B(new_n275), .Z(new_n276));
  OAI21_X1  g075(.A(new_n202), .B1(new_n271), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n264), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n265), .A2(new_n270), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n278), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT83), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n278), .A2(new_n279), .ZN(new_n282));
  INV_X1    g081(.A(new_n276), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT83), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n271), .A2(new_n276), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .A4(new_n202), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n282), .A2(KEYINPUT6), .A3(new_n283), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n281), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AND2_X1   g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290));
  INV_X1    g089(.A(G169gat), .ZN(new_n291));
  INV_X1    g090(.A(G176gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n290), .B1(new_n293), .B2(KEYINPUT26), .ZN(new_n294));
  NOR2_X1   g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT26), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT28), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(G190gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT27), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G183gat), .ZN(new_n304));
  INV_X1    g103(.A(G183gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT27), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n302), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT67), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT27), .B(G183gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n310), .A2(KEYINPUT67), .A3(new_n302), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT66), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G183gat), .ZN(new_n314));
  AOI21_X1  g113(.A(G190gat), .B1(new_n314), .B2(KEYINPUT27), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n303), .A3(G183gat), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT28), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n300), .B1(new_n312), .B2(new_n318), .ZN(new_n319));
  OR2_X1    g118(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n290), .B1(new_n320), .B2(new_n295), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT24), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n299), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G190gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n305), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  AND2_X1   g126(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n328));
  NOR2_X1   g127(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n293), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n321), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT25), .ZN(new_n332));
  OR3_X1    g131(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n333), .A2(new_n323), .A3(new_n326), .A4(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT25), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n335), .A2(new_n336), .A3(new_n330), .A4(new_n321), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n230), .B1(new_n319), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G227gat), .A2(G233gat), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n321), .A2(new_n336), .A3(new_n330), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n341), .A2(new_n335), .B1(new_n331), .B2(KEYINPUT25), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n294), .A2(new_n297), .B1(G183gat), .B2(G190gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n309), .A2(new_n311), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n343), .B1(new_n344), .B2(new_n317), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n248), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n339), .A2(new_n340), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT71), .B1(new_n347), .B2(KEYINPUT34), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT34), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n339), .A2(new_n350), .A3(new_n340), .A4(new_n346), .ZN(new_n351));
  OR2_X1    g150(.A1(new_n351), .A2(KEYINPUT72), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n347), .A2(KEYINPUT71), .A3(KEYINPUT34), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(KEYINPUT72), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n349), .A2(new_n352), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n340), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n248), .A2(new_n342), .A3(new_n345), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n342), .A2(new_n345), .B1(new_n229), .B2(new_n222), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT32), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT33), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G15gat), .B(G43gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(G71gat), .B(G99gat), .ZN(new_n364));
  XOR2_X1   g163(.A(new_n363), .B(new_n364), .Z(new_n365));
  NAND3_X1  g164(.A1(new_n360), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n365), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n359), .B(KEYINPUT32), .C1(new_n361), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n355), .A2(new_n369), .ZN(new_n370));
  XOR2_X1   g169(.A(G211gat), .B(G218gat), .Z(new_n371));
  XOR2_X1   g170(.A(G197gat), .B(G204gat), .Z(new_n372));
  AOI21_X1  g171(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G211gat), .B(G218gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(G197gat), .B(G204gat), .ZN(new_n376));
  INV_X1    g175(.A(G211gat), .ZN(new_n377));
  INV_X1    g176(.A(G218gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n375), .B(new_n376), .C1(KEYINPUT22), .C2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT29), .B1(new_n374), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n256), .B1(new_n381), .B2(KEYINPUT79), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n374), .A2(new_n380), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT29), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n383), .A2(KEYINPUT79), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n245), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G228gat), .A2(G233gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n257), .A2(new_n384), .ZN(new_n388));
  INV_X1    g187(.A(new_n383), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n245), .B1(new_n381), .B2(KEYINPUT3), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT78), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n388), .A2(new_n389), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT78), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n397), .B(new_n245), .C1(new_n381), .C2(KEYINPUT3), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n395), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n387), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n386), .A2(KEYINPUT80), .A3(new_n390), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n393), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  XOR2_X1   g201(.A(G78gat), .B(G106gat), .Z(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(G22gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT31), .B(G50gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n393), .A2(new_n400), .A3(new_n401), .A4(new_n406), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n347), .A2(KEYINPUT71), .A3(KEYINPUT34), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n411), .A2(new_n348), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT72), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n351), .B(new_n413), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n412), .A2(new_n414), .A3(new_n368), .A4(new_n366), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n370), .A2(new_n410), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(G226gat), .A2(G233gat), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n342), .A2(new_n345), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n418), .B1(new_n419), .B2(new_n384), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n417), .B1(new_n342), .B2(new_n345), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n389), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n419), .A2(new_n418), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT29), .B1(new_n342), .B2(new_n345), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n423), .B(new_n383), .C1(new_n418), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  XOR2_X1   g225(.A(G64gat), .B(G92gat), .Z(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(KEYINPUT74), .ZN(new_n428));
  XNOR2_X1  g227(.A(G8gat), .B(G36gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n422), .A2(new_n425), .A3(new_n430), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(KEYINPUT30), .A3(new_n433), .ZN(new_n434));
  OR3_X1    g233(.A1(new_n426), .A2(KEYINPUT30), .A3(new_n431), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NOR3_X1   g235(.A1(new_n416), .A2(new_n436), .A3(KEYINPUT35), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n289), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT87), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT87), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n289), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n416), .A2(KEYINPUT88), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT88), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n370), .A2(new_n410), .A3(new_n415), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n288), .B1(new_n277), .B2(new_n280), .ZN(new_n446));
  INV_X1    g245(.A(new_n436), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT35), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n439), .A2(new_n441), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n252), .A2(new_n258), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n269), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n266), .A2(new_n267), .A3(new_n254), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT39), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT81), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT81), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n453), .A2(new_n456), .A3(KEYINPUT39), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n452), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n458), .B(new_n276), .C1(KEYINPUT39), .C2(new_n452), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT40), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT82), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n459), .B(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(new_n284), .A3(new_n436), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT84), .B(KEYINPUT37), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT85), .B1(new_n426), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT85), .ZN(new_n466));
  INV_X1    g265(.A(new_n464), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n422), .A2(new_n425), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT38), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n430), .B1(new_n426), .B2(KEYINPUT37), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT86), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n469), .A2(new_n471), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT38), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n469), .A2(KEYINPUT86), .A3(new_n470), .A4(new_n471), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n474), .A2(new_n476), .A3(new_n477), .A4(new_n433), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n463), .B(new_n410), .C1(new_n478), .C2(new_n289), .ZN(new_n479));
  INV_X1    g278(.A(new_n370), .ZN(new_n480));
  INV_X1    g279(.A(new_n415), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  XOR2_X1   g281(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT36), .ZN(new_n485));
  OAI22_X1  g284(.A1(new_n480), .A2(new_n481), .B1(KEYINPUT73), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n410), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n484), .A2(new_n486), .B1(new_n448), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n479), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n450), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT89), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT89), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n450), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT14), .ZN(new_n495));
  NOR2_X1   g294(.A1(G29gat), .A2(G36gat), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT92), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT92), .B1(G29gat), .B2(G36gat), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n498), .B(new_n500), .ZN(new_n501));
  XOR2_X1   g300(.A(G43gat), .B(G50gat), .Z(new_n502));
  INV_X1    g301(.A(KEYINPUT15), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n502), .A2(new_n503), .B1(G29gat), .B2(G36gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n502), .A2(new_n503), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT94), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT17), .ZN(new_n509));
  INV_X1    g308(.A(new_n506), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n505), .B(new_n510), .ZN(new_n511));
  OR2_X1    g310(.A1(new_n508), .A2(KEYINPUT17), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n508), .A2(KEYINPUT17), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(G85gat), .A2(G92gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(KEYINPUT7), .ZN(new_n517));
  INV_X1    g316(.A(G99gat), .ZN(new_n518));
  INV_X1    g317(.A(G106gat), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT8), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n517), .B(new_n520), .C1(G85gat), .C2(G92gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(G99gat), .B(G106gat), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n521), .B(new_n522), .Z(new_n523));
  NAND2_X1  g322(.A1(new_n515), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT100), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT100), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n515), .A2(new_n526), .A3(new_n523), .ZN(new_n527));
  NAND2_X1  g326(.A1(G232gat), .A2(G233gat), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n528), .B(KEYINPUT99), .Z(new_n529));
  INV_X1    g328(.A(KEYINPUT41), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n521), .B(new_n522), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n531), .B1(new_n507), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n525), .A2(new_n527), .A3(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(G134gat), .B(G162gat), .Z(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n535), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n525), .A2(new_n537), .A3(new_n527), .A4(new_n533), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G190gat), .B(G218gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT101), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n529), .A2(new_n530), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n541), .B(new_n542), .Z(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n536), .A2(new_n543), .A3(new_n538), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(G8gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(G15gat), .B(G22gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT16), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n550), .B1(new_n551), .B2(G1gat), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT93), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n549), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n552), .B1(G1gat), .B2(new_n550), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(G57gat), .B(G64gat), .Z(new_n557));
  INV_X1    g356(.A(G71gat), .ZN(new_n558));
  INV_X1    g357(.A(G78gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n557), .B(KEYINPUT97), .C1(KEYINPUT9), .C2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G71gat), .B(G78gat), .Z(new_n562));
  OR2_X1    g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n562), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n565), .A2(KEYINPUT21), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(KEYINPUT21), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n556), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n568), .B1(new_n556), .B2(new_n566), .ZN(new_n569));
  XNOR2_X1  g368(.A(G183gat), .B(G211gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT98), .ZN(new_n571));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n569), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G127gat), .B(G155gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n574), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n580));
  XNOR2_X1  g379(.A(G113gat), .B(G141gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G169gat), .B(G197gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n584), .B(KEYINPUT12), .Z(new_n585));
  INV_X1    g384(.A(new_n556), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n511), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n587), .B1(new_n515), .B2(new_n586), .ZN(new_n588));
  NAND2_X1  g387(.A1(G229gat), .A2(G233gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(KEYINPUT95), .A2(KEYINPUT18), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n588), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  OR3_X1    g391(.A1(new_n507), .A2(KEYINPUT96), .A3(new_n556), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT96), .B1(new_n507), .B2(new_n556), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n593), .B(new_n594), .C1(new_n586), .C2(new_n511), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n589), .B(KEYINPUT13), .Z(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n591), .B1(new_n588), .B2(new_n589), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n585), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n585), .ZN(new_n603));
  OAI211_X1 g402(.A(KEYINPUT91), .B(new_n603), .C1(new_n598), .C2(new_n599), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G176gat), .B(G204gat), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT104), .ZN(new_n607));
  XNOR2_X1  g406(.A(G120gat), .B(G148gat), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n607), .B(new_n608), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G230gat), .A2(G233gat), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n563), .A2(new_n564), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n523), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n565), .A2(new_n532), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT10), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n565), .A2(KEYINPUT10), .A3(new_n532), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n612), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n610), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT105), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI211_X1 g422(.A(KEYINPUT105), .B(new_n610), .C1(new_n619), .C2(new_n620), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT103), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n609), .B1(new_n620), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n627), .B1(new_n626), .B2(new_n620), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n617), .A2(new_n618), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT102), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n612), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n617), .A2(new_n618), .A3(KEYINPUT102), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n625), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(KEYINPUT106), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT106), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n625), .A2(new_n637), .A3(new_n634), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NOR4_X1   g438(.A1(new_n548), .A2(new_n579), .A3(new_n605), .A4(new_n639), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n494), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n446), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(G1gat), .ZN(G1324gat));
  INV_X1    g443(.A(KEYINPUT42), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n641), .A2(new_n436), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT107), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT16), .B(G8gat), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n645), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n646), .A2(new_n645), .A3(new_n649), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n651), .B1(new_n648), .B2(G8gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(G1325gat));
  AOI21_X1  g452(.A(G15gat), .B1(new_n641), .B2(new_n482), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n486), .A2(G15gat), .A3(new_n484), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n654), .B1(new_n641), .B2(new_n655), .ZN(G1326gat));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n487), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT108), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT43), .B(G22gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(G1327gat));
  NOR3_X1   g459(.A1(new_n605), .A2(new_n639), .A3(new_n578), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n491), .A2(new_n493), .A3(new_n548), .A4(new_n661), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n662), .A2(G29gat), .A3(new_n446), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n663), .B(KEYINPUT45), .Z(new_n664));
  INV_X1    g463(.A(new_n661), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n491), .A2(new_n493), .A3(new_n548), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(KEYINPUT44), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n547), .B1(new_n450), .B2(new_n489), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n665), .B1(new_n667), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(G29gat), .B1(new_n673), .B2(new_n446), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n664), .A2(new_n674), .ZN(G1328gat));
  OAI21_X1  g474(.A(G36gat), .B1(new_n673), .B2(new_n447), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n447), .A2(G36gat), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT46), .B1(new_n662), .B2(new_n677), .ZN(new_n678));
  OR3_X1    g477(.A1(new_n662), .A2(KEYINPUT46), .A3(new_n677), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n676), .A2(new_n678), .A3(new_n679), .ZN(G1329gat));
  INV_X1    g479(.A(KEYINPUT109), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n484), .A2(new_n486), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n673), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(G43gat), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n662), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n686), .A2(new_n684), .A3(new_n482), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(new_n683), .B2(new_n684), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT47), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  OAI221_X1 g489(.A(new_n687), .B1(new_n681), .B2(KEYINPUT47), .C1(new_n683), .C2(new_n684), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(G1330gat));
  INV_X1    g491(.A(G50gat), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n693), .B1(new_n672), .B2(new_n487), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n494), .A2(KEYINPUT111), .A3(new_n548), .A4(new_n661), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT111), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n662), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n410), .A2(G50gat), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT112), .B1(new_n694), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT48), .B1(new_n701), .B2(KEYINPUT110), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT112), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n670), .B1(new_n666), .B2(KEYINPUT44), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n704), .A2(new_n410), .A3(new_n665), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n703), .B(new_n701), .C1(new_n705), .C2(new_n693), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n700), .A2(new_n702), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n702), .B1(new_n700), .B2(new_n706), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(G1331gat));
  NOR2_X1   g508(.A1(new_n548), .A2(new_n579), .ZN(new_n710));
  AND4_X1   g509(.A1(new_n490), .A2(new_n605), .A3(new_n710), .A4(new_n639), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n642), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n436), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n715));
  XOR2_X1   g514(.A(KEYINPUT49), .B(G64gat), .Z(new_n716));
  OAI21_X1  g515(.A(new_n715), .B1(new_n714), .B2(new_n716), .ZN(G1333gat));
  AOI21_X1  g516(.A(G71gat), .B1(new_n711), .B2(new_n482), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n682), .A2(new_n558), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n711), .B2(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g520(.A1(new_n711), .A2(new_n487), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT113), .B(G78gat), .Z(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1335gat));
  NAND2_X1  g523(.A1(new_n667), .A2(new_n671), .ZN(new_n725));
  INV_X1    g524(.A(new_n604), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n588), .A2(new_n589), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n590), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n728), .A2(new_n597), .A3(new_n592), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n603), .B1(new_n729), .B2(KEYINPUT91), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(new_n578), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n725), .A2(new_n639), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733), .B2(new_n446), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n668), .A2(new_n732), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT51), .Z(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n639), .ZN(new_n737));
  OR2_X1    g536(.A1(new_n446), .A2(G85gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n734), .B1(new_n737), .B2(new_n738), .ZN(G1336gat));
  OAI21_X1  g538(.A(G92gat), .B1(new_n733), .B2(new_n447), .ZN(new_n740));
  INV_X1    g539(.A(new_n639), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n741), .A2(G92gat), .A3(new_n447), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(KEYINPUT114), .Z(new_n743));
  NAND2_X1  g542(.A1(new_n736), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g545(.A(G99gat), .B1(new_n733), .B2(new_n682), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n639), .A2(new_n518), .A3(new_n482), .ZN(new_n748));
  XOR2_X1   g547(.A(new_n748), .B(KEYINPUT115), .Z(new_n749));
  NAND2_X1  g548(.A1(new_n736), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n750), .ZN(G1338gat));
  INV_X1    g550(.A(KEYINPUT116), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n733), .A2(new_n410), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n753), .B2(new_n519), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n736), .A2(new_n519), .A3(new_n487), .A4(new_n639), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(new_n753), .B2(new_n519), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n754), .A2(new_n756), .A3(KEYINPUT53), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n758));
  OAI221_X1 g557(.A(new_n755), .B1(new_n752), .B2(new_n758), .C1(new_n753), .C2(new_n519), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(G1339gat));
  NOR2_X1   g559(.A1(new_n588), .A2(new_n589), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT117), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n589), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n556), .B1(new_n509), .B2(new_n514), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n762), .B(new_n764), .C1(new_n765), .C2(new_n587), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n596), .B2(new_n595), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n584), .B1(new_n763), .B2(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n728), .A2(new_n597), .A3(new_n592), .A4(new_n603), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n639), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT54), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n609), .B1(new_n619), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n629), .A2(new_n630), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n775), .A2(new_n632), .A3(new_n611), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT54), .B1(new_n629), .B2(new_n611), .ZN(new_n777));
  OAI211_X1 g576(.A(KEYINPUT55), .B(new_n774), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n634), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AOI22_X1  g581(.A1(new_n772), .A2(KEYINPUT118), .B1(new_n731), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n639), .A2(new_n771), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n548), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n548), .A2(new_n771), .A3(new_n782), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n579), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n710), .A2(new_n605), .A3(new_n741), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n446), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n416), .A2(new_n436), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT119), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT119), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n791), .A2(new_n795), .A3(new_n792), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(G113gat), .B1(new_n797), .B2(new_n605), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n445), .A2(new_n436), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n791), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n801), .A2(new_n204), .A3(new_n731), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n798), .A2(new_n802), .ZN(G1340gat));
  NAND3_X1  g602(.A1(new_n801), .A2(new_n206), .A3(new_n639), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n794), .A2(new_n639), .A3(new_n796), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n805), .A2(KEYINPUT120), .A3(G120gat), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT120), .B1(new_n805), .B2(G120gat), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n804), .B1(new_n806), .B2(new_n807), .ZN(G1341gat));
  INV_X1    g607(.A(G127gat), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n797), .A2(new_n809), .A3(new_n579), .ZN(new_n810));
  AOI21_X1  g609(.A(G127gat), .B1(new_n801), .B2(new_n578), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n810), .A2(new_n811), .ZN(G1342gat));
  NOR3_X1   g611(.A1(new_n800), .A2(G134gat), .A3(new_n547), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT56), .ZN(new_n814));
  OAI21_X1  g613(.A(G134gat), .B1(new_n797), .B2(new_n547), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(G1343gat));
  AND2_X1   g615(.A1(new_n778), .A2(new_n634), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n777), .B1(new_n632), .B2(new_n631), .ZN(new_n818));
  INV_X1    g617(.A(new_n774), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n780), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n602), .A2(new_n817), .A3(new_n604), .A4(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n770), .B1(new_n636), .B2(new_n638), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n821), .B1(new_n822), .B2(new_n784), .ZN(new_n823));
  INV_X1    g622(.A(new_n785), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n547), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n578), .B1(new_n825), .B2(new_n787), .ZN(new_n826));
  INV_X1    g625(.A(new_n790), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n487), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n820), .A2(KEYINPUT121), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT121), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n781), .A2(new_n831), .A3(new_n780), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n817), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n605), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n547), .B1(new_n834), .B2(new_n822), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n578), .B1(new_n835), .B2(new_n787), .ZN(new_n836));
  OAI211_X1 g635(.A(KEYINPUT57), .B(new_n487), .C1(new_n836), .C2(new_n827), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT122), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n828), .A2(new_n829), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n831), .B1(new_n781), .B2(new_n780), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n779), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n731), .A2(new_n832), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n548), .B1(new_n842), .B2(new_n772), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n579), .B1(new_n843), .B2(new_n788), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n410), .B1(new_n844), .B2(new_n790), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n845), .A2(KEYINPUT122), .A3(KEYINPUT57), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n839), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n682), .A2(new_n642), .A3(new_n447), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n847), .A2(new_n731), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(G141gat), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n828), .A2(new_n848), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n234), .A3(new_n731), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n851), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n848), .B1(new_n839), .B2(new_n846), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n234), .B1(new_n856), .B2(new_n731), .ZN(new_n857));
  INV_X1    g656(.A(new_n854), .ZN(new_n858));
  OAI21_X1  g657(.A(KEYINPUT58), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n855), .A2(new_n859), .ZN(G1344gat));
  NAND3_X1  g659(.A1(new_n853), .A2(new_n236), .A3(new_n639), .ZN(new_n861));
  AOI211_X1 g660(.A(KEYINPUT59), .B(new_n236), .C1(new_n856), .C2(new_n639), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863));
  AOI211_X1 g662(.A(KEYINPUT57), .B(new_n410), .C1(new_n844), .C2(new_n790), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n864), .B1(KEYINPUT57), .B2(new_n828), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n639), .A3(new_n849), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n863), .B1(new_n866), .B2(G148gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n861), .B1(new_n862), .B2(new_n867), .ZN(G1345gat));
  AOI21_X1  g667(.A(G155gat), .B1(new_n853), .B2(new_n578), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n578), .A2(G155gat), .ZN(new_n870));
  XOR2_X1   g669(.A(new_n870), .B(KEYINPUT123), .Z(new_n871));
  AOI21_X1  g670(.A(new_n869), .B1(new_n856), .B2(new_n871), .ZN(G1346gat));
  AOI21_X1  g671(.A(G162gat), .B1(new_n853), .B2(new_n548), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n547), .A2(new_n232), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n856), .B2(new_n874), .ZN(G1347gat));
  NAND2_X1  g674(.A1(new_n789), .A2(new_n790), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n642), .A2(new_n447), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n416), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(G169gat), .B1(new_n880), .B2(new_n605), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n878), .A2(new_n445), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n291), .A3(new_n731), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(KEYINPUT124), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT124), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n881), .A2(new_n886), .A3(new_n883), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(G1348gat));
  AOI21_X1  g687(.A(G176gat), .B1(new_n882), .B2(new_n639), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n741), .A2(new_n292), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n879), .B2(new_n890), .ZN(G1349gat));
  OAI21_X1  g690(.A(G183gat), .B1(new_n880), .B2(new_n579), .ZN(new_n892));
  OR2_X1    g691(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n578), .A2(new_n310), .ZN(new_n894));
  AOI22_X1  g693(.A1(new_n882), .A2(new_n894), .B1(KEYINPUT125), .B2(KEYINPUT60), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n893), .B1(new_n892), .B2(new_n895), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(G1350gat));
  NAND3_X1  g697(.A1(new_n882), .A2(new_n324), .A3(new_n548), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n879), .A2(new_n548), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(G190gat), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n901), .A2(KEYINPUT61), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(KEYINPUT61), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(G1351gat));
  NAND2_X1  g703(.A1(new_n682), .A2(new_n877), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n828), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(G197gat), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n907), .A3(new_n731), .ZN(new_n908));
  INV_X1    g707(.A(new_n905), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n865), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(KEYINPUT126), .A3(new_n731), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(G197gat), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT126), .B1(new_n910), .B2(new_n731), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n908), .B1(new_n912), .B2(new_n913), .ZN(G1352gat));
  NOR4_X1   g713(.A1(new_n828), .A2(G204gat), .A3(new_n741), .A4(new_n905), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT62), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n865), .A2(new_n639), .A3(new_n909), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G204gat), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1353gat));
  NAND3_X1  g718(.A1(new_n906), .A2(new_n377), .A3(new_n578), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n828), .A2(KEYINPUT57), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n845), .A2(new_n829), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n921), .A2(new_n578), .A3(new_n922), .A4(new_n909), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(KEYINPUT127), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT127), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n865), .A2(new_n925), .A3(new_n578), .A4(new_n909), .ZN(new_n926));
  AND4_X1   g725(.A1(KEYINPUT63), .A2(new_n924), .A3(G211gat), .A4(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n377), .B1(new_n923), .B2(KEYINPUT127), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT63), .B1(new_n928), .B2(new_n926), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n920), .B1(new_n927), .B2(new_n929), .ZN(G1354gat));
  AOI21_X1  g729(.A(G218gat), .B1(new_n906), .B2(new_n548), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n547), .A2(new_n378), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(new_n910), .B2(new_n932), .ZN(G1355gat));
endmodule


