//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n786, new_n788, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G141gat), .B(G148gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(KEYINPUT2), .ZN(new_n208));
  INV_X1    g007(.A(G141gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(G148gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT73), .B(G141gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n210), .B1(new_n211), .B2(G148gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n204), .B1(new_n213), .B2(new_n205), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n208), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G134gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G127gat), .ZN(new_n217));
  INV_X1    g016(.A(G127gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G134gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G113gat), .B(G120gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(KEYINPUT1), .ZN(new_n222));
  INV_X1    g021(.A(G120gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G113gat), .ZN(new_n224));
  INV_X1    g023(.A(G113gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G120gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G127gat), .B(G134gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n222), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT75), .B1(new_n215), .B2(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n222), .A2(new_n230), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n209), .A2(KEYINPUT73), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT73), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G141gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n236), .A3(G148gat), .ZN(new_n237));
  INV_X1    g036(.A(G148gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G141gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n205), .A2(new_n213), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n203), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n238), .A2(G141gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n213), .B1(new_n210), .B2(new_n243), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n240), .A2(new_n242), .B1(new_n244), .B2(new_n206), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT75), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n233), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT4), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n232), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(G225gat), .A2(G233gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT74), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n237), .A2(new_n239), .B1(new_n203), .B2(new_n241), .ZN(new_n253));
  XNOR2_X1  g052(.A(G155gat), .B(G162gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n209), .A2(G148gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n254), .B1(new_n213), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT3), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n208), .B(new_n259), .C1(new_n212), .C2(new_n214), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n260), .A3(new_n231), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n215), .A2(new_n231), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT4), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n249), .A2(new_n252), .A3(new_n261), .A4(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n215), .A2(new_n231), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n232), .A2(new_n247), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT76), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n266), .A2(new_n267), .A3(new_n251), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n267), .B1(new_n266), .B2(new_n251), .ZN(new_n269));
  OAI211_X1 g068(.A(KEYINPUT5), .B(new_n264), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n232), .A2(new_n247), .A3(KEYINPUT4), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT78), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n272), .B1(new_n262), .B2(new_n248), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n232), .A2(new_n247), .A3(new_n272), .A4(KEYINPUT4), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n261), .A2(new_n276), .A3(new_n252), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n274), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n270), .A2(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(G1gat), .B(G29gat), .Z(new_n280));
  XNOR2_X1  g079(.A(G57gat), .B(G85gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n202), .B1(new_n279), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n284), .ZN(new_n286));
  AOI211_X1 g085(.A(KEYINPUT83), .B(new_n286), .C1(new_n270), .C2(new_n278), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT82), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n274), .A2(new_n261), .A3(new_n275), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT39), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n291), .A3(new_n251), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(new_n286), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT39), .B1(new_n266), .B2(new_n251), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n294), .B1(new_n290), .B2(new_n251), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n289), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT40), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT40), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n289), .B(new_n298), .C1(new_n293), .C2(new_n295), .ZN(new_n299));
  INV_X1    g098(.A(G226gat), .ZN(new_n300));
  INV_X1    g099(.A(G233gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(KEYINPUT29), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT25), .ZN(new_n305));
  OR2_X1    g104(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n306));
  INV_X1    g105(.A(G176gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n306), .A2(KEYINPUT23), .A3(new_n307), .A4(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT24), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G183gat), .ZN(new_n313));
  INV_X1    g112(.A(G190gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n312), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(G169gat), .A2(G176gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT23), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n309), .A2(new_n317), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n318), .B1(KEYINPUT23), .B2(new_n320), .ZN(new_n324));
  INV_X1    g123(.A(G169gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n325), .A2(new_n307), .A3(KEYINPUT23), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT25), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(G183gat), .A2(G190gat), .ZN(new_n329));
  AND2_X1   g128(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n329), .B1(new_n330), .B2(G190gat), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT65), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n310), .A2(new_n332), .A3(new_n311), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n332), .B1(new_n310), .B2(new_n311), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n331), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n305), .A2(new_n323), .B1(new_n328), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT27), .B(G183gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n338), .A3(new_n314), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n313), .A2(KEYINPUT27), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT27), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G183gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n342), .A3(new_n314), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT28), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n344), .A2(KEYINPUT66), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT26), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n318), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n348), .B1(new_n318), .B2(new_n349), .ZN(new_n350));
  AND4_X1   g149(.A1(new_n310), .A2(new_n339), .A3(new_n346), .A4(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n304), .B1(new_n336), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G211gat), .B(G218gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT70), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(G211gat), .ZN(new_n356));
  INV_X1    g155(.A(G218gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G211gat), .A2(G218gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(KEYINPUT70), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n355), .A2(KEYINPUT69), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G197gat), .ZN(new_n362));
  INV_X1    g161(.A(G204gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(G197gat), .A2(G204gat), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT22), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n364), .A2(new_n365), .B1(new_n366), .B2(new_n359), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n361), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n367), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n369), .A2(new_n355), .A3(KEYINPUT69), .A4(new_n360), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n323), .A2(new_n305), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n328), .A2(new_n335), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n339), .A2(new_n346), .A3(new_n310), .A4(new_n350), .ZN(new_n375));
  INV_X1    g174(.A(new_n302), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n352), .A2(new_n371), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n371), .B1(new_n352), .B2(new_n377), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(G8gat), .B(G36gat), .Z(new_n381));
  XNOR2_X1  g180(.A(G64gat), .B(G92gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT30), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT71), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n378), .B2(new_n379), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n352), .A2(new_n377), .ZN(new_n389));
  INV_X1    g188(.A(new_n371), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n352), .A2(new_n377), .A3(new_n371), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(KEYINPUT71), .A3(new_n392), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n383), .B(KEYINPUT72), .Z(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n388), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n380), .A2(KEYINPUT30), .A3(new_n383), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n386), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n288), .A2(new_n297), .A3(new_n299), .A4(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G78gat), .B(G106gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(G22gat), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(G228gat), .A2(G233gat), .ZN(new_n403));
  XOR2_X1   g202(.A(new_n403), .B(KEYINPUT80), .Z(new_n404));
  INV_X1    g203(.A(KEYINPUT29), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n371), .B1(new_n405), .B2(new_n260), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n355), .A2(new_n360), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n369), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n355), .A2(new_n360), .A3(new_n367), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n405), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n245), .B1(new_n410), .B2(new_n259), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n404), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT29), .B1(new_n368), .B2(new_n370), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n215), .B1(new_n413), .B2(KEYINPUT3), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n260), .A2(new_n405), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n390), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n403), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n414), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  XOR2_X1   g217(.A(KEYINPUT31), .B(G50gat), .Z(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n412), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n420), .B1(new_n412), .B2(new_n418), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n402), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n414), .A2(new_n416), .A3(new_n417), .ZN(new_n424));
  INV_X1    g223(.A(new_n404), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n259), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n215), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n425), .B1(new_n427), .B2(new_n416), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n419), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n418), .A3(new_n420), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n401), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n423), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n278), .ZN(new_n434));
  INV_X1    g233(.A(new_n269), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n266), .A2(new_n267), .A3(new_n251), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n264), .A2(KEYINPUT5), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n434), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT83), .B1(new_n439), .B2(new_n286), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n442), .B1(new_n439), .B2(new_n286), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n286), .B1(new_n270), .B2(new_n278), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n202), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n440), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n279), .A2(new_n284), .A3(new_n442), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OR3_X1    g247(.A1(new_n391), .A2(KEYINPUT84), .A3(new_n371), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n380), .A2(KEYINPUT84), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(new_n450), .A3(KEYINPUT37), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT37), .ZN(new_n452));
  AOI211_X1 g251(.A(KEYINPUT38), .B(new_n394), .C1(new_n380), .C2(new_n452), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n451), .A2(new_n453), .B1(new_n383), .B2(new_n380), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT85), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n388), .A2(new_n393), .A3(KEYINPUT37), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n383), .B1(new_n380), .B2(new_n452), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n455), .B1(new_n458), .B2(KEYINPUT38), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT38), .ZN(new_n460));
  AOI211_X1 g259(.A(KEYINPUT85), .B(new_n460), .C1(new_n456), .C2(new_n457), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n454), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n399), .B(new_n433), .C1(new_n448), .C2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT36), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT67), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n465), .B1(new_n336), .B2(new_n351), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n374), .A2(KEYINPUT67), .A3(new_n375), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n467), .A3(new_n231), .ZN(new_n468));
  INV_X1    g267(.A(G227gat), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n469), .A2(new_n301), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n465), .B(new_n233), .C1(new_n336), .C2(new_n351), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT33), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(G71gat), .B(G99gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(KEYINPUT68), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(G15gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(G43gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n468), .A2(new_n471), .ZN(new_n481));
  INV_X1    g280(.A(new_n470), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT34), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT34), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n481), .A2(new_n485), .A3(new_n482), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n480), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT32), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n478), .B1(new_n472), .B2(new_n473), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n485), .B1(new_n481), .B2(new_n482), .ZN(new_n491));
  AOI211_X1 g290(.A(KEYINPUT34), .B(new_n470), .C1(new_n468), .C2(new_n471), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n487), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n489), .B1(new_n487), .B2(new_n493), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n464), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n493), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n488), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n487), .A2(new_n489), .A3(new_n493), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(KEYINPUT36), .A3(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n268), .A2(new_n269), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n264), .A2(KEYINPUT5), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n278), .B(new_n286), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n441), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n447), .B1(new_n505), .B2(new_n444), .ZN(new_n506));
  INV_X1    g305(.A(new_n398), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n423), .A2(new_n431), .A3(KEYINPUT81), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT81), .B1(new_n423), .B2(new_n431), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n496), .A2(new_n501), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n494), .A2(new_n495), .A3(new_n398), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n432), .A2(KEYINPUT35), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n448), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n433), .A3(new_n500), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT35), .B1(new_n516), .B2(new_n508), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n463), .A2(new_n512), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G229gat), .A2(G233gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT13), .ZN(new_n520));
  XNOR2_X1  g319(.A(G15gat), .B(G22gat), .ZN(new_n521));
  INV_X1    g320(.A(G1gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT16), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(G1gat), .B2(new_n521), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(G8gat), .ZN(new_n526));
  INV_X1    g325(.A(G8gat), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n524), .B(new_n527), .C1(G1gat), .C2(new_n521), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G29gat), .ZN(new_n530));
  INV_X1    g329(.A(G36gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(new_n531), .A3(KEYINPUT14), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT14), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(G29gat), .B2(G36gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(G29gat), .A2(G36gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT15), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n532), .A2(new_n534), .A3(KEYINPUT15), .A4(new_n535), .ZN(new_n539));
  XNOR2_X1  g338(.A(G43gat), .B(G50gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n539), .A2(new_n540), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n529), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n526), .A2(new_n528), .A3(new_n541), .A4(new_n542), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n520), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n529), .A2(new_n543), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(KEYINPUT17), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT17), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n541), .A2(new_n549), .A3(new_n542), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n529), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n547), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(new_n519), .ZN(new_n554));
  XNOR2_X1  g353(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n546), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT87), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n553), .A2(new_n557), .A3(KEYINPUT18), .A4(new_n519), .ZN(new_n558));
  INV_X1    g357(.A(new_n550), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n549), .B1(new_n541), .B2(new_n542), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n552), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n561), .A2(KEYINPUT18), .A3(new_n519), .A4(new_n544), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT87), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G113gat), .B(G141gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(G197gat), .ZN(new_n566));
  XOR2_X1   g365(.A(KEYINPUT11), .B(G169gat), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT12), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n556), .A2(new_n564), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n569), .B1(new_n556), .B2(new_n564), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n518), .A2(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(G155gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(G183gat), .B(G211gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G71gat), .A2(G78gat), .ZN(new_n580));
  OR2_X1    g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(G57gat), .B(G64gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT9), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n580), .B(new_n581), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(new_n580), .ZN(new_n585));
  INV_X1    g384(.A(G57gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(G64gat), .ZN(new_n587));
  INV_X1    g386(.A(G64gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(G57gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n580), .A2(new_n583), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n585), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n584), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT88), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n584), .A2(KEYINPUT88), .A3(new_n592), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n529), .B1(new_n598), .B2(KEYINPUT21), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT21), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(G231gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n603), .A2(new_n301), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n597), .B(new_n601), .C1(new_n603), .C2(new_n301), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n218), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n605), .A2(new_n218), .A3(new_n606), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n600), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n605), .A2(new_n218), .A3(new_n606), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n611), .A2(new_n607), .A3(new_n599), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n579), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n608), .A2(new_n600), .A3(new_n609), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n599), .B1(new_n611), .B2(new_n607), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(new_n615), .A3(new_n578), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G85gat), .A2(G92gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT7), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(KEYINPUT89), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT90), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n621), .B1(new_n618), .B2(KEYINPUT7), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT7), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n623), .A2(KEYINPUT90), .A3(G85gat), .A4(G92gat), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT89), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n618), .A2(new_n625), .A3(KEYINPUT7), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n620), .A2(new_n622), .A3(new_n624), .A4(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(G99gat), .B(G106gat), .Z(new_n628));
  NAND2_X1  g427(.A1(G99gat), .A2(G106gat), .ZN(new_n629));
  INV_X1    g428(.A(G85gat), .ZN(new_n630));
  INV_X1    g429(.A(G92gat), .ZN(new_n631));
  AOI22_X1  g430(.A1(KEYINPUT8), .A2(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n627), .A2(new_n628), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n628), .B1(new_n627), .B2(new_n632), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  AND2_X1   g435(.A1(G232gat), .A2(G233gat), .ZN(new_n637));
  AOI22_X1  g436(.A1(new_n636), .A2(new_n543), .B1(KEYINPUT41), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n551), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n638), .B1(new_n639), .B2(new_n636), .ZN(new_n640));
  XOR2_X1   g439(.A(G190gat), .B(G218gat), .Z(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n641), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n638), .B(new_n643), .C1(new_n639), .C2(new_n636), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n637), .A2(KEYINPUT41), .ZN(new_n646));
  XNOR2_X1  g445(.A(G134gat), .B(G162gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n642), .A2(new_n648), .A3(new_n644), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n617), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n628), .A2(KEYINPUT91), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n654), .B1(new_n627), .B2(new_n632), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(new_n593), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n627), .A2(new_n632), .A3(new_n654), .ZN(new_n657));
  AOI22_X1  g456(.A1(new_n635), .A2(new_n597), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT10), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n597), .A2(new_n659), .ZN(new_n660));
  AOI22_X1  g459(.A1(new_n658), .A2(new_n659), .B1(new_n660), .B2(new_n636), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT92), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n635), .A2(new_n597), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n656), .A2(new_n657), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n664), .A2(new_n659), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n660), .A2(new_n636), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT92), .ZN(new_n669));
  NAND2_X1  g468(.A1(G230gat), .A2(G233gat), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n663), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n658), .A2(new_n670), .ZN(new_n672));
  XNOR2_X1  g471(.A(G120gat), .B(G148gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(G176gat), .B(G204gat), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n673), .B(new_n674), .Z(new_n675));
  AND2_X1   g474(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n670), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n672), .B1(new_n661), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n675), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n653), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n506), .A2(KEYINPUT93), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n506), .A2(KEYINPUT93), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n574), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT94), .B(G1gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1324gat));
  NAND2_X1  g488(.A1(new_n574), .A2(new_n683), .ZN(new_n690));
  OAI21_X1  g489(.A(KEYINPUT95), .B1(new_n690), .B2(new_n507), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n463), .A2(new_n512), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n515), .A2(new_n517), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n572), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n570), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n694), .A2(new_n696), .A3(new_n683), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT95), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n697), .A2(new_n698), .A3(new_n398), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n691), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT16), .B(G8gat), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(KEYINPUT96), .Z(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OR4_X1    g504(.A1(new_n704), .A2(new_n690), .A3(new_n507), .A4(new_n701), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n691), .A2(G8gat), .A3(new_n699), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT97), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n705), .B(new_n706), .C1(new_n709), .C2(new_n710), .ZN(G1325gat));
  NOR2_X1   g510(.A1(new_n494), .A2(new_n495), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  OR3_X1    g512(.A1(new_n690), .A2(G15gat), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n496), .A2(new_n501), .ZN(new_n715));
  OAI21_X1  g514(.A(G15gat), .B1(new_n690), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(G1326gat));
  NAND3_X1  g516(.A1(new_n574), .A2(new_n511), .A3(new_n683), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT43), .B(G22gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1327gat));
  AND3_X1   g519(.A1(new_n642), .A2(new_n648), .A3(new_n644), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n648), .B1(new_n642), .B2(new_n644), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n694), .A2(KEYINPUT44), .A3(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(new_n518), .B2(new_n652), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n617), .B(KEYINPUT98), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n682), .B(KEYINPUT99), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n729), .A2(new_n730), .A3(new_n573), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n727), .A2(new_n686), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n530), .B1(new_n732), .B2(KEYINPUT100), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(KEYINPUT100), .B2(new_n732), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n617), .A2(new_n652), .A3(new_n682), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n574), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n736), .A2(new_n530), .A3(new_n686), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT45), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n734), .A2(new_n738), .ZN(G1328gat));
  INV_X1    g538(.A(KEYINPUT46), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n507), .A2(G36gat), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n736), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT102), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n727), .A2(new_n398), .A3(new_n731), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G36gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n736), .A2(new_n741), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT46), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n748), .A2(KEYINPUT101), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n748), .A2(KEYINPUT101), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n744), .B(new_n746), .C1(new_n749), .C2(new_n750), .ZN(G1329gat));
  INV_X1    g550(.A(KEYINPUT103), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT47), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n715), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n724), .A2(new_n726), .A3(new_n755), .A4(new_n731), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(G43gat), .ZN(new_n757));
  INV_X1    g556(.A(G43gat), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n736), .A2(new_n758), .A3(new_n712), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n754), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT103), .A2(KEYINPUT47), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(G1330gat));
  NAND3_X1  g561(.A1(new_n727), .A2(new_n432), .A3(new_n731), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n763), .A2(G50gat), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n574), .A2(new_n735), .ZN(new_n765));
  INV_X1    g564(.A(new_n511), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n765), .A2(G50gat), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT48), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n727), .A2(new_n511), .A3(new_n731), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n767), .B1(new_n770), .B2(G50gat), .ZN(new_n771));
  OAI22_X1  g570(.A1(new_n764), .A2(new_n769), .B1(new_n771), .B2(KEYINPUT48), .ZN(G1331gat));
  AOI21_X1  g571(.A(new_n723), .B1(new_n616), .B2(new_n613), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n730), .A2(new_n573), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT104), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n694), .ZN(new_n776));
  INV_X1    g575(.A(new_n686), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(new_n586), .ZN(G1332gat));
  AOI211_X1 g578(.A(new_n507), .B(new_n776), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n780));
  NOR2_X1   g579(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n780), .B(new_n781), .ZN(G1333gat));
  NOR3_X1   g581(.A1(new_n776), .A2(new_n713), .A3(G71gat), .ZN(new_n783));
  INV_X1    g582(.A(new_n776), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n755), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n783), .B1(G71gat), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g586(.A1(new_n776), .A2(new_n766), .ZN(new_n788));
  XNOR2_X1  g587(.A(KEYINPUT105), .B(G78gat), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(G1335gat));
  INV_X1    g589(.A(new_n682), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n696), .A2(new_n617), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n724), .A2(new_n726), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT106), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n724), .A2(new_n726), .A3(KEYINPUT106), .A4(new_n792), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n795), .A2(new_n686), .A3(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n696), .A2(new_n617), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n694), .A2(new_n723), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n694), .A2(KEYINPUT51), .A3(new_n723), .A4(new_n798), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n686), .A2(new_n630), .A3(new_n682), .ZN(new_n806));
  OAI22_X1  g605(.A1(new_n797), .A2(new_n630), .B1(new_n805), .B2(new_n806), .ZN(G1336gat));
  INV_X1    g606(.A(new_n730), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n507), .A2(G92gat), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI211_X1 g609(.A(new_n808), .B(new_n810), .C1(new_n801), .C2(new_n803), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n813), .B(G92gat), .C1(new_n793), .C2(new_n507), .ZN(new_n814));
  NAND2_X1  g613(.A1(KEYINPUT107), .A2(KEYINPUT52), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n795), .A2(new_n398), .A3(new_n796), .ZN(new_n817));
  AOI22_X1  g616(.A1(new_n817), .A2(G92gat), .B1(new_n811), .B2(KEYINPUT107), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n816), .B1(new_n818), .B2(new_n813), .ZN(G1337gat));
  NAND3_X1  g618(.A1(new_n795), .A2(new_n755), .A3(new_n796), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(G99gat), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n713), .A2(G99gat), .A3(new_n791), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(KEYINPUT108), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n821), .B1(new_n823), .B2(new_n805), .ZN(G1338gat));
  NOR2_X1   g623(.A1(new_n433), .A2(G106gat), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  AOI211_X1 g625(.A(new_n808), .B(new_n826), .C1(new_n801), .C2(new_n803), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(G106gat), .B1(new_n793), .B2(new_n433), .ZN(new_n829));
  XOR2_X1   g628(.A(KEYINPUT109), .B(KEYINPUT53), .Z(new_n830));
  NAND3_X1  g629(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n795), .A2(new_n511), .A3(new_n796), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n827), .B1(new_n832), .B2(G106gat), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n831), .B1(new_n833), .B2(new_n834), .ZN(G1339gat));
  INV_X1    g634(.A(KEYINPUT110), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n617), .A2(new_n695), .A3(new_n570), .A4(new_n652), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(new_n682), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n773), .A2(KEYINPUT110), .A3(new_n573), .A4(new_n791), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n544), .A2(new_n545), .A3(new_n520), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT113), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n841), .B(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT112), .B1(new_n553), .B2(new_n519), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n561), .A2(new_n544), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT112), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n845), .A2(new_n846), .A3(G229gat), .A4(G233gat), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n843), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n568), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n682), .A2(new_n570), .A3(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT111), .ZN(new_n851));
  AOI211_X1 g650(.A(KEYINPUT54), .B(new_n678), .C1(new_n666), .C2(new_n667), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n852), .B2(new_n675), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n668), .A2(new_n854), .A3(new_n670), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(KEYINPUT111), .A3(new_n680), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n854), .B1(new_n661), .B2(new_n678), .ZN(new_n857));
  AOI22_X1  g656(.A1(new_n853), .A2(new_n856), .B1(new_n671), .B2(new_n857), .ZN(new_n858));
  OAI22_X1  g657(.A1(new_n858), .A2(KEYINPUT55), .B1(new_n571), .B2(new_n572), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n670), .B1(new_n661), .B2(new_n662), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n668), .A2(KEYINPUT92), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n857), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n852), .A2(new_n851), .A3(new_n675), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT111), .B1(new_n855), .B2(new_n680), .ZN(new_n864));
  OAI211_X1 g663(.A(KEYINPUT55), .B(new_n862), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n677), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n850), .B1(new_n859), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n723), .B1(new_n858), .B2(KEYINPUT55), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n868), .A2(new_n866), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n849), .A2(new_n570), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n849), .A2(new_n570), .A3(KEYINPUT114), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI22_X1  g673(.A1(new_n867), .A2(new_n652), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n840), .B1(new_n875), .B2(new_n729), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n686), .A2(new_n513), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n432), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(G113gat), .B1(new_n880), .B2(new_n696), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n876), .A2(new_n766), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n877), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n573), .A2(new_n225), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n881), .B1(new_n886), .B2(new_n887), .ZN(G1340gat));
  AOI21_X1  g687(.A(G120gat), .B1(new_n880), .B2(new_n682), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n808), .A2(new_n223), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n886), .B2(new_n890), .ZN(G1341gat));
  OAI21_X1  g690(.A(G127gat), .B1(new_n885), .B2(new_n728), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n880), .A2(new_n218), .A3(new_n617), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1342gat));
  NOR3_X1   g693(.A1(new_n879), .A2(G134gat), .A3(new_n652), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT56), .ZN(new_n896));
  OAI21_X1  g695(.A(G134gat), .B1(new_n885), .B2(new_n652), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1343gat));
  NOR3_X1   g697(.A1(new_n777), .A2(new_n755), .A3(new_n398), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT57), .B1(new_n876), .B2(new_n432), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n511), .A2(KEYINPUT57), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT55), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n904), .A2(new_n696), .A3(new_n677), .A4(new_n865), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n723), .B1(new_n905), .B2(new_n850), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n872), .A2(new_n873), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n907), .A2(new_n866), .A3(new_n868), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n616), .B(new_n613), .C1(new_n906), .C2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n901), .B1(new_n909), .B2(new_n840), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n696), .B(new_n899), .C1(new_n900), .C2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT116), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n211), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n867), .A2(new_n652), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n869), .A2(new_n874), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n617), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n838), .A2(new_n839), .ZN(new_n918));
  OAI211_X1 g717(.A(KEYINPUT57), .B(new_n511), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n728), .B1(new_n906), .B2(new_n908), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n433), .B1(new_n920), .B2(new_n840), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n919), .B1(new_n921), .B2(KEYINPUT57), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n922), .A2(KEYINPUT116), .A3(new_n696), .A4(new_n899), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n913), .A2(new_n914), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n876), .A2(new_n432), .ZN(new_n925));
  INV_X1    g724(.A(new_n899), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n573), .A2(G141gat), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT58), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n911), .A2(new_n914), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n921), .A2(new_n899), .A3(new_n928), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT115), .ZN(new_n933));
  OAI21_X1  g732(.A(KEYINPUT58), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n930), .A2(new_n934), .ZN(G1344gat));
  NAND3_X1  g734(.A1(new_n927), .A2(new_n238), .A3(new_n682), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT57), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n925), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n926), .B1(new_n938), .B2(new_n919), .ZN(new_n939));
  AOI211_X1 g738(.A(KEYINPUT59), .B(new_n238), .C1(new_n939), .C2(new_n682), .ZN(new_n940));
  XOR2_X1   g739(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n941));
  NAND2_X1  g740(.A1(new_n925), .A2(KEYINPUT57), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n837), .A2(new_n682), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT118), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n937), .B(new_n511), .C1(new_n944), .C2(new_n917), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n942), .A2(new_n682), .A3(new_n899), .A4(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n941), .B1(new_n946), .B2(G148gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n936), .B1(new_n940), .B2(new_n947), .ZN(G1345gat));
  AOI21_X1  g747(.A(G155gat), .B1(new_n927), .B2(new_n617), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n729), .A2(G155gat), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT119), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n949), .B1(new_n939), .B2(new_n951), .ZN(G1346gat));
  NOR4_X1   g751(.A1(new_n925), .A2(G162gat), .A3(new_n926), .A4(new_n652), .ZN(new_n953));
  XOR2_X1   g752(.A(new_n953), .B(KEYINPUT120), .Z(new_n954));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n723), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(G162gat), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1347gat));
  NOR2_X1   g756(.A1(new_n516), .A2(new_n507), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n876), .A2(new_n777), .A3(new_n958), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n959), .A2(new_n306), .A3(new_n308), .A4(new_n696), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n686), .A2(new_n507), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(new_n712), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n882), .A2(new_n573), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n960), .B1(new_n325), .B2(new_n963), .ZN(G1348gat));
  NAND3_X1  g763(.A1(new_n959), .A2(new_n307), .A3(new_n682), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n882), .A2(new_n808), .A3(new_n962), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n965), .B1(new_n307), .B2(new_n966), .ZN(G1349gat));
  INV_X1    g766(.A(new_n962), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n883), .A2(new_n729), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(G183gat), .ZN(new_n970));
  NOR2_X1   g769(.A1(KEYINPUT121), .A2(KEYINPUT60), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n617), .A2(new_n337), .ZN(new_n973));
  AOI22_X1  g772(.A1(new_n959), .A2(new_n973), .B1(KEYINPUT121), .B2(KEYINPUT60), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n970), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n972), .B1(new_n970), .B2(new_n974), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n975), .A2(new_n976), .ZN(G1350gat));
  NAND3_X1  g776(.A1(new_n959), .A2(new_n314), .A3(new_n723), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n876), .A2(new_n968), .A3(new_n766), .A4(new_n723), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT61), .ZN(new_n980));
  AND4_X1   g779(.A1(KEYINPUT122), .A2(new_n979), .A3(new_n980), .A4(G190gat), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT122), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n314), .B1(new_n982), .B2(KEYINPUT61), .ZN(new_n983));
  AOI22_X1  g782(.A1(new_n979), .A2(new_n983), .B1(KEYINPUT122), .B2(new_n980), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n978), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(KEYINPUT123), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT123), .ZN(new_n987));
  OAI211_X1 g786(.A(new_n987), .B(new_n978), .C1(new_n981), .C2(new_n984), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n986), .A2(new_n988), .ZN(G1351gat));
  NAND2_X1  g788(.A1(new_n961), .A2(new_n715), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n990), .B(KEYINPUT124), .ZN(new_n991));
  NAND4_X1  g790(.A1(new_n942), .A2(new_n991), .A3(new_n696), .A4(new_n945), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n362), .B1(new_n992), .B2(KEYINPUT125), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n993), .B1(KEYINPUT125), .B2(new_n992), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n686), .B1(new_n920), .B2(new_n840), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n755), .A2(new_n507), .A3(new_n433), .ZN(new_n996));
  NAND4_X1  g795(.A1(new_n995), .A2(new_n362), .A3(new_n696), .A4(new_n996), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n994), .A2(new_n997), .ZN(G1352gat));
  NAND2_X1  g797(.A1(new_n995), .A2(new_n996), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n682), .A2(new_n363), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT126), .ZN(new_n1001));
  OAI22_X1  g800(.A1(new_n999), .A2(new_n1000), .B1(new_n1001), .B2(KEYINPUT62), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1001), .A2(KEYINPUT62), .ZN(new_n1003));
  OR2_X1    g802(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n942), .A2(new_n945), .A3(new_n991), .ZN(new_n1005));
  OAI21_X1  g804(.A(G204gat), .B1(new_n1005), .B2(new_n808), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n1004), .A2(new_n1006), .A3(new_n1007), .ZN(G1353gat));
  NAND2_X1  g807(.A1(new_n942), .A2(new_n945), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n961), .A2(new_n715), .A3(new_n617), .ZN(new_n1010));
  OAI21_X1  g809(.A(G211gat), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OR2_X1    g810(.A1(new_n1011), .A2(KEYINPUT63), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1011), .A2(KEYINPUT63), .ZN(new_n1013));
  NAND4_X1  g812(.A1(new_n995), .A2(new_n356), .A3(new_n617), .A4(new_n996), .ZN(new_n1014));
  XOR2_X1   g813(.A(new_n1014), .B(KEYINPUT127), .Z(new_n1015));
  NAND3_X1  g814(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .ZN(G1354gat));
  OAI21_X1  g815(.A(G218gat), .B1(new_n1005), .B2(new_n652), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n723), .A2(new_n357), .ZN(new_n1018));
  OAI21_X1  g817(.A(new_n1017), .B1(new_n999), .B2(new_n1018), .ZN(G1355gat));
endmodule


