//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027, new_n1028;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n202));
  XNOR2_X1  g001(.A(G1gat), .B(G29gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT0), .ZN(new_n204));
  XNOR2_X1  g003(.A(G57gat), .B(G85gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT5), .ZN(new_n208));
  OR2_X1    g007(.A1(KEYINPUT73), .A2(G148gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(KEYINPUT73), .A2(G148gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(G141gat), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G141gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G148gat), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215));
  INV_X1    g014(.A(G155gat), .ZN(new_n216));
  INV_X1    g015(.A(G162gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G148gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G141gat), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT2), .B1(new_n213), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n216), .A2(new_n217), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(new_n219), .ZN(new_n225));
  OAI22_X1  g024(.A1(new_n214), .A2(new_n220), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G113gat), .B(G120gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  XNOR2_X1  g027(.A(G127gat), .B(G134gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n229), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(KEYINPUT1), .B2(new_n227), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n211), .A2(new_n213), .B1(new_n219), .B2(new_n218), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n213), .A2(new_n222), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n225), .B1(new_n236), .B2(new_n215), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(new_n230), .A3(new_n232), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G225gat), .A2(G233gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n208), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n238), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(KEYINPUT3), .B1(new_n235), .B2(new_n237), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n246), .A3(new_n233), .ZN(new_n247));
  INV_X1    g046(.A(new_n233), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n248), .A2(new_n238), .A3(KEYINPUT4), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT74), .B(KEYINPUT4), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n250), .B1(new_n226), .B2(new_n233), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n247), .A2(new_n249), .A3(new_n241), .A4(new_n251), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n243), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n250), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n248), .A2(new_n238), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n239), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n255), .B(new_n208), .C1(new_n256), .C2(KEYINPUT4), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n247), .A2(new_n241), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI211_X1 g058(.A(KEYINPUT6), .B(new_n207), .C1(new_n253), .C2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n207), .B1(new_n253), .B2(new_n259), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT6), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n243), .A2(new_n252), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n263), .B(new_n206), .C1(new_n258), .C2(new_n257), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n261), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G8gat), .B(G36gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(G64gat), .B(G92gat), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n266), .B(new_n267), .Z(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G197gat), .B(G204gat), .ZN(new_n270));
  INV_X1    g069(.A(G211gat), .ZN(new_n271));
  INV_X1    g070(.A(G218gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT71), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G218gat), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n271), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT70), .B(KEYINPUT22), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n270), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G211gat), .B(G218gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n279), .B(new_n270), .C1(new_n276), .C2(new_n277), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G183gat), .ZN(new_n286));
  INV_X1    g085(.A(G190gat), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT24), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT24), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n289), .A2(G183gat), .A3(G190gat), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n288), .A2(new_n290), .B1(new_n286), .B2(new_n287), .ZN(new_n291));
  INV_X1    g090(.A(G169gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT23), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT25), .B1(new_n293), .B2(G176gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n295), .B1(KEYINPUT23), .B2(new_n296), .ZN(new_n297));
  NOR3_X1   g096(.A1(new_n291), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  AND2_X1   g097(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n293), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT66), .B1(new_n301), .B2(new_n297), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n303), .A2(G169gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT65), .ZN(new_n305));
  INV_X1    g104(.A(G176gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n304), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n296), .A2(KEYINPUT23), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n292), .A2(new_n306), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT66), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n309), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NOR3_X1   g115(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n288), .A2(new_n290), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n302), .A2(new_n314), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT25), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n298), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G226gat), .A2(G233gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT26), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT68), .B1(new_n295), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT68), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n327), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n296), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n330), .B1(new_n325), .B2(new_n295), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n329), .A2(new_n331), .B1(G183gat), .B2(G190gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n286), .A2(KEYINPUT27), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT27), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(G183gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n335), .A3(new_n287), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT28), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT27), .B(G183gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n339), .A2(KEYINPUT28), .A3(new_n287), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n332), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n323), .A2(new_n324), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n309), .A2(new_n312), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n345), .A2(KEYINPUT66), .B1(new_n318), .B2(new_n319), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT25), .B1(new_n346), .B2(new_n314), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT67), .B1(new_n347), .B2(new_n298), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n342), .A2(KEYINPUT69), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT69), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n332), .A2(new_n350), .A3(new_n341), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n321), .A2(new_n322), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT67), .ZN(new_n354));
  INV_X1    g153(.A(new_n298), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n348), .A2(new_n352), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n324), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(KEYINPUT29), .ZN(new_n359));
  AOI211_X1 g158(.A(new_n285), .B(new_n344), .C1(new_n357), .C2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n283), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n348), .A2(new_n356), .A3(new_n358), .A4(new_n352), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n359), .B1(new_n323), .B2(new_n343), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n269), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n362), .A2(new_n363), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n283), .ZN(new_n367));
  INV_X1    g166(.A(new_n351), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n350), .B1(new_n332), .B2(new_n341), .ZN(new_n369));
  OAI22_X1  g168(.A1(new_n323), .A2(new_n354), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n347), .A2(KEYINPUT67), .A3(new_n298), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n359), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n344), .ZN(new_n373));
  INV_X1    g172(.A(new_n285), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n367), .A2(new_n375), .A3(new_n268), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n365), .A2(KEYINPUT30), .A3(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n360), .A2(new_n364), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT30), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(new_n379), .A3(new_n268), .ZN(new_n380));
  AOI221_X4 g179(.A(new_n202), .B1(new_n260), .B2(new_n265), .C1(new_n377), .C2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n377), .A2(new_n380), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n265), .A2(new_n260), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT75), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G78gat), .B(G106gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(KEYINPUT77), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G228gat), .A2(G233gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT29), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT3), .B1(new_n283), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT29), .B1(new_n238), .B2(new_n244), .ZN(new_n393));
  OAI221_X1 g192(.A(new_n390), .B1(new_n238), .B2(new_n392), .C1(new_n285), .C2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n283), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT78), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n281), .A2(new_n396), .A3(new_n282), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n391), .B1(new_n281), .B2(new_n396), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT79), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  XOR2_X1   g198(.A(KEYINPUT70), .B(KEYINPUT22), .Z(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT71), .B(G218gat), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n400), .B1(new_n271), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n279), .B1(new_n402), .B2(new_n270), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT29), .B1(new_n403), .B2(KEYINPUT78), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT79), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n281), .A2(new_n396), .A3(new_n282), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n399), .A2(new_n244), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n395), .B1(new_n408), .B2(new_n226), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n394), .B1(new_n409), .B2(new_n390), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(G22gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT76), .B(KEYINPUT31), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(G50gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(G22gat), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n415), .B(new_n394), .C1(new_n409), .C2(new_n390), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n411), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n414), .B1(new_n411), .B2(new_n416), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n388), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n411), .A2(new_n416), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n413), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n411), .A2(new_n414), .A3(new_n416), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n387), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n385), .A2(new_n424), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n419), .A2(new_n423), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n265), .A2(new_n376), .A3(new_n260), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n367), .A2(new_n375), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n269), .B1(new_n428), .B2(KEYINPUT37), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n344), .B1(new_n357), .B2(new_n359), .ZN(new_n431));
  OAI22_X1  g230(.A1(new_n431), .A2(new_n374), .B1(new_n366), .B2(new_n283), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT38), .B1(new_n432), .B2(KEYINPUT37), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n427), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n428), .A2(KEYINPUT37), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT38), .B1(new_n435), .B2(new_n429), .ZN(new_n436));
  INV_X1    g235(.A(new_n382), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n247), .B(new_n255), .C1(new_n256), .C2(KEYINPUT4), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n242), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n240), .A2(new_n242), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT39), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n438), .A2(new_n441), .A3(new_n242), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n206), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT40), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n261), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n446), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT80), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT80), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n445), .A2(new_n450), .A3(new_n446), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n447), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n434), .A2(new_n436), .B1(new_n437), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT36), .ZN(new_n454));
  XOR2_X1   g253(.A(G15gat), .B(G43gat), .Z(new_n455));
  XNOR2_X1  g254(.A(G71gat), .B(G99gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n455), .B(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n357), .A2(new_n233), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n348), .A2(new_n356), .A3(new_n248), .A4(new_n352), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(G227gat), .A2(G233gat), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT33), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n458), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n459), .A2(new_n462), .A3(new_n460), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT34), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT34), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n459), .A2(new_n469), .A3(new_n462), .A4(new_n460), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n464), .A2(KEYINPUT32), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n462), .B1(new_n459), .B2(new_n460), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n457), .B1(new_n475), .B2(KEYINPUT33), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n476), .A2(new_n468), .A3(new_n470), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n472), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n474), .B1(new_n472), .B2(new_n477), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n454), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n472), .A2(new_n477), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n473), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n483), .A2(KEYINPUT36), .A3(new_n478), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n426), .A2(new_n453), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n419), .A2(new_n423), .A3(new_n483), .A4(new_n478), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT35), .B1(new_n486), .B2(new_n385), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n479), .A2(new_n480), .ZN(new_n488));
  INV_X1    g287(.A(new_n383), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n437), .A2(KEYINPUT35), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n426), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n425), .A2(new_n485), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G15gat), .B(G22gat), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT16), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n493), .B1(new_n494), .B2(G1gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(KEYINPUT84), .A2(G8gat), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n495), .B(new_n496), .C1(G1gat), .C2(new_n493), .ZN(new_n497));
  NOR2_X1   g296(.A1(KEYINPUT84), .A2(G8gat), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n498), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G43gat), .B(G50gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT15), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT81), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n502), .A2(KEYINPUT15), .ZN(new_n506));
  INV_X1    g305(.A(G29gat), .ZN(new_n507));
  INV_X1    g306(.A(G36gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT14), .ZN(new_n509));
  NAND2_X1  g308(.A1(G29gat), .A2(G36gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT14), .B1(new_n507), .B2(new_n508), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n502), .A2(KEYINPUT81), .A3(KEYINPUT15), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n505), .A2(new_n506), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n513), .A2(new_n503), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT17), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT83), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT82), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n515), .A2(new_n516), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n521), .B1(new_n515), .B2(new_n516), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n520), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n515), .A2(new_n516), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT82), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n515), .A2(new_n516), .A3(new_n521), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n528), .A2(new_n520), .A3(new_n525), .A4(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n519), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n528), .A2(new_n529), .A3(new_n500), .A4(new_n499), .ZN(new_n533));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n532), .A2(KEYINPUT18), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT18), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n528), .A2(new_n525), .A3(new_n529), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT83), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n518), .B1(new_n540), .B2(new_n530), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n538), .B1(new_n541), .B2(new_n535), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n501), .B1(new_n522), .B2(new_n523), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n533), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n534), .B(KEYINPUT13), .Z(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n537), .A2(new_n542), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT85), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n537), .A2(new_n548), .A3(new_n546), .ZN(new_n549));
  XNOR2_X1  g348(.A(G113gat), .B(G141gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(G197gat), .ZN(new_n551));
  XOR2_X1   g350(.A(KEYINPUT11), .B(G169gat), .Z(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT12), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n547), .A2(new_n549), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n546), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n530), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n535), .B1(new_n558), .B2(new_n519), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n557), .B1(new_n559), .B2(KEYINPUT18), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n560), .B(new_n542), .C1(new_n548), .C2(new_n554), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n492), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT92), .ZN(new_n564));
  XNOR2_X1  g363(.A(G120gat), .B(G148gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(G176gat), .B(G204gat), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n565), .B(new_n566), .Z(new_n567));
  INV_X1    g366(.A(G57gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(G64gat), .ZN(new_n569));
  INV_X1    g368(.A(G64gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(G57gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G71gat), .A2(G78gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT87), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT86), .ZN(new_n578));
  NOR2_X1   g377(.A1(G71gat), .A2(G78gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n578), .B1(new_n580), .B2(new_n573), .ZN(new_n581));
  INV_X1    g380(.A(new_n573), .ZN(new_n582));
  NOR3_X1   g381(.A1(new_n582), .A2(new_n579), .A3(KEYINPUT86), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n576), .B(new_n577), .C1(new_n581), .C2(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n582), .A2(new_n579), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT87), .B1(new_n576), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n580), .A2(new_n578), .A3(new_n573), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT86), .B1(new_n582), .B2(new_n579), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n587), .A2(new_n588), .B1(new_n572), .B2(new_n575), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n584), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(G85gat), .ZN(new_n591));
  INV_X1    g390(.A(G92gat), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT7), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT7), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(G85gat), .A3(G92gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G99gat), .B(G106gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(G99gat), .A2(G106gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n598), .B1(new_n591), .B2(new_n592), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n597), .B1(new_n596), .B2(new_n599), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n590), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n596), .A2(new_n599), .ZN(new_n605));
  INV_X1    g404(.A(new_n597), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(new_n600), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n576), .B1(new_n581), .B2(new_n583), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n569), .A2(new_n571), .B1(new_n574), .B2(new_n573), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n580), .A2(new_n573), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n577), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n608), .A2(new_n613), .A3(new_n584), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n604), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G230gat), .A2(G233gat), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n604), .A2(new_n614), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n590), .A2(new_n603), .A3(KEYINPUT10), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n616), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n567), .B1(new_n618), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n616), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n625), .B1(new_n620), .B2(new_n621), .ZN(new_n626));
  INV_X1    g425(.A(new_n567), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n617), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n564), .B1(new_n624), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n618), .A2(new_n623), .A3(new_n567), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n627), .B1(new_n617), .B2(new_n626), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n631), .A3(KEYINPUT92), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n590), .A2(KEYINPUT21), .ZN(new_n635));
  AND2_X1   g434(.A1(G231gat), .A2(G233gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(G127gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n590), .A2(KEYINPUT21), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n501), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n638), .A2(new_n641), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT88), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(G155gat), .ZN(new_n646));
  XOR2_X1   g445(.A(G183gat), .B(G211gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n642), .A2(new_n643), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n648), .B1(new_n642), .B2(new_n643), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n522), .A2(new_n523), .A3(new_n608), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT89), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT41), .ZN(new_n655));
  INV_X1    g454(.A(G232gat), .ZN(new_n656));
  INV_X1    g455(.A(G233gat), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  OR3_X1    g457(.A1(new_n653), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n654), .B1(new_n653), .B2(new_n658), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n558), .A2(new_n517), .A3(new_n608), .ZN(new_n662));
  XOR2_X1   g461(.A(G190gat), .B(G218gat), .Z(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n661), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n664), .B1(new_n661), .B2(new_n662), .ZN(new_n666));
  XNOR2_X1  g465(.A(G134gat), .B(G162gat), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n667), .B(new_n668), .Z(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  OAI22_X1  g469(.A1(new_n665), .A2(new_n666), .B1(KEYINPUT90), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n661), .A2(new_n662), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n663), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n661), .A2(new_n662), .A3(new_n664), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n669), .B(KEYINPUT90), .Z(new_n675));
  NAND3_X1  g474(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT91), .B1(new_n652), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n677), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT91), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n651), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n563), .A2(new_n634), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n383), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT93), .B(G1gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1324gat));
  NOR2_X1   g485(.A1(new_n683), .A2(new_n382), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n688), .A2(G8gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT16), .B(G8gat), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT42), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(KEYINPUT42), .B2(new_n691), .ZN(G1325gat));
  NAND2_X1  g492(.A1(new_n481), .A2(new_n484), .ZN(new_n694));
  OAI21_X1  g493(.A(G15gat), .B1(new_n683), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n488), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n696), .A2(G15gat), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n683), .B2(new_n697), .ZN(G1326gat));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n426), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT94), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT43), .B(G22gat), .Z(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1327gat));
  NAND3_X1  g501(.A1(new_n652), .A2(new_n634), .A3(new_n677), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT95), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n563), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n706), .A2(new_n507), .A3(new_n489), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT45), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n487), .A2(new_n491), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n426), .A2(new_n453), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(new_n425), .A3(new_n694), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n679), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT97), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT97), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n715), .B(KEYINPUT44), .C1(new_n492), .C2(new_n679), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT99), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n709), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT98), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n425), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n385), .A2(KEYINPUT98), .A3(new_n424), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(new_n485), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n487), .A2(KEYINPUT99), .A3(new_n491), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n719), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n725), .A2(new_n713), .A3(new_n677), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n717), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n633), .B(KEYINPUT96), .Z(new_n728));
  NOR3_X1   g527(.A1(new_n728), .A2(new_n651), .A3(new_n562), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(G29gat), .B1(new_n730), .B2(new_n383), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n708), .A2(new_n731), .ZN(G1328gat));
  NOR3_X1   g531(.A1(new_n705), .A2(G36gat), .A3(new_n382), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT46), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n730), .A2(new_n382), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n735), .A2(KEYINPUT100), .ZN(new_n736));
  OAI21_X1  g535(.A(G36gat), .B1(new_n735), .B2(KEYINPUT100), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(G1329gat));
  NOR3_X1   g537(.A1(new_n705), .A2(G43gat), .A3(new_n696), .ZN(new_n739));
  INV_X1    g538(.A(new_n694), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n727), .A2(new_n740), .A3(new_n729), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n739), .B1(new_n741), .B2(G43gat), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT101), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1330gat));
  OAI21_X1  g545(.A(G50gat), .B1(new_n730), .B2(new_n426), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT48), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n426), .A2(G50gat), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT102), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n706), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT104), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n748), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n747), .B(new_n754), .C1(new_n753), .C2(new_n752), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n751), .A2(KEYINPUT103), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n751), .A2(KEYINPUT103), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n747), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n755), .B1(new_n758), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g558(.A1(new_n682), .A2(new_n562), .A3(new_n728), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT105), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n725), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(new_n383), .ZN(new_n763));
  XNOR2_X1  g562(.A(KEYINPUT106), .B(G57gat), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(G1332gat));
  NOR2_X1   g564(.A1(new_n762), .A2(new_n382), .ZN(new_n766));
  NOR2_X1   g565(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n767));
  AND2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n766), .B2(new_n767), .ZN(G1333gat));
  OAI21_X1  g569(.A(G71gat), .B1(new_n762), .B2(new_n694), .ZN(new_n771));
  OR2_X1    g570(.A1(new_n696), .A2(G71gat), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n762), .B2(new_n772), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n773), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g573(.A1(new_n762), .A2(new_n426), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n775), .B(G78gat), .Z(G1335gat));
  NAND2_X1  g575(.A1(new_n556), .A2(new_n561), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n651), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n633), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT107), .B1(new_n727), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT107), .ZN(new_n782));
  AOI211_X1 g581(.A(new_n782), .B(new_n779), .C1(new_n717), .C2(new_n726), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n591), .B1(new_n784), .B2(new_n489), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n634), .A2(G85gat), .A3(new_n383), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n725), .A2(new_n677), .A3(new_n778), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n725), .A2(KEYINPUT51), .A3(new_n677), .A4(new_n778), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n789), .A2(KEYINPUT108), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT108), .B1(new_n789), .B2(new_n790), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n786), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT109), .B1(new_n785), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n781), .A2(new_n783), .A3(new_n383), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n796), .B(new_n793), .C1(new_n797), .C2(new_n591), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n798), .ZN(G1336gat));
  NAND2_X1  g598(.A1(new_n789), .A2(new_n790), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n728), .ZN(new_n802));
  NOR4_X1   g601(.A1(new_n801), .A2(G92gat), .A3(new_n382), .A4(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n727), .A2(new_n780), .ZN(new_n805));
  OAI21_X1  g604(.A(G92gat), .B1(new_n805), .B2(new_n382), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n804), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n784), .A2(new_n437), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n803), .B1(new_n809), .B2(G92gat), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n808), .B1(new_n810), .B2(new_n807), .ZN(G1337gat));
  INV_X1    g610(.A(G99gat), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n488), .A2(new_n812), .A3(new_n633), .ZN(new_n813));
  XOR2_X1   g612(.A(new_n813), .B(KEYINPUT110), .Z(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n791), .B2(new_n792), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n781), .A2(new_n783), .A3(new_n694), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n815), .B1(new_n816), .B2(new_n812), .ZN(G1338gat));
  OAI21_X1  g616(.A(G106gat), .B1(new_n805), .B2(new_n426), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n802), .A2(new_n426), .A3(G106gat), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT53), .B1(new_n800), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  XOR2_X1   g620(.A(new_n819), .B(KEYINPUT111), .Z(new_n822));
  NOR2_X1   g621(.A1(new_n801), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n784), .A2(new_n424), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n823), .B1(new_n824), .B2(G106gat), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n821), .B1(new_n825), .B2(new_n826), .ZN(G1339gat));
  NAND4_X1  g626(.A1(new_n678), .A2(new_n562), .A3(new_n634), .A4(new_n681), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n567), .B1(new_n626), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n620), .A2(new_n621), .A3(new_n625), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n623), .A2(KEYINPUT54), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT112), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n626), .A2(new_n830), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT112), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n836), .A2(new_n837), .A3(new_n833), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n832), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n630), .B1(new_n839), .B2(KEYINPUT55), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841));
  AOI211_X1 g640(.A(new_n841), .B(new_n832), .C1(new_n835), .C2(new_n838), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n534), .B1(new_n532), .B2(new_n533), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n544), .A2(new_n545), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n553), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n537), .A2(new_n542), .A3(new_n546), .A4(new_n554), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n843), .A2(new_n677), .A3(new_n848), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n633), .A2(new_n846), .A3(new_n847), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n850), .B1(new_n843), .B2(new_n777), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n679), .B1(new_n851), .B2(KEYINPUT113), .ZN(new_n852));
  INV_X1    g651(.A(new_n850), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n834), .A2(KEYINPUT112), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n837), .B1(new_n836), .B2(new_n833), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n831), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n841), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n839), .A2(KEYINPUT55), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n630), .A3(new_n858), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n853), .B(KEYINPUT113), .C1(new_n562), .C2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n849), .B1(new_n852), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n651), .B1(new_n862), .B2(KEYINPUT114), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT114), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n864), .B(new_n849), .C1(new_n852), .C2(new_n861), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n829), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n424), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n437), .A2(new_n383), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n488), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(G113gat), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n869), .A2(new_n870), .A3(new_n562), .ZN(new_n871));
  NOR4_X1   g670(.A1(new_n866), .A2(new_n383), .A3(new_n437), .A4(new_n486), .ZN(new_n872));
  AOI21_X1  g671(.A(G113gat), .B1(new_n872), .B2(new_n777), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n871), .A2(new_n873), .ZN(G1340gat));
  INV_X1    g673(.A(G120gat), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n869), .A2(new_n875), .A3(new_n802), .ZN(new_n876));
  AOI21_X1  g675(.A(G120gat), .B1(new_n872), .B2(new_n633), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(G1341gat));
  OAI21_X1  g677(.A(G127gat), .B1(new_n869), .B2(new_n652), .ZN(new_n879));
  INV_X1    g678(.A(G127gat), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n872), .A2(new_n880), .A3(new_n651), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n882), .B(KEYINPUT115), .Z(G1342gat));
  INV_X1    g682(.A(G134gat), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n872), .A2(new_n884), .A3(new_n677), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n885), .A2(KEYINPUT56), .ZN(new_n886));
  OAI21_X1  g685(.A(G134gat), .B1(new_n869), .B2(new_n679), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(KEYINPUT56), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT116), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n886), .A2(new_n891), .A3(new_n887), .A4(new_n888), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(G1343gat));
  INV_X1    g692(.A(new_n868), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n740), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n426), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n853), .B1(new_n562), .B2(new_n859), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n677), .B1(new_n900), .B2(KEYINPUT118), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n851), .A2(new_n902), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(new_n849), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n652), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n899), .B1(new_n906), .B2(new_n828), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n897), .B1(new_n866), .B2(new_n426), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT117), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT113), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n677), .B1(new_n900), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n905), .B1(new_n912), .B2(new_n860), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n652), .B1(new_n913), .B2(new_n864), .ZN(new_n914));
  INV_X1    g713(.A(new_n865), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n828), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT57), .B1(new_n916), .B2(new_n424), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(KEYINPUT117), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n896), .B1(new_n910), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n212), .B1(new_n919), .B2(new_n777), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n866), .A2(new_n383), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n740), .A2(new_n437), .A3(new_n426), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n562), .A2(G141gat), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT119), .ZN(new_n927));
  OAI21_X1  g726(.A(KEYINPUT58), .B1(new_n920), .B2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n907), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n929), .B1(new_n917), .B2(KEYINPUT117), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n908), .A2(new_n909), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n777), .B(new_n895), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(G141gat), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT58), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n933), .A2(KEYINPUT119), .A3(new_n934), .A4(new_n926), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n928), .A2(new_n935), .ZN(G1344gat));
  NAND4_X1  g735(.A1(new_n924), .A2(new_n209), .A3(new_n210), .A4(new_n633), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n633), .B1(new_n895), .B2(KEYINPUT120), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n862), .A2(KEYINPUT114), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(new_n652), .A3(new_n865), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n899), .B1(new_n940), .B2(new_n828), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n843), .A2(new_n677), .A3(KEYINPUT121), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n942), .A2(new_n848), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT121), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n944), .B1(new_n679), .B2(new_n859), .ZN(new_n945));
  AOI22_X1  g744(.A1(new_n901), .A2(new_n903), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n828), .B1(new_n946), .B2(new_n651), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT57), .B1(new_n947), .B2(new_n424), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n941), .A2(new_n948), .ZN(new_n949));
  AOI211_X1 g748(.A(new_n938), .B(new_n949), .C1(KEYINPUT120), .C2(new_n895), .ZN(new_n950));
  NAND2_X1  g749(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n951));
  AOI22_X1  g750(.A1(new_n919), .A2(new_n633), .B1(new_n209), .B2(new_n210), .ZN(new_n952));
  OAI221_X1 g751(.A(new_n937), .B1(new_n950), .B2(new_n951), .C1(new_n952), .C2(KEYINPUT59), .ZN(G1345gat));
  AOI21_X1  g752(.A(new_n216), .B1(new_n919), .B2(new_n651), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n923), .A2(G155gat), .A3(new_n652), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n954), .A2(new_n955), .ZN(G1346gat));
  AOI21_X1  g755(.A(new_n217), .B1(new_n919), .B2(new_n677), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n923), .A2(G162gat), .A3(new_n679), .ZN(new_n958));
  OAI21_X1  g757(.A(KEYINPUT122), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n677), .B(new_n895), .C1(new_n930), .C2(new_n931), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(G162gat), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT122), .ZN(new_n962));
  INV_X1    g761(.A(new_n958), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n959), .A2(new_n964), .ZN(G1347gat));
  NOR2_X1   g764(.A1(new_n382), .A2(new_n489), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n696), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n867), .A2(new_n968), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n969), .A2(new_n292), .A3(new_n562), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n866), .A2(new_n489), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n486), .A2(new_n382), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(new_n777), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n970), .B1(new_n292), .B2(new_n975), .ZN(G1348gat));
  OAI21_X1  g775(.A(new_n306), .B1(new_n973), .B2(new_n634), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n728), .B1(new_n300), .B2(new_n299), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n977), .B1(new_n969), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n979), .B(KEYINPUT123), .ZN(G1349gat));
  OAI21_X1  g779(.A(G183gat), .B1(new_n969), .B2(new_n652), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n651), .A2(new_n339), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n981), .B1(new_n973), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n983), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g783(.A1(new_n974), .A2(new_n287), .A3(new_n677), .ZN(new_n985));
  OAI21_X1  g784(.A(G190gat), .B1(new_n969), .B2(new_n679), .ZN(new_n986));
  AND2_X1   g785(.A1(new_n986), .A2(KEYINPUT61), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n986), .A2(KEYINPUT61), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(G1351gat));
  INV_X1    g788(.A(KEYINPUT124), .ZN(new_n990));
  NOR3_X1   g789(.A1(new_n949), .A2(new_n740), .A3(new_n967), .ZN(new_n991));
  INV_X1    g790(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n990), .B1(new_n992), .B2(new_n562), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n991), .A2(KEYINPUT124), .A3(new_n777), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n993), .A2(G197gat), .A3(new_n994), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n740), .A2(new_n382), .A3(new_n426), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n971), .A2(new_n996), .ZN(new_n997));
  OR2_X1    g796(.A1(new_n562), .A2(G197gat), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(G1352gat));
  NOR3_X1   g798(.A1(new_n997), .A2(G204gat), .A3(new_n634), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT62), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g801(.A(G204gat), .B1(new_n992), .B2(new_n802), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1004));
  AND2_X1   g803(.A1(new_n1004), .A2(KEYINPUT125), .ZN(new_n1005));
  NOR2_X1   g804(.A1(new_n1004), .A2(KEYINPUT125), .ZN(new_n1006));
  OAI211_X1 g805(.A(new_n1002), .B(new_n1003), .C1(new_n1005), .C2(new_n1006), .ZN(G1353gat));
  INV_X1    g806(.A(KEYINPUT127), .ZN(new_n1008));
  NOR2_X1   g807(.A1(new_n740), .A2(new_n967), .ZN(new_n1009));
  OAI211_X1 g808(.A(new_n651), .B(new_n1009), .C1(new_n941), .C2(new_n948), .ZN(new_n1010));
  INV_X1    g809(.A(KEYINPUT126), .ZN(new_n1011));
  INV_X1    g810(.A(KEYINPUT63), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AND3_X1   g812(.A1(new_n1010), .A2(G211gat), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g813(.A(new_n1013), .B1(new_n1010), .B2(G211gat), .ZN(new_n1015));
  NOR2_X1   g814(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1016));
  NOR3_X1   g815(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  NOR3_X1   g816(.A1(new_n997), .A2(G211gat), .A3(new_n652), .ZN(new_n1018));
  OAI21_X1  g817(.A(new_n1008), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g818(.A(new_n1018), .ZN(new_n1020));
  INV_X1    g819(.A(new_n1016), .ZN(new_n1021));
  AND2_X1   g820(.A1(new_n1010), .A2(G211gat), .ZN(new_n1022));
  OAI21_X1  g821(.A(new_n1021), .B1(new_n1022), .B2(new_n1013), .ZN(new_n1023));
  OAI211_X1 g822(.A(KEYINPUT127), .B(new_n1020), .C1(new_n1023), .C2(new_n1014), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1019), .A2(new_n1024), .ZN(G1354gat));
  INV_X1    g824(.A(new_n997), .ZN(new_n1026));
  AOI21_X1  g825(.A(G218gat), .B1(new_n1026), .B2(new_n677), .ZN(new_n1027));
  NOR2_X1   g826(.A1(new_n679), .A2(new_n401), .ZN(new_n1028));
  AOI21_X1  g827(.A(new_n1027), .B1(new_n991), .B2(new_n1028), .ZN(G1355gat));
endmodule


