

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n527, n528, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U561 ( .A(n788), .B(KEYINPUT98), .ZN(n546) );
  INV_X1 U562 ( .A(KEYINPUT94), .ZN(n528) );
  AND2_X1 U563 ( .A1(n729), .A2(G2067), .ZN(n728) );
  AND2_X1 U564 ( .A1(n597), .A2(n596), .ZN(n599) );
  AND2_X1 U565 ( .A1(n595), .A2(n594), .ZN(n596) );
  INV_X2 U566 ( .A(G2104), .ZN(n577) );
  INV_X1 U567 ( .A(G2105), .ZN(n538) );
  XNOR2_X2 U568 ( .A(n527), .B(KEYINPUT103), .ZN(n556) );
  NAND2_X1 U569 ( .A1(n548), .A2(n549), .ZN(n527) );
  XNOR2_X1 U570 ( .A(n732), .B(n528), .ZN(n746) );
  NOR2_X1 U571 ( .A1(n749), .A2(n748), .ZN(n754) );
  NOR2_X1 U572 ( .A1(G651), .A2(n687), .ZN(n693) );
  NOR2_X2 U573 ( .A1(n821), .A2(G1966), .ZN(n766) );
  XOR2_X1 U574 ( .A(KEYINPUT107), .B(n870), .Z(n871) );
  AND2_X1 U575 ( .A1(n773), .A2(n772), .ZN(n775) );
  XOR2_X1 U576 ( .A(KEYINPUT97), .B(n785), .Z(n786) );
  NOR2_X1 U577 ( .A1(n754), .A2(n1023), .ZN(n756) );
  XNOR2_X1 U578 ( .A(n582), .B(KEYINPUT17), .ZN(n600) );
  AND2_X1 U579 ( .A1(G2105), .A2(G126), .ZN(n550) );
  BUF_X1 U580 ( .A(n724), .Z(G164) );
  BUF_X1 U581 ( .A(n790), .Z(n530) );
  XNOR2_X1 U582 ( .A(n732), .B(KEYINPUT94), .ZN(n531) );
  OR2_X1 U583 ( .A1(n1036), .A2(n733), .ZN(n741) );
  NOR2_X1 U584 ( .A1(n559), .A2(n535), .ZN(n558) );
  NOR2_X1 U585 ( .A1(n536), .A2(n561), .ZN(n559) );
  AND2_X1 U586 ( .A1(n768), .A2(G1996), .ZN(n737) );
  INV_X1 U587 ( .A(KEYINPUT28), .ZN(n755) );
  NOR2_X1 U588 ( .A1(n532), .A2(n543), .ZN(n542) );
  NOR2_X1 U589 ( .A1(KEYINPUT32), .A2(G8), .ZN(n543) );
  INV_X1 U590 ( .A(KEYINPUT101), .ZN(n817) );
  NOR2_X1 U591 ( .A1(n555), .A2(n823), .ZN(n554) );
  NAND2_X1 U592 ( .A1(n558), .A2(n533), .ZN(n553) );
  INV_X1 U593 ( .A(G651), .ZN(n569) );
  NOR2_X2 U594 ( .A1(n687), .A2(n569), .ZN(n680) );
  AND2_X2 U595 ( .A1(n538), .A2(G2104), .ZN(n607) );
  BUF_X1 U596 ( .A(n603), .Z(n925) );
  BUF_X1 U597 ( .A(n600), .Z(n930) );
  XNOR2_X1 U598 ( .A(n639), .B(n638), .ZN(n1036) );
  NOR2_X1 U599 ( .A1(n637), .A2(n636), .ZN(n639) );
  NAND2_X1 U600 ( .A1(n577), .A2(n550), .ZN(n593) );
  NOR2_X1 U601 ( .A1(n586), .A2(n585), .ZN(n726) );
  XOR2_X1 U602 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NOR2_X1 U603 ( .A1(n794), .A2(n793), .ZN(n532) );
  OR2_X1 U604 ( .A1(n560), .A2(KEYINPUT104), .ZN(n533) );
  AND2_X1 U605 ( .A1(n562), .A2(KEYINPUT104), .ZN(n534) );
  INV_X1 U606 ( .A(n1026), .ZN(n745) );
  AND2_X1 U607 ( .A1(n869), .A2(n1022), .ZN(n535) );
  AND2_X1 U608 ( .A1(n855), .A2(n864), .ZN(n536) );
  NOR2_X1 U609 ( .A1(n821), .A2(n807), .ZN(n537) );
  NAND2_X1 U610 ( .A1(KEYINPUT32), .A2(G8), .ZN(n545) );
  INV_X1 U611 ( .A(KEYINPUT104), .ZN(n561) );
  NAND2_X1 U612 ( .A1(n540), .A2(n539), .ZN(n544) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n539) );
  NAND2_X1 U614 ( .A1(n541), .A2(KEYINPUT32), .ZN(n540) );
  INV_X1 U615 ( .A(n546), .ZN(n541) );
  NAND2_X1 U616 ( .A1(n544), .A2(n542), .ZN(n804) );
  XNOR2_X1 U617 ( .A(n818), .B(n817), .ZN(n548) );
  NAND2_X1 U618 ( .A1(n798), .A2(n821), .ZN(n549) );
  AND2_X1 U619 ( .A1(n577), .A2(G2105), .ZN(n603) );
  NAND2_X1 U620 ( .A1(n551), .A2(n557), .ZN(n857) );
  NAND2_X1 U621 ( .A1(n552), .A2(n553), .ZN(n551) );
  NAND2_X1 U622 ( .A1(n556), .A2(n554), .ZN(n552) );
  NAND2_X1 U623 ( .A1(n556), .A2(n534), .ZN(n557) );
  INV_X1 U624 ( .A(n558), .ZN(n555) );
  INV_X1 U625 ( .A(n536), .ZN(n560) );
  INV_X1 U626 ( .A(n823), .ZN(n562) );
  INV_X1 U627 ( .A(G168), .ZN(n772) );
  INV_X1 U628 ( .A(KEYINPUT96), .ZN(n774) );
  INV_X1 U629 ( .A(KEYINPUT105), .ZN(n856) );
  INV_X1 U630 ( .A(KEYINPUT70), .ZN(n638) );
  BUF_X1 U631 ( .A(n607), .Z(n929) );
  BUF_X1 U632 ( .A(n726), .Z(G160) );
  XOR2_X1 U633 ( .A(G543), .B(KEYINPUT0), .Z(n687) );
  NAND2_X1 U634 ( .A1(G51), .A2(n693), .ZN(n566) );
  NOR2_X1 U635 ( .A1(G543), .A2(n569), .ZN(n564) );
  XNOR2_X1 U636 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n563) );
  XNOR2_X2 U637 ( .A(n564), .B(n563), .ZN(n692) );
  NAND2_X1 U638 ( .A1(G63), .A2(n692), .ZN(n565) );
  NAND2_X1 U639 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U640 ( .A(KEYINPUT6), .B(n567), .ZN(n574) );
  NOR2_X4 U641 ( .A1(G543), .A2(G651), .ZN(n677) );
  NAND2_X1 U642 ( .A1(n677), .A2(G89), .ZN(n568) );
  XNOR2_X1 U643 ( .A(n568), .B(KEYINPUT4), .ZN(n571) );
  NAND2_X1 U644 ( .A1(G76), .A2(n680), .ZN(n570) );
  NAND2_X1 U645 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U646 ( .A(n572), .B(KEYINPUT5), .Z(n573) );
  NOR2_X1 U647 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U648 ( .A(KEYINPUT7), .B(n575), .Z(n576) );
  XNOR2_X1 U649 ( .A(KEYINPUT72), .B(n576), .ZN(G168) );
  NAND2_X1 U650 ( .A1(G125), .A2(n603), .ZN(n578) );
  XNOR2_X1 U651 ( .A(n578), .B(KEYINPUT66), .ZN(n581) );
  NAND2_X1 U652 ( .A1(G101), .A2(n607), .ZN(n579) );
  XOR2_X1 U653 ( .A(KEYINPUT23), .B(n579), .Z(n580) );
  NAND2_X1 U654 ( .A1(n581), .A2(n580), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n538), .A2(n577), .ZN(n582) );
  NAND2_X1 U656 ( .A1(n600), .A2(G137), .ZN(n584) );
  AND2_X4 U657 ( .A1(G2105), .A2(G2104), .ZN(n926) );
  NAND2_X1 U658 ( .A1(n926), .A2(G113), .ZN(n583) );
  NAND2_X1 U659 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U660 ( .A1(G85), .A2(n677), .ZN(n588) );
  NAND2_X1 U661 ( .A1(G72), .A2(n680), .ZN(n587) );
  NAND2_X1 U662 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U663 ( .A1(G47), .A2(n693), .ZN(n590) );
  NAND2_X1 U664 ( .A1(G60), .A2(n692), .ZN(n589) );
  NAND2_X1 U665 ( .A1(n590), .A2(n589), .ZN(n591) );
  OR2_X1 U666 ( .A1(n592), .A2(n591), .ZN(G290) );
  XNOR2_X1 U667 ( .A(n593), .B(KEYINPUT86), .ZN(n597) );
  NAND2_X1 U668 ( .A1(G102), .A2(n607), .ZN(n595) );
  NAND2_X1 U669 ( .A1(G114), .A2(n926), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n600), .A2(G138), .ZN(n598) );
  AND2_X2 U671 ( .A1(n599), .A2(n598), .ZN(n724) );
  AND2_X1 U672 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U673 ( .A1(G111), .A2(n926), .ZN(n602) );
  NAND2_X1 U674 ( .A1(G135), .A2(n930), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n602), .A2(n601), .ZN(n606) );
  NAND2_X1 U676 ( .A1(n925), .A2(G123), .ZN(n604) );
  XOR2_X1 U677 ( .A(KEYINPUT18), .B(n604), .Z(n605) );
  NOR2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U679 ( .A1(n929), .A2(G99), .ZN(n608) );
  NAND2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n978) );
  XNOR2_X1 U681 ( .A(G2096), .B(n978), .ZN(n610) );
  OR2_X1 U682 ( .A1(G2100), .A2(n610), .ZN(G156) );
  INV_X1 U683 ( .A(G108), .ZN(G238) );
  INV_X1 U684 ( .A(G120), .ZN(G236) );
  INV_X1 U685 ( .A(G69), .ZN(G235) );
  INV_X1 U686 ( .A(G132), .ZN(G219) );
  INV_X1 U687 ( .A(G82), .ZN(G220) );
  NAND2_X1 U688 ( .A1(G52), .A2(n693), .ZN(n612) );
  NAND2_X1 U689 ( .A1(G64), .A2(n692), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n618) );
  NAND2_X1 U691 ( .A1(n680), .A2(G77), .ZN(n613) );
  XNOR2_X1 U692 ( .A(n613), .B(KEYINPUT68), .ZN(n615) );
  NAND2_X1 U693 ( .A1(G90), .A2(n677), .ZN(n614) );
  NAND2_X1 U694 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U695 ( .A(KEYINPUT9), .B(n616), .Z(n617) );
  NOR2_X1 U696 ( .A1(n618), .A2(n617), .ZN(G171) );
  NAND2_X1 U697 ( .A1(G75), .A2(n680), .ZN(n620) );
  NAND2_X1 U698 ( .A1(G50), .A2(n693), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n623) );
  NAND2_X1 U700 ( .A1(n677), .A2(G88), .ZN(n621) );
  XOR2_X1 U701 ( .A(KEYINPUT80), .B(n621), .Z(n622) );
  NOR2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n692), .A2(G62), .ZN(n624) );
  NAND2_X1 U704 ( .A1(n625), .A2(n624), .ZN(G303) );
  NAND2_X1 U705 ( .A1(G7), .A2(G661), .ZN(n626) );
  XNOR2_X1 U706 ( .A(n626), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U707 ( .A(G223), .ZN(n874) );
  NAND2_X1 U708 ( .A1(n874), .A2(G567), .ZN(n627) );
  XOR2_X1 U709 ( .A(KEYINPUT11), .B(n627), .Z(G234) );
  INV_X1 U710 ( .A(G860), .ZN(n660) );
  NAND2_X1 U711 ( .A1(G81), .A2(n677), .ZN(n628) );
  XOR2_X1 U712 ( .A(KEYINPUT12), .B(n628), .Z(n629) );
  XNOR2_X1 U713 ( .A(n629), .B(KEYINPUT69), .ZN(n631) );
  NAND2_X1 U714 ( .A1(G68), .A2(n680), .ZN(n630) );
  NAND2_X1 U715 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U716 ( .A(n632), .B(KEYINPUT13), .ZN(n634) );
  NAND2_X1 U717 ( .A1(G43), .A2(n693), .ZN(n633) );
  NAND2_X1 U718 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n692), .A2(G56), .ZN(n635) );
  XOR2_X1 U720 ( .A(KEYINPUT14), .B(n635), .Z(n636) );
  OR2_X1 U721 ( .A1(n660), .A2(n1036), .ZN(n640) );
  XOR2_X1 U722 ( .A(KEYINPUT71), .B(n640), .Z(G153) );
  INV_X1 U723 ( .A(G171), .ZN(G301) );
  NAND2_X1 U724 ( .A1(G868), .A2(G301), .ZN(n649) );
  NAND2_X1 U725 ( .A1(G54), .A2(n693), .ZN(n642) );
  NAND2_X1 U726 ( .A1(G66), .A2(n692), .ZN(n641) );
  NAND2_X1 U727 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U728 ( .A1(G92), .A2(n677), .ZN(n644) );
  NAND2_X1 U729 ( .A1(G79), .A2(n680), .ZN(n643) );
  NAND2_X1 U730 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U731 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U732 ( .A(n647), .B(KEYINPUT15), .ZN(n1026) );
  INV_X1 U733 ( .A(G868), .ZN(n656) );
  NAND2_X1 U734 ( .A1(n1026), .A2(n656), .ZN(n648) );
  NAND2_X1 U735 ( .A1(n649), .A2(n648), .ZN(G284) );
  NAND2_X1 U736 ( .A1(G91), .A2(n677), .ZN(n651) );
  NAND2_X1 U737 ( .A1(G78), .A2(n680), .ZN(n650) );
  NAND2_X1 U738 ( .A1(n651), .A2(n650), .ZN(n655) );
  NAND2_X1 U739 ( .A1(G53), .A2(n693), .ZN(n653) );
  NAND2_X1 U740 ( .A1(G65), .A2(n692), .ZN(n652) );
  NAND2_X1 U741 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U742 ( .A1(n655), .A2(n654), .ZN(n1023) );
  INV_X1 U743 ( .A(n1023), .ZN(G299) );
  NOR2_X1 U744 ( .A1(G286), .A2(n656), .ZN(n657) );
  XOR2_X1 U745 ( .A(KEYINPUT73), .B(n657), .Z(n659) );
  NOR2_X1 U746 ( .A1(G868), .A2(G299), .ZN(n658) );
  NOR2_X1 U747 ( .A1(n659), .A2(n658), .ZN(G297) );
  NAND2_X1 U748 ( .A1(n660), .A2(G559), .ZN(n661) );
  NAND2_X1 U749 ( .A1(n661), .A2(n745), .ZN(n662) );
  XNOR2_X1 U750 ( .A(n662), .B(KEYINPUT16), .ZN(n663) );
  XNOR2_X1 U751 ( .A(KEYINPUT74), .B(n663), .ZN(G148) );
  NOR2_X1 U752 ( .A1(n1036), .A2(G868), .ZN(n666) );
  NAND2_X1 U753 ( .A1(G868), .A2(n745), .ZN(n664) );
  NOR2_X1 U754 ( .A1(G559), .A2(n664), .ZN(n665) );
  NOR2_X1 U755 ( .A1(n666), .A2(n665), .ZN(G282) );
  NAND2_X1 U756 ( .A1(G55), .A2(n693), .ZN(n668) );
  NAND2_X1 U757 ( .A1(G67), .A2(n692), .ZN(n667) );
  NAND2_X1 U758 ( .A1(n668), .A2(n667), .ZN(n672) );
  NAND2_X1 U759 ( .A1(G93), .A2(n677), .ZN(n670) );
  NAND2_X1 U760 ( .A1(G80), .A2(n680), .ZN(n669) );
  NAND2_X1 U761 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U762 ( .A1(n672), .A2(n671), .ZN(n705) );
  XOR2_X1 U763 ( .A(n1036), .B(KEYINPUT75), .Z(n674) );
  NAND2_X1 U764 ( .A1(G559), .A2(n745), .ZN(n673) );
  XNOR2_X1 U765 ( .A(n674), .B(n673), .ZN(n702) );
  XNOR2_X1 U766 ( .A(KEYINPUT76), .B(n702), .ZN(n675) );
  NOR2_X1 U767 ( .A1(G860), .A2(n675), .ZN(n676) );
  XNOR2_X1 U768 ( .A(n705), .B(n676), .ZN(G145) );
  NAND2_X1 U769 ( .A1(G86), .A2(n677), .ZN(n679) );
  NAND2_X1 U770 ( .A1(G48), .A2(n693), .ZN(n678) );
  NAND2_X1 U771 ( .A1(n679), .A2(n678), .ZN(n684) );
  NAND2_X1 U772 ( .A1(G73), .A2(n680), .ZN(n681) );
  XNOR2_X1 U773 ( .A(n681), .B(KEYINPUT2), .ZN(n682) );
  XNOR2_X1 U774 ( .A(n682), .B(KEYINPUT79), .ZN(n683) );
  NOR2_X1 U775 ( .A1(n684), .A2(n683), .ZN(n686) );
  NAND2_X1 U776 ( .A1(n692), .A2(G61), .ZN(n685) );
  NAND2_X1 U777 ( .A1(n686), .A2(n685), .ZN(G305) );
  INV_X1 U778 ( .A(G303), .ZN(G166) );
  NAND2_X1 U779 ( .A1(n687), .A2(G87), .ZN(n688) );
  XNOR2_X1 U780 ( .A(n688), .B(KEYINPUT78), .ZN(n690) );
  NAND2_X1 U781 ( .A1(G74), .A2(G651), .ZN(n689) );
  NAND2_X1 U782 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U783 ( .A1(n692), .A2(n691), .ZN(n696) );
  NAND2_X1 U784 ( .A1(G49), .A2(n693), .ZN(n694) );
  XOR2_X1 U785 ( .A(KEYINPUT77), .B(n694), .Z(n695) );
  NAND2_X1 U786 ( .A1(n696), .A2(n695), .ZN(G288) );
  XNOR2_X1 U787 ( .A(G166), .B(KEYINPUT19), .ZN(n698) );
  XNOR2_X1 U788 ( .A(G290), .B(n1023), .ZN(n697) );
  XNOR2_X1 U789 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U790 ( .A(n705), .B(n699), .ZN(n700) );
  XNOR2_X1 U791 ( .A(n700), .B(G288), .ZN(n701) );
  XNOR2_X1 U792 ( .A(G305), .B(n701), .ZN(n944) );
  XNOR2_X1 U793 ( .A(n702), .B(n944), .ZN(n703) );
  NAND2_X1 U794 ( .A1(n703), .A2(G868), .ZN(n704) );
  XNOR2_X1 U795 ( .A(n704), .B(KEYINPUT81), .ZN(n707) );
  NOR2_X1 U796 ( .A1(n705), .A2(G868), .ZN(n706) );
  NOR2_X1 U797 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U798 ( .A(KEYINPUT82), .B(n708), .Z(G295) );
  NAND2_X1 U799 ( .A1(G2084), .A2(G2078), .ZN(n709) );
  XNOR2_X1 U800 ( .A(n709), .B(KEYINPUT83), .ZN(n710) );
  XNOR2_X1 U801 ( .A(KEYINPUT20), .B(n710), .ZN(n711) );
  NAND2_X1 U802 ( .A1(n711), .A2(G2090), .ZN(n712) );
  XNOR2_X1 U803 ( .A(KEYINPUT21), .B(n712), .ZN(n713) );
  NAND2_X1 U804 ( .A1(n713), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U805 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U806 ( .A1(G220), .A2(G219), .ZN(n714) );
  XOR2_X1 U807 ( .A(KEYINPUT22), .B(n714), .Z(n715) );
  NOR2_X1 U808 ( .A1(G218), .A2(n715), .ZN(n716) );
  NAND2_X1 U809 ( .A1(G96), .A2(n716), .ZN(n879) );
  NAND2_X1 U810 ( .A1(n879), .A2(G2106), .ZN(n722) );
  NOR2_X1 U811 ( .A1(G235), .A2(G236), .ZN(n717) );
  XNOR2_X1 U812 ( .A(KEYINPUT84), .B(n717), .ZN(n718) );
  NAND2_X1 U813 ( .A1(n718), .A2(G57), .ZN(n719) );
  NOR2_X1 U814 ( .A1(n719), .A2(G238), .ZN(n720) );
  XNOR2_X1 U815 ( .A(n720), .B(KEYINPUT85), .ZN(n878) );
  NAND2_X1 U816 ( .A1(n878), .A2(G567), .ZN(n721) );
  NAND2_X1 U817 ( .A1(n722), .A2(n721), .ZN(n900) );
  NAND2_X1 U818 ( .A1(G661), .A2(G483), .ZN(n723) );
  NOR2_X1 U819 ( .A1(n900), .A2(n723), .ZN(n877) );
  NAND2_X1 U820 ( .A1(n877), .A2(G36), .ZN(G176) );
  NOR2_X2 U821 ( .A1(n724), .A2(G1384), .ZN(n725) );
  XNOR2_X1 U822 ( .A(n725), .B(KEYINPUT65), .ZN(n842) );
  NAND2_X1 U823 ( .A1(n726), .A2(G40), .ZN(n843) );
  NOR2_X2 U824 ( .A1(n842), .A2(n843), .ZN(n727) );
  XNOR2_X2 U825 ( .A(n727), .B(KEYINPUT64), .ZN(n729) );
  XNOR2_X1 U826 ( .A(n728), .B(KEYINPUT93), .ZN(n731) );
  INV_X2 U827 ( .A(n729), .ZN(n765) );
  NAND2_X1 U828 ( .A1(G1348), .A2(n765), .ZN(n730) );
  NAND2_X1 U829 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U830 ( .A1(n531), .A2(n1026), .ZN(n743) );
  XNOR2_X1 U831 ( .A(KEYINPUT26), .B(KEYINPUT92), .ZN(n736) );
  NOR2_X1 U832 ( .A1(G1996), .A2(n736), .ZN(n733) );
  INV_X1 U833 ( .A(G1341), .ZN(n1059) );
  NAND2_X1 U834 ( .A1(n1059), .A2(n736), .ZN(n735) );
  INV_X2 U835 ( .A(n765), .ZN(n768) );
  INV_X1 U836 ( .A(n768), .ZN(n734) );
  NAND2_X1 U837 ( .A1(n735), .A2(n734), .ZN(n739) );
  NAND2_X1 U838 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U839 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U840 ( .A1(n741), .A2(n740), .ZN(n742) );
  AND2_X1 U841 ( .A1(n743), .A2(n742), .ZN(n753) );
  NAND2_X1 U842 ( .A1(n746), .A2(n745), .ZN(n751) );
  NAND2_X1 U843 ( .A1(G2072), .A2(n768), .ZN(n747) );
  XNOR2_X1 U844 ( .A(n747), .B(KEYINPUT27), .ZN(n749) );
  INV_X1 U845 ( .A(G1956), .ZN(n1058) );
  NOR2_X1 U846 ( .A1(n768), .A2(n1058), .ZN(n748) );
  NAND2_X1 U847 ( .A1(n754), .A2(n1023), .ZN(n750) );
  NAND2_X1 U848 ( .A1(n751), .A2(n750), .ZN(n752) );
  OR2_X2 U849 ( .A1(n753), .A2(n752), .ZN(n758) );
  XNOR2_X1 U850 ( .A(n756), .B(n755), .ZN(n757) );
  NAND2_X1 U851 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U852 ( .A(n759), .B(KEYINPUT29), .ZN(n763) );
  XOR2_X1 U853 ( .A(KEYINPUT25), .B(G2078), .Z(n1003) );
  NAND2_X1 U854 ( .A1(n1003), .A2(n768), .ZN(n761) );
  NAND2_X1 U855 ( .A1(n734), .A2(G1961), .ZN(n760) );
  NAND2_X1 U856 ( .A1(n761), .A2(n760), .ZN(n776) );
  NOR2_X1 U857 ( .A1(G301), .A2(n776), .ZN(n762) );
  NOR2_X1 U858 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U859 ( .A(n764), .B(KEYINPUT95), .ZN(n781) );
  NAND2_X2 U860 ( .A1(n765), .A2(G8), .ZN(n821) );
  XNOR2_X1 U861 ( .A(n766), .B(KEYINPUT91), .ZN(n789) );
  INV_X1 U862 ( .A(G8), .ZN(n769) );
  INV_X1 U863 ( .A(G2084), .ZN(n767) );
  AND2_X1 U864 ( .A1(n768), .A2(n767), .ZN(n791) );
  NOR2_X1 U865 ( .A1(n769), .A2(n791), .ZN(n770) );
  AND2_X1 U866 ( .A1(n789), .A2(n770), .ZN(n771) );
  XNOR2_X1 U867 ( .A(n771), .B(KEYINPUT30), .ZN(n773) );
  XNOR2_X1 U868 ( .A(n775), .B(n774), .ZN(n778) );
  NAND2_X1 U869 ( .A1(G301), .A2(n776), .ZN(n777) );
  NAND2_X1 U870 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U871 ( .A(n779), .B(KEYINPUT31), .ZN(n780) );
  NAND2_X1 U872 ( .A1(n781), .A2(n780), .ZN(n790) );
  NAND2_X1 U873 ( .A1(n790), .A2(G286), .ZN(n787) );
  NOR2_X1 U874 ( .A1(n734), .A2(G2090), .ZN(n783) );
  NOR2_X1 U875 ( .A1(G1971), .A2(n821), .ZN(n782) );
  NOR2_X1 U876 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U877 ( .A1(n784), .A2(G303), .ZN(n785) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n788) );
  INV_X1 U879 ( .A(n789), .ZN(n794) );
  NAND2_X1 U880 ( .A1(G8), .A2(n791), .ZN(n792) );
  NAND2_X1 U881 ( .A1(n530), .A2(n792), .ZN(n793) );
  NOR2_X1 U882 ( .A1(G2090), .A2(G303), .ZN(n795) );
  NAND2_X1 U883 ( .A1(G8), .A2(n795), .ZN(n796) );
  NAND2_X1 U884 ( .A1(n804), .A2(n796), .ZN(n797) );
  XNOR2_X1 U885 ( .A(n797), .B(KEYINPUT102), .ZN(n798) );
  OR2_X1 U886 ( .A1(G1971), .A2(G303), .ZN(n800) );
  NOR2_X1 U887 ( .A1(G288), .A2(G1976), .ZN(n799) );
  XNOR2_X1 U888 ( .A(n799), .B(KEYINPUT99), .ZN(n806) );
  AND2_X1 U889 ( .A1(n800), .A2(n806), .ZN(n802) );
  INV_X1 U890 ( .A(KEYINPUT33), .ZN(n801) );
  AND2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U892 ( .A1(n804), .A2(n803), .ZN(n816) );
  INV_X1 U893 ( .A(KEYINPUT100), .ZN(n807) );
  NAND2_X1 U894 ( .A1(G1976), .A2(G288), .ZN(n1024) );
  AND2_X1 U895 ( .A1(n537), .A2(n1024), .ZN(n805) );
  NOR2_X1 U896 ( .A1(KEYINPUT33), .A2(n805), .ZN(n814) );
  INV_X1 U897 ( .A(n806), .ZN(n1033) );
  NAND2_X1 U898 ( .A1(n807), .A2(n1033), .ZN(n810) );
  NAND2_X1 U899 ( .A1(n1033), .A2(KEYINPUT33), .ZN(n808) );
  NAND2_X1 U900 ( .A1(n808), .A2(KEYINPUT100), .ZN(n809) );
  NAND2_X1 U901 ( .A1(n810), .A2(n809), .ZN(n811) );
  OR2_X1 U902 ( .A1(n821), .A2(n811), .ZN(n812) );
  XOR2_X1 U903 ( .A(G1981), .B(G305), .Z(n1018) );
  NAND2_X1 U904 ( .A1(n812), .A2(n1018), .ZN(n813) );
  NOR2_X1 U905 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U906 ( .A1(n816), .A2(n815), .ZN(n818) );
  NOR2_X1 U907 ( .A1(G1981), .A2(G305), .ZN(n819) );
  XOR2_X1 U908 ( .A(n819), .B(KEYINPUT24), .Z(n820) );
  NOR2_X1 U909 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U910 ( .A(n822), .B(KEYINPUT90), .ZN(n823) );
  NAND2_X1 U911 ( .A1(G105), .A2(n929), .ZN(n824) );
  XNOR2_X1 U912 ( .A(n824), .B(KEYINPUT38), .ZN(n831) );
  NAND2_X1 U913 ( .A1(G117), .A2(n926), .ZN(n826) );
  NAND2_X1 U914 ( .A1(G141), .A2(n930), .ZN(n825) );
  NAND2_X1 U915 ( .A1(n826), .A2(n825), .ZN(n829) );
  NAND2_X1 U916 ( .A1(n925), .A2(G129), .ZN(n827) );
  XOR2_X1 U917 ( .A(KEYINPUT88), .B(n827), .Z(n828) );
  NOR2_X1 U918 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U919 ( .A1(n831), .A2(n830), .ZN(n910) );
  NAND2_X1 U920 ( .A1(G1996), .A2(n910), .ZN(n840) );
  NAND2_X1 U921 ( .A1(G95), .A2(n929), .ZN(n833) );
  NAND2_X1 U922 ( .A1(G131), .A2(n930), .ZN(n832) );
  NAND2_X1 U923 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U924 ( .A(KEYINPUT87), .B(n834), .ZN(n838) );
  NAND2_X1 U925 ( .A1(n925), .A2(G119), .ZN(n836) );
  NAND2_X1 U926 ( .A1(G107), .A2(n926), .ZN(n835) );
  AND2_X1 U927 ( .A1(n836), .A2(n835), .ZN(n837) );
  NAND2_X1 U928 ( .A1(n838), .A2(n837), .ZN(n909) );
  NAND2_X1 U929 ( .A1(G1991), .A2(n909), .ZN(n839) );
  NAND2_X1 U930 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U931 ( .A(KEYINPUT89), .B(n841), .ZN(n984) );
  INV_X1 U932 ( .A(n842), .ZN(n844) );
  NOR2_X1 U933 ( .A1(n844), .A2(n843), .ZN(n869) );
  INV_X1 U934 ( .A(n869), .ZN(n845) );
  NOR2_X1 U935 ( .A1(n984), .A2(n845), .ZN(n860) );
  INV_X1 U936 ( .A(n860), .ZN(n855) );
  XNOR2_X1 U937 ( .A(G2067), .B(KEYINPUT37), .ZN(n866) );
  NAND2_X1 U938 ( .A1(G104), .A2(n929), .ZN(n847) );
  NAND2_X1 U939 ( .A1(G140), .A2(n930), .ZN(n846) );
  NAND2_X1 U940 ( .A1(n847), .A2(n846), .ZN(n848) );
  XNOR2_X1 U941 ( .A(KEYINPUT34), .B(n848), .ZN(n853) );
  NAND2_X1 U942 ( .A1(G128), .A2(n925), .ZN(n850) );
  NAND2_X1 U943 ( .A1(G116), .A2(n926), .ZN(n849) );
  NAND2_X1 U944 ( .A1(n850), .A2(n849), .ZN(n851) );
  XOR2_X1 U945 ( .A(KEYINPUT35), .B(n851), .Z(n852) );
  NOR2_X1 U946 ( .A1(n853), .A2(n852), .ZN(n854) );
  XNOR2_X1 U947 ( .A(KEYINPUT36), .B(n854), .ZN(n939) );
  NOR2_X1 U948 ( .A1(n866), .A2(n939), .ZN(n980) );
  NAND2_X1 U949 ( .A1(n869), .A2(n980), .ZN(n864) );
  XNOR2_X1 U950 ( .A(G1986), .B(G290), .ZN(n1022) );
  XNOR2_X1 U951 ( .A(n857), .B(n856), .ZN(n872) );
  NOR2_X1 U952 ( .A1(G1996), .A2(n910), .ZN(n972) );
  NOR2_X1 U953 ( .A1(G1986), .A2(G290), .ZN(n858) );
  NOR2_X1 U954 ( .A1(G1991), .A2(n909), .ZN(n977) );
  NOR2_X1 U955 ( .A1(n858), .A2(n977), .ZN(n859) );
  NOR2_X1 U956 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U957 ( .A(n861), .B(KEYINPUT106), .ZN(n862) );
  NOR2_X1 U958 ( .A1(n972), .A2(n862), .ZN(n863) );
  XNOR2_X1 U959 ( .A(KEYINPUT39), .B(n863), .ZN(n865) );
  NAND2_X1 U960 ( .A1(n865), .A2(n864), .ZN(n867) );
  NAND2_X1 U961 ( .A1(n866), .A2(n939), .ZN(n974) );
  NAND2_X1 U962 ( .A1(n867), .A2(n974), .ZN(n868) );
  NAND2_X1 U963 ( .A1(n869), .A2(n868), .ZN(n870) );
  NAND2_X1 U964 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U965 ( .A(n873), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U966 ( .A1(G2106), .A2(n874), .ZN(G217) );
  AND2_X1 U967 ( .A1(G15), .A2(G2), .ZN(n875) );
  NAND2_X1 U968 ( .A1(G661), .A2(n875), .ZN(G259) );
  NAND2_X1 U969 ( .A1(G3), .A2(G1), .ZN(n876) );
  NAND2_X1 U970 ( .A1(n877), .A2(n876), .ZN(G188) );
  INV_X1 U972 ( .A(G96), .ZN(G221) );
  INV_X1 U973 ( .A(G57), .ZN(G237) );
  NOR2_X1 U974 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U975 ( .A(n880), .B(KEYINPUT110), .ZN(G325) );
  INV_X1 U976 ( .A(G325), .ZN(G261) );
  XOR2_X1 U977 ( .A(KEYINPUT111), .B(G2090), .Z(n882) );
  XNOR2_X1 U978 ( .A(G2067), .B(G2084), .ZN(n881) );
  XNOR2_X1 U979 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U980 ( .A(n883), .B(G2100), .Z(n885) );
  XNOR2_X1 U981 ( .A(G2078), .B(G2072), .ZN(n884) );
  XNOR2_X1 U982 ( .A(n885), .B(n884), .ZN(n889) );
  XOR2_X1 U983 ( .A(G2096), .B(G2678), .Z(n887) );
  XNOR2_X1 U984 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U986 ( .A(n889), .B(n888), .Z(G227) );
  XNOR2_X1 U987 ( .A(G1996), .B(KEYINPUT112), .ZN(n899) );
  XOR2_X1 U988 ( .A(G1991), .B(G1976), .Z(n891) );
  XNOR2_X1 U989 ( .A(G1981), .B(G1966), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n891), .B(n890), .ZN(n895) );
  XOR2_X1 U991 ( .A(G1971), .B(G1956), .Z(n893) );
  XNOR2_X1 U992 ( .A(G1986), .B(G1961), .ZN(n892) );
  XNOR2_X1 U993 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U994 ( .A(n895), .B(n894), .Z(n897) );
  XNOR2_X1 U995 ( .A(G2474), .B(KEYINPUT41), .ZN(n896) );
  XNOR2_X1 U996 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(G229) );
  INV_X1 U998 ( .A(n900), .ZN(G319) );
  NAND2_X1 U999 ( .A1(n925), .A2(G124), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n901), .B(KEYINPUT44), .ZN(n903) );
  NAND2_X1 U1001 ( .A1(G112), .A2(n926), .ZN(n902) );
  NAND2_X1 U1002 ( .A1(n903), .A2(n902), .ZN(n907) );
  NAND2_X1 U1003 ( .A1(G100), .A2(n929), .ZN(n905) );
  NAND2_X1 U1004 ( .A1(G136), .A2(n930), .ZN(n904) );
  NAND2_X1 U1005 ( .A1(n905), .A2(n904), .ZN(n906) );
  NOR2_X1 U1006 ( .A1(n907), .A2(n906), .ZN(G162) );
  XOR2_X1 U1007 ( .A(G164), .B(G162), .Z(n908) );
  XNOR2_X1 U1008 ( .A(n909), .B(n908), .ZN(n916) );
  XNOR2_X1 U1009 ( .A(G160), .B(n910), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(n911), .B(n978), .ZN(n912) );
  XOR2_X1 U1011 ( .A(n912), .B(KEYINPUT48), .Z(n914) );
  XNOR2_X1 U1012 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(n914), .B(n913), .ZN(n915) );
  XOR2_X1 U1014 ( .A(n916), .B(n915), .Z(n938) );
  NAND2_X1 U1015 ( .A1(G103), .A2(n929), .ZN(n918) );
  NAND2_X1 U1016 ( .A1(G139), .A2(n930), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n923) );
  NAND2_X1 U1018 ( .A1(G127), .A2(n925), .ZN(n920) );
  NAND2_X1 U1019 ( .A1(G115), .A2(n926), .ZN(n919) );
  NAND2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1021 ( .A(KEYINPUT47), .B(n921), .Z(n922) );
  NOR2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1023 ( .A(KEYINPUT113), .B(n924), .Z(n966) );
  NAND2_X1 U1024 ( .A1(G130), .A2(n925), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(G118), .A2(n926), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n935) );
  NAND2_X1 U1027 ( .A1(G106), .A2(n929), .ZN(n932) );
  NAND2_X1 U1028 ( .A1(G142), .A2(n930), .ZN(n931) );
  NAND2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1030 ( .A(KEYINPUT45), .B(n933), .Z(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(n966), .B(n936), .ZN(n937) );
  XNOR2_X1 U1033 ( .A(n938), .B(n937), .ZN(n940) );
  XNOR2_X1 U1034 ( .A(n940), .B(n939), .ZN(n941) );
  NOR2_X1 U1035 ( .A1(G37), .A2(n941), .ZN(G395) );
  XOR2_X1 U1036 ( .A(KEYINPUT115), .B(n1036), .Z(n943) );
  XNOR2_X1 U1037 ( .A(G171), .B(n745), .ZN(n942) );
  XNOR2_X1 U1038 ( .A(n943), .B(n942), .ZN(n945) );
  XNOR2_X1 U1039 ( .A(n945), .B(n944), .ZN(n946) );
  XOR2_X1 U1040 ( .A(n946), .B(G286), .Z(n947) );
  NOR2_X1 U1041 ( .A1(G37), .A2(n947), .ZN(G397) );
  XNOR2_X1 U1042 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n949) );
  NOR2_X1 U1043 ( .A1(G227), .A2(G229), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(n949), .B(n948), .ZN(n962) );
  XNOR2_X1 U1045 ( .A(G2451), .B(G2427), .ZN(n959) );
  XOR2_X1 U1046 ( .A(G2430), .B(G2443), .Z(n951) );
  XNOR2_X1 U1047 ( .A(G2435), .B(KEYINPUT109), .ZN(n950) );
  XNOR2_X1 U1048 ( .A(n951), .B(n950), .ZN(n955) );
  XOR2_X1 U1049 ( .A(G2438), .B(G2454), .Z(n953) );
  XNOR2_X1 U1050 ( .A(G1348), .B(G1341), .ZN(n952) );
  XNOR2_X1 U1051 ( .A(n953), .B(n952), .ZN(n954) );
  XOR2_X1 U1052 ( .A(n955), .B(n954), .Z(n957) );
  XNOR2_X1 U1053 ( .A(G2446), .B(KEYINPUT108), .ZN(n956) );
  XNOR2_X1 U1054 ( .A(n957), .B(n956), .ZN(n958) );
  XNOR2_X1 U1055 ( .A(n959), .B(n958), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n960), .A2(G14), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(G319), .A2(n965), .ZN(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(G395), .A2(G397), .ZN(n963) );
  NAND2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(G225) );
  INV_X1 U1061 ( .A(G225), .ZN(G308) );
  INV_X1 U1062 ( .A(n965), .ZN(G401) );
  INV_X1 U1063 ( .A(KEYINPUT55), .ZN(n1012) );
  XNOR2_X1 U1064 ( .A(G2072), .B(n966), .ZN(n967) );
  XNOR2_X1 U1065 ( .A(n967), .B(KEYINPUT119), .ZN(n969) );
  XOR2_X1 U1066 ( .A(G2078), .B(G164), .Z(n968) );
  NOR2_X1 U1067 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1068 ( .A(KEYINPUT50), .B(n970), .Z(n989) );
  XOR2_X1 U1069 ( .A(G2090), .B(G162), .Z(n971) );
  NOR2_X1 U1070 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1071 ( .A(KEYINPUT51), .B(n973), .Z(n975) );
  NAND2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n986) );
  XOR2_X1 U1073 ( .A(G160), .B(G2084), .Z(n976) );
  NOR2_X1 U1074 ( .A1(n977), .A2(n976), .ZN(n979) );
  NAND2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1077 ( .A(KEYINPUT117), .B(n982), .Z(n983) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1080 ( .A(KEYINPUT118), .B(n987), .Z(n988) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1082 ( .A(n990), .B(KEYINPUT52), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(n991), .B(KEYINPUT120), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n1012), .A2(n992), .ZN(n993) );
  NAND2_X1 U1085 ( .A1(n993), .A2(G29), .ZN(n1046) );
  XOR2_X1 U1086 ( .A(G2084), .B(G34), .Z(n994) );
  XNOR2_X1 U1087 ( .A(KEYINPUT54), .B(n994), .ZN(n1010) );
  XNOR2_X1 U1088 ( .A(G2090), .B(G35), .ZN(n1008) );
  XNOR2_X1 U1089 ( .A(G2067), .B(G26), .ZN(n996) );
  XNOR2_X1 U1090 ( .A(G32), .B(G1996), .ZN(n995) );
  NOR2_X1 U1091 ( .A1(n996), .A2(n995), .ZN(n1002) );
  XOR2_X1 U1092 ( .A(G2072), .B(G33), .Z(n997) );
  NAND2_X1 U1093 ( .A1(n997), .A2(G28), .ZN(n1000) );
  XOR2_X1 U1094 ( .A(G25), .B(G1991), .Z(n998) );
  XNOR2_X1 U1095 ( .A(KEYINPUT121), .B(n998), .ZN(n999) );
  NOR2_X1 U1096 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1097 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XNOR2_X1 U1098 ( .A(G27), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1099 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1100 ( .A(KEYINPUT53), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1101 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1103 ( .A(n1011), .B(KEYINPUT122), .ZN(n1013) );
  XNOR2_X1 U1104 ( .A(n1013), .B(n1012), .ZN(n1015) );
  INV_X1 U1105 ( .A(G29), .ZN(n1014) );
  NAND2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1107 ( .A1(G11), .A2(n1016), .ZN(n1044) );
  XNOR2_X1 U1108 ( .A(G16), .B(KEYINPUT56), .ZN(n1017) );
  XNOR2_X1 U1109 ( .A(n1017), .B(KEYINPUT123), .ZN(n1042) );
  XNOR2_X1 U1110 ( .A(G1966), .B(G168), .ZN(n1019) );
  NAND2_X1 U1111 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1112 ( .A(KEYINPUT57), .B(n1020), .ZN(n1035) );
  XNOR2_X1 U1113 ( .A(G1971), .B(G303), .ZN(n1021) );
  NOR2_X1 U1114 ( .A1(n1022), .A2(n1021), .ZN(n1031) );
  XNOR2_X1 U1115 ( .A(n1023), .B(G1956), .ZN(n1025) );
  NAND2_X1 U1116 ( .A1(n1025), .A2(n1024), .ZN(n1029) );
  XNOR2_X1 U1117 ( .A(G1348), .B(n1026), .ZN(n1027) );
  XNOR2_X1 U1118 ( .A(KEYINPUT124), .B(n1027), .ZN(n1028) );
  NOR2_X1 U1119 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1120 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1121 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1122 ( .A1(n1035), .A2(n1034), .ZN(n1040) );
  XNOR2_X1 U1123 ( .A(G171), .B(G1961), .ZN(n1038) );
  XNOR2_X1 U1124 ( .A(n1059), .B(n1036), .ZN(n1037) );
  NAND2_X1 U1125 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NOR2_X1 U1126 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  NOR2_X1 U1127 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  NOR2_X1 U1128 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  NAND2_X1 U1129 ( .A1(n1046), .A2(n1045), .ZN(n1074) );
  XNOR2_X1 U1130 ( .A(G1986), .B(G24), .ZN(n1051) );
  XNOR2_X1 U1131 ( .A(G1971), .B(G22), .ZN(n1048) );
  XNOR2_X1 U1132 ( .A(G1976), .B(G23), .ZN(n1047) );
  NOR2_X1 U1133 ( .A1(n1048), .A2(n1047), .ZN(n1049) );
  XNOR2_X1 U1134 ( .A(KEYINPUT127), .B(n1049), .ZN(n1050) );
  NOR2_X1 U1135 ( .A1(n1051), .A2(n1050), .ZN(n1052) );
  XNOR2_X1 U1136 ( .A(KEYINPUT58), .B(n1052), .ZN(n1056) );
  XNOR2_X1 U1137 ( .A(G1966), .B(G21), .ZN(n1054) );
  XNOR2_X1 U1138 ( .A(G5), .B(G1961), .ZN(n1053) );
  NOR2_X1 U1139 ( .A1(n1054), .A2(n1053), .ZN(n1055) );
  NAND2_X1 U1140 ( .A1(n1056), .A2(n1055), .ZN(n1070) );
  XOR2_X1 U1141 ( .A(G1348), .B(KEYINPUT59), .Z(n1057) );
  XNOR2_X1 U1142 ( .A(G4), .B(n1057), .ZN(n1066) );
  XNOR2_X1 U1143 ( .A(n1058), .B(G20), .ZN(n1061) );
  XNOR2_X1 U1144 ( .A(n1059), .B(G19), .ZN(n1060) );
  NAND2_X1 U1145 ( .A1(n1061), .A2(n1060), .ZN(n1063) );
  XNOR2_X1 U1146 ( .A(G6), .B(G1981), .ZN(n1062) );
  NOR2_X1 U1147 ( .A1(n1063), .A2(n1062), .ZN(n1064) );
  XNOR2_X1 U1148 ( .A(n1064), .B(KEYINPUT125), .ZN(n1065) );
  NOR2_X1 U1149 ( .A1(n1066), .A2(n1065), .ZN(n1067) );
  XOR2_X1 U1150 ( .A(KEYINPUT60), .B(n1067), .Z(n1068) );
  XNOR2_X1 U1151 ( .A(KEYINPUT126), .B(n1068), .ZN(n1069) );
  NOR2_X1 U1152 ( .A1(n1070), .A2(n1069), .ZN(n1071) );
  XOR2_X1 U1153 ( .A(KEYINPUT61), .B(n1071), .Z(n1072) );
  NOR2_X1 U1154 ( .A1(G16), .A2(n1072), .ZN(n1073) );
  NOR2_X1 U1155 ( .A1(n1074), .A2(n1073), .ZN(n1075) );
  XNOR2_X1 U1156 ( .A(n1075), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1157 ( .A(G311), .ZN(G150) );
endmodule

