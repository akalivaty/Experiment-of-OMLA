//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  XNOR2_X1  g000(.A(G110), .B(G122), .ZN(new_n187));
  OR2_X1    g001(.A1(new_n187), .A2(KEYINPUT85), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(KEYINPUT85), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT8), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(KEYINPUT8), .A3(new_n189), .ZN(new_n193));
  INV_X1    g007(.A(G104), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT3), .B1(new_n194), .B2(G107), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n196));
  INV_X1    g010(.A(G107), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(G104), .ZN(new_n198));
  INV_X1    g012(.A(G101), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n194), .A2(G107), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n195), .A2(new_n198), .A3(new_n199), .A4(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n197), .A2(G104), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n194), .A2(G107), .ZN(new_n203));
  OAI21_X1  g017(.A(G101), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  XOR2_X1   g020(.A(G116), .B(G119), .Z(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT2), .B(G113), .ZN(new_n208));
  OR2_X1    g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT5), .ZN(new_n210));
  INV_X1    g024(.A(G119), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(G116), .ZN(new_n212));
  OAI211_X1 g026(.A(G113), .B(new_n212), .C1(new_n207), .C2(new_n210), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n206), .A2(new_n209), .A3(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n206), .B1(new_n209), .B2(new_n213), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n192), .B(new_n193), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G953), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n217), .A2(G224), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT7), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G143), .ZN(new_n223));
  INV_X1    g037(.A(G143), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G146), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G128), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G128), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT1), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n232), .B1(G143), .B2(new_n222), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n226), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n223), .A2(new_n225), .A3(new_n232), .A4(G128), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G125), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G143), .B(G146), .ZN(new_n239));
  NAND2_X1  g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OR2_X1    g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n242), .A2(new_n240), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n241), .B1(new_n243), .B2(new_n239), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G125), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n238), .A2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n219), .A2(KEYINPUT87), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n221), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  AOI211_X1 g063(.A(new_n247), .B(new_n220), .C1(new_n238), .C2(new_n245), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n216), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OR2_X1    g065(.A1(new_n251), .A2(KEYINPUT88), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT84), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n214), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n195), .A2(new_n198), .A3(new_n200), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G101), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(KEYINPUT4), .A3(new_n201), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT77), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n207), .B(new_n208), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT77), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n256), .A2(new_n260), .A3(KEYINPUT4), .A4(new_n201), .ZN(new_n261));
  OR2_X1    g075(.A1(new_n256), .A2(KEYINPUT4), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n258), .A2(new_n259), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n213), .A2(new_n209), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT84), .B1(new_n264), .B2(new_n205), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n254), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n251), .A2(KEYINPUT88), .B1(new_n266), .B2(new_n190), .ZN(new_n267));
  AOI21_X1  g081(.A(G902), .B1(new_n252), .B2(new_n267), .ZN(new_n268));
  XOR2_X1   g082(.A(new_n246), .B(new_n218), .Z(new_n269));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n254), .A2(new_n263), .A3(new_n265), .ZN(new_n271));
  XOR2_X1   g085(.A(new_n190), .B(KEYINPUT86), .Z(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n254), .A2(new_n263), .A3(new_n190), .A4(new_n265), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT6), .B1(new_n271), .B2(new_n272), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n269), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n268), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(G210), .B1(G237), .B2(G902), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT89), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n268), .A2(new_n277), .A3(new_n279), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n268), .A2(new_n277), .A3(new_n279), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT89), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(G237), .A2(G953), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G214), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n224), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(G143), .A3(G214), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(KEYINPUT18), .A2(G131), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n290), .A2(KEYINPUT18), .A3(G131), .A4(new_n291), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G140), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G125), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n237), .A2(G140), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n222), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n298), .A2(new_n299), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G146), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n301), .A2(KEYINPUT90), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT90), .B1(new_n301), .B2(new_n303), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n296), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G131), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n290), .A2(new_n307), .A3(new_n291), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT91), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n292), .A2(G131), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT91), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n290), .A2(new_n311), .A3(new_n307), .A4(new_n291), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n309), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT73), .A4(KEYINPUT16), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT16), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(new_n298), .B2(KEYINPUT16), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n314), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G146), .ZN(new_n319));
  OR2_X1    g133(.A1(new_n302), .A2(KEYINPUT19), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n302), .A2(KEYINPUT19), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n222), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n306), .B1(new_n313), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(G113), .B(G122), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(new_n194), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT17), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n309), .A2(new_n310), .A3(new_n329), .A4(new_n312), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n222), .B(new_n314), .C1(new_n315), .C2(new_n317), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n292), .A2(KEYINPUT17), .A3(G131), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n330), .A2(new_n331), .A3(new_n319), .A4(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(new_n326), .A3(new_n306), .ZN(new_n334));
  AOI21_X1  g148(.A(G475), .B1(new_n328), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G902), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n335), .A2(KEYINPUT20), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT20), .B1(new_n335), .B2(new_n336), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n334), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n326), .B1(new_n333), .B2(new_n306), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n336), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G475), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G952), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n345), .A2(KEYINPUT95), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n345), .A2(KEYINPUT95), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n217), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n348), .B1(G234), .B2(G237), .ZN(new_n349));
  XOR2_X1   g163(.A(new_n349), .B(KEYINPUT96), .Z(new_n350));
  XOR2_X1   g164(.A(KEYINPUT21), .B(G898), .Z(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  AOI211_X1 g166(.A(new_n336), .B(new_n217), .C1(G234), .C2(G237), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT92), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT66), .B(G128), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n356), .B1(new_n357), .B2(new_n224), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n231), .A2(KEYINPUT92), .A3(G143), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n227), .A2(G143), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT13), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n363), .A2(new_n365), .A3(G134), .ZN(new_n366));
  INV_X1    g180(.A(G134), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n360), .B(new_n362), .C1(new_n364), .C2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G122), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(G116), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(G116), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(new_n197), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n366), .A2(new_n368), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT14), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n372), .B1(new_n370), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT93), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT94), .B1(new_n371), .B2(KEYINPUT14), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT94), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n370), .A2(new_n381), .A3(new_n376), .ZN(new_n382));
  OAI211_X1 g196(.A(KEYINPUT93), .B(new_n372), .C1(new_n370), .C2(new_n376), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n379), .A2(new_n380), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G107), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n373), .A2(new_n197), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n367), .B1(new_n360), .B2(new_n362), .ZN(new_n387));
  AOI211_X1 g201(.A(G134), .B(new_n361), .C1(new_n358), .C2(new_n359), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n385), .B(new_n386), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  XOR2_X1   g203(.A(KEYINPUT9), .B(G234), .Z(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G217), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n391), .A2(new_n392), .A3(G953), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n375), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n393), .B1(new_n375), .B2(new_n389), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n336), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G478), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(KEYINPUT15), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  OAI221_X1 g214(.A(new_n336), .B1(KEYINPUT15), .B2(new_n398), .C1(new_n395), .C2(new_n396), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n344), .A2(new_n355), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(G214), .B1(G237), .B2(G902), .ZN(new_n404));
  INV_X1    g218(.A(G221), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n405), .B1(new_n390), .B2(new_n336), .ZN(new_n406));
  XNOR2_X1  g220(.A(G110), .B(G140), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n217), .A2(G227), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n407), .B(new_n408), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n258), .A2(new_n244), .A3(new_n261), .A4(new_n262), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT78), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n256), .A2(KEYINPUT4), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(KEYINPUT77), .B2(new_n257), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n414), .A2(KEYINPUT78), .A3(new_n244), .A4(new_n261), .ZN(new_n415));
  INV_X1    g229(.A(G137), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n416), .B1(KEYINPUT11), .B2(G134), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT64), .B(G137), .ZN(new_n418));
  AND2_X1   g232(.A1(KEYINPUT11), .A2(G134), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT11), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n367), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n307), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  AND2_X1   g237(.A1(KEYINPUT64), .A2(G137), .ZN(new_n424));
  NOR2_X1   g238(.A1(KEYINPUT64), .A2(G137), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n419), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(G137), .B1(new_n421), .B2(new_n367), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n426), .A2(new_n307), .A3(new_n422), .A4(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT79), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n235), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n239), .A2(KEYINPUT79), .A3(new_n232), .A4(G128), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n226), .B1(new_n233), .B2(new_n227), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n206), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT10), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n437), .B1(new_n234), .B2(new_n235), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n436), .A2(new_n437), .B1(new_n206), .B2(new_n438), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n412), .A2(new_n415), .A3(new_n430), .A4(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT80), .B1(new_n206), .B2(new_n236), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT80), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n205), .A2(new_n442), .A3(new_n234), .A4(new_n235), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n436), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n430), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT12), .ZN(new_n447));
  OR2_X1    g261(.A1(new_n447), .A2(KEYINPUT81), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(KEYINPUT81), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n446), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n444), .A2(KEYINPUT81), .A3(new_n447), .A4(new_n445), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n440), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n409), .B1(new_n452), .B2(KEYINPUT82), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT82), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n440), .A2(new_n450), .A3(new_n454), .A4(new_n451), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n440), .A2(new_n409), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n412), .A2(new_n439), .A3(new_n415), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n445), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n453), .A2(new_n455), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(G469), .B1(new_n460), .B2(G902), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n409), .B1(new_n459), .B2(new_n440), .ZN(new_n462));
  AND4_X1   g276(.A1(new_n440), .A2(new_n450), .A3(new_n451), .A4(new_n409), .ZN(new_n463));
  OR2_X1    g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(KEYINPUT83), .A2(G469), .ZN(new_n465));
  OR2_X1    g279(.A1(KEYINPUT83), .A2(G469), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n464), .A2(new_n336), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n406), .B1(new_n461), .B2(new_n467), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n287), .A2(new_n403), .A3(new_n404), .A4(new_n468), .ZN(new_n469));
  XOR2_X1   g283(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n470));
  NAND2_X1  g284(.A1(new_n288), .A2(G210), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n470), .B(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT26), .B(G101), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n472), .B(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n244), .B1(new_n423), .B2(new_n429), .ZN(new_n475));
  INV_X1    g289(.A(new_n259), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n367), .B1(new_n424), .B2(new_n425), .ZN(new_n477));
  NAND2_X1  g291(.A1(G134), .A2(G137), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(G131), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT65), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT65), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n477), .A2(new_n481), .A3(G131), .A4(new_n478), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n480), .A2(new_n236), .A3(new_n428), .A4(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n475), .A2(new_n476), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n476), .B1(new_n475), .B2(new_n483), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT28), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT69), .ZN(new_n488));
  AND4_X1   g302(.A1(new_n428), .A2(new_n480), .A3(new_n236), .A4(new_n482), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n426), .A2(new_n422), .A3(new_n427), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G131), .ZN(new_n491));
  OR2_X1    g305(.A1(new_n243), .A2(new_n239), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n491), .A2(new_n428), .B1(new_n492), .B2(new_n241), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT70), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT70), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n475), .A2(new_n495), .A3(new_n483), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n496), .A3(new_n476), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT28), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT69), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n500), .B(KEYINPUT28), .C1(new_n485), .C2(new_n486), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n488), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n474), .B1(new_n502), .B2(KEYINPUT29), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT71), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n487), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n487), .A2(new_n504), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n499), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n336), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT30), .B1(new_n489), .B2(new_n493), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT30), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n475), .A2(new_n510), .A3(new_n483), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n485), .B1(new_n512), .B2(new_n259), .ZN(new_n513));
  INV_X1    g327(.A(new_n474), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT29), .B1(new_n503), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(G472), .B1(new_n508), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(G472), .A2(G902), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n475), .A2(new_n510), .A3(new_n483), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n510), .B1(new_n475), .B2(new_n483), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n259), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n522), .A2(new_n474), .A3(new_n484), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n523), .A2(KEYINPUT31), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(KEYINPUT68), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT68), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n522), .A2(new_n526), .A3(new_n474), .A4(new_n484), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n524), .B1(new_n528), .B2(KEYINPUT31), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n502), .A2(new_n514), .ZN(new_n530));
  AOI211_X1 g344(.A(KEYINPUT32), .B(new_n519), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT32), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n526), .B1(new_n513), .B2(new_n474), .ZN(new_n533));
  INV_X1    g347(.A(new_n527), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT31), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n524), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n530), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n532), .B1(new_n537), .B2(new_n518), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n517), .B1(new_n531), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n229), .A2(G128), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n541));
  OAI211_X1 g355(.A(KEYINPUT23), .B(G119), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT72), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT23), .B1(new_n227), .B2(G119), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n544), .B1(new_n211), .B2(G128), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT72), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n231), .A2(new_n546), .A3(KEYINPUT23), .A4(G119), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n543), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G110), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n319), .A2(new_n331), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n211), .A2(G128), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n551), .B1(new_n357), .B2(new_n211), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT24), .B(G110), .ZN(new_n553));
  OR2_X1    g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n549), .A2(new_n550), .A3(new_n554), .ZN(new_n555));
  XOR2_X1   g369(.A(KEYINPUT74), .B(G110), .Z(new_n556));
  NAND4_X1  g370(.A1(new_n543), .A2(new_n545), .A3(new_n547), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n552), .A2(new_n553), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n301), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n560), .B1(new_n318), .B2(G146), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT76), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT76), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n555), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT75), .B(KEYINPUT22), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(G137), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n217), .A2(G221), .A3(G234), .ZN(new_n569));
  XOR2_X1   g383(.A(new_n568), .B(new_n569), .Z(new_n570));
  NAND3_X1  g384(.A1(new_n564), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n570), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n572), .A2(new_n565), .A3(new_n555), .A4(new_n562), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT25), .B1(new_n574), .B2(G902), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n392), .B1(G234), .B2(new_n336), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n571), .A2(new_n573), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT25), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n578), .A3(new_n336), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n575), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n576), .A2(G902), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n539), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n469), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(new_n199), .ZN(G3));
  INV_X1    g401(.A(G472), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n588), .B1(new_n537), .B2(new_n336), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n537), .A2(new_n518), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n468), .A2(new_n590), .A3(new_n591), .A4(new_n584), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n395), .A2(new_n396), .A3(KEYINPUT33), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT33), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n375), .A2(new_n389), .ZN(new_n596));
  INV_X1    g410(.A(new_n393), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n595), .B1(new_n598), .B2(new_n394), .ZN(new_n599));
  OAI211_X1 g413(.A(G478), .B(new_n336), .C1(new_n594), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(KEYINPUT97), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n397), .A2(new_n398), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT33), .B1(new_n395), .B2(new_n396), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n598), .A2(new_n595), .A3(new_n394), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n605), .A2(new_n606), .A3(G478), .A4(new_n336), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n601), .A2(new_n602), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n344), .ZN(new_n609));
  INV_X1    g423(.A(new_n355), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n279), .B1(new_n268), .B2(new_n277), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n610), .B(new_n404), .C1(new_n285), .C2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n593), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT34), .B(G104), .ZN(new_n615));
  XOR2_X1   g429(.A(new_n615), .B(KEYINPUT98), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n614), .B(new_n616), .ZN(G6));
  INV_X1    g431(.A(new_n402), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n612), .A2(new_n618), .A3(new_n344), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n592), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT35), .B(G107), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G9));
  AOI21_X1  g437(.A(new_n578), .B1(new_n577), .B2(new_n336), .ZN(new_n624));
  AOI211_X1 g438(.A(KEYINPUT25), .B(G902), .C1(new_n571), .C2(new_n573), .ZN(new_n625));
  INV_X1    g439(.A(new_n576), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n572), .A2(KEYINPUT36), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(new_n563), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n581), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT99), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n580), .A2(new_n633), .A3(new_n630), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(new_n591), .A3(new_n590), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n469), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT37), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G110), .ZN(G12));
  INV_X1    g453(.A(G900), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n353), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n350), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n339), .A2(new_n402), .A3(new_n343), .A4(new_n643), .ZN(new_n644));
  AOI211_X1 g458(.A(new_n406), .B(new_n644), .C1(new_n461), .C2(new_n467), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n404), .B1(new_n285), .B2(new_n611), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n539), .A2(new_n645), .A3(new_n647), .A4(new_n635), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  INV_X1    g463(.A(KEYINPUT100), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n284), .A2(new_n650), .A3(new_n286), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n650), .B1(new_n284), .B2(new_n286), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT38), .ZN(new_n653));
  OR3_X1    g467(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n653), .B1(new_n651), .B2(new_n652), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n624), .A2(new_n625), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n631), .B1(new_n658), .B2(new_n576), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n344), .A2(new_n402), .A3(new_n404), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT102), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n514), .B1(new_n485), .B2(new_n486), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n528), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(G472), .B1(new_n665), .B2(G902), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n666), .B1(new_n531), .B2(new_n538), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI211_X1 g483(.A(KEYINPUT101), .B(new_n666), .C1(new_n531), .C2(new_n538), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n642), .B(KEYINPUT103), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT39), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n468), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT40), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n657), .A2(new_n663), .A3(new_n671), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G143), .ZN(G45));
  NAND3_X1  g491(.A1(new_n539), .A2(new_n647), .A3(new_n635), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n608), .A2(new_n344), .A3(new_n643), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT104), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n608), .A2(new_n681), .A3(new_n344), .A4(new_n643), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n680), .A2(new_n468), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n222), .ZN(G48));
  INV_X1    g499(.A(new_n406), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n336), .B1(new_n462), .B2(new_n463), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(G469), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n467), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n539), .A2(new_n613), .A3(new_n584), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  NOR3_X1   g507(.A1(new_n585), .A2(new_n620), .A3(new_n689), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n694), .B(G116), .Z(G18));
  NAND4_X1  g509(.A1(new_n539), .A2(new_n647), .A3(new_n635), .A4(new_n690), .ZN(new_n696));
  INV_X1    g510(.A(new_n403), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(new_n211), .ZN(G21));
  NAND2_X1  g513(.A1(new_n507), .A2(new_n514), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n519), .B1(new_n529), .B2(new_n700), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n589), .A2(new_n583), .A3(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n612), .A2(new_n618), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n702), .A2(new_n344), .A3(new_n703), .A4(new_n690), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G122), .ZN(G24));
  NOR3_X1   g519(.A1(new_n589), .A2(new_n659), .A3(new_n701), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n689), .A2(new_n646), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n706), .A2(new_n680), .A3(new_n707), .A4(new_n682), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT105), .B(G125), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G27));
  OAI21_X1  g524(.A(KEYINPUT106), .B1(new_n531), .B2(new_n538), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n502), .A2(new_n514), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT31), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n713), .B1(new_n525), .B2(new_n527), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n712), .A2(new_n714), .A3(new_n524), .ZN(new_n715));
  OAI21_X1  g529(.A(KEYINPUT32), .B1(new_n715), .B2(new_n519), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n537), .A2(new_n532), .A3(new_n518), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n711), .A2(new_n719), .A3(new_n517), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n720), .A2(KEYINPUT42), .A3(new_n584), .ZN(new_n721));
  INV_X1    g535(.A(new_n404), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n284), .B2(new_n286), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n680), .A2(new_n723), .A3(new_n468), .A4(new_n682), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n721), .A2(KEYINPUT107), .A3(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n720), .A2(KEYINPUT42), .A3(new_n584), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n727), .B1(new_n728), .B2(new_n724), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT42), .ZN(new_n730));
  AND4_X1   g544(.A1(new_n539), .A2(new_n584), .A3(new_n468), .A4(new_n723), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n680), .A2(new_n682), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  AOI22_X1  g548(.A1(new_n726), .A2(new_n729), .B1(new_n730), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n307), .ZN(G33));
  INV_X1    g550(.A(new_n644), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n731), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G134), .ZN(G36));
  NAND2_X1  g553(.A1(G469), .A2(G902), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n453), .A2(new_n455), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n456), .B1(new_n445), .B2(new_n458), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n460), .A2(KEYINPUT45), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(G469), .A3(new_n745), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n746), .A2(KEYINPUT108), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(KEYINPUT108), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n740), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT46), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT109), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n746), .B(KEYINPUT108), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n753), .A2(new_n754), .A3(KEYINPUT46), .A4(new_n740), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n751), .A2(new_n752), .A3(new_n467), .A4(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n686), .A3(new_n673), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n756), .A2(KEYINPUT110), .A3(new_n686), .A4(new_n673), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n344), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n608), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT43), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n590), .A2(new_n591), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n766), .A3(new_n660), .ZN(new_n767));
  XOR2_X1   g581(.A(new_n767), .B(KEYINPUT44), .Z(new_n768));
  INV_X1    g582(.A(new_n723), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n761), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G137), .ZN(G39));
  NOR3_X1   g586(.A1(new_n769), .A2(new_n539), .A3(new_n584), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n756), .A2(KEYINPUT47), .A3(new_n686), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT47), .B1(new_n756), .B2(new_n686), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n733), .B(new_n773), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G140), .ZN(G42));
  NAND2_X1  g592(.A1(new_n467), .A2(new_n688), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT49), .ZN(new_n780));
  NOR4_X1   g594(.A1(new_n657), .A2(new_n406), .A3(new_n763), .A4(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n669), .A2(new_n670), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n781), .A2(new_n584), .A3(new_n404), .A4(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT113), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n691), .B(new_n704), .C1(new_n696), .C2(new_n697), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n694), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n344), .A2(new_n642), .ZN(new_n787));
  XOR2_X1   g601(.A(new_n402), .B(KEYINPUT111), .Z(new_n788));
  NAND4_X1  g602(.A1(new_n539), .A2(new_n635), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n706), .A2(new_n680), .A3(new_n682), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n468), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n769), .A2(new_n792), .ZN(new_n793));
  AOI22_X1  g607(.A1(new_n791), .A2(new_n793), .B1(new_n731), .B2(new_n737), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n469), .B1(new_n585), .B2(new_n636), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n609), .B1(new_n788), .B2(new_n344), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(new_n610), .A3(new_n287), .A4(new_n404), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n592), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n786), .A2(new_n794), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n734), .A2(new_n730), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT107), .B1(new_n721), .B2(new_n725), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n728), .A2(new_n727), .A3(new_n724), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT112), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n648), .B(new_n708), .C1(new_n678), .C2(new_n683), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n792), .A2(new_n642), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n661), .B1(new_n283), .B2(new_n281), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n671), .A2(new_n659), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n808), .A2(KEYINPUT52), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT52), .B1(new_n808), .B2(new_n811), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n806), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n815));
  INV_X1    g629(.A(new_n811), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n815), .B1(new_n816), .B2(new_n807), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n808), .A2(KEYINPUT52), .A3(new_n811), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(KEYINPUT112), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n805), .B1(new_n814), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n784), .B1(new_n820), .B2(KEYINPUT53), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n800), .B(new_n804), .C1(new_n813), .C2(new_n812), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n786), .A2(new_n794), .A3(new_n799), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n735), .A2(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n812), .A2(new_n813), .A3(new_n806), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT112), .B1(new_n817), .B2(new_n818), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(KEYINPUT113), .A3(new_n823), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n821), .A2(new_n824), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT54), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n833), .A2(KEYINPUT51), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(KEYINPUT51), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n702), .A2(new_n690), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n837));
  INV_X1    g651(.A(new_n350), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n765), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n763), .A2(new_n764), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT43), .B1(new_n608), .B2(new_n762), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT116), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n836), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n404), .B1(new_n654), .B2(new_n655), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n769), .A2(new_n689), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n839), .B2(new_n843), .ZN(new_n849));
  AOI22_X1  g663(.A1(new_n846), .A2(KEYINPUT50), .B1(new_n706), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT50), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n844), .A2(new_n851), .A3(new_n845), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n583), .A2(new_n350), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n782), .A2(new_n847), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n782), .A2(KEYINPUT117), .A3(new_n847), .A4(new_n853), .ZN(new_n857));
  INV_X1    g671(.A(new_n608), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n856), .A2(new_n762), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n850), .A2(new_n852), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n860), .B(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n756), .A2(new_n686), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT47), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n467), .A2(new_n406), .A3(new_n688), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n865), .A2(new_n774), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n723), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n839), .A2(new_n843), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n702), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n834), .B(new_n835), .C1(new_n862), .C2(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(KEYINPUT51), .B(new_n860), .C1(new_n868), .C2(new_n870), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n720), .A2(new_n584), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n849), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT119), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT48), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n870), .A2(new_n646), .A3(new_n689), .ZN(new_n878));
  INV_X1    g692(.A(new_n609), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n856), .A2(new_n857), .ZN(new_n880));
  AOI211_X1 g694(.A(new_n348), .B(new_n878), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n873), .A2(new_n877), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT114), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n822), .A2(new_n883), .A3(new_n823), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n883), .B1(new_n822), .B2(new_n823), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n887));
  OAI211_X1 g701(.A(KEYINPUT53), .B(new_n826), .C1(new_n827), .C2(new_n828), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AND4_X1   g703(.A1(new_n832), .A2(new_n872), .A3(new_n882), .A4(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(G952), .A2(G953), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n783), .B1(new_n890), .B2(new_n891), .ZN(G75));
  NOR2_X1   g706(.A1(new_n812), .A2(new_n813), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n823), .B1(new_n805), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT114), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n822), .A2(new_n883), .A3(new_n823), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(new_n888), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(G210), .A3(G902), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT56), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n275), .A2(new_n276), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n269), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT55), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n898), .A2(new_n899), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n903), .B1(new_n898), .B2(new_n899), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n217), .A2(G952), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(G51));
  XOR2_X1   g721(.A(new_n740), .B(KEYINPUT57), .Z(new_n908));
  AOI21_X1  g722(.A(new_n887), .B1(new_n886), .B2(new_n888), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n897), .A2(KEYINPUT54), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n464), .ZN(new_n912));
  INV_X1    g726(.A(new_n753), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n897), .A2(G902), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n906), .B1(new_n912), .B2(new_n914), .ZN(G54));
  AND2_X1   g729(.A1(KEYINPUT58), .A2(G475), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n916), .A2(KEYINPUT120), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(KEYINPUT120), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n897), .A2(G902), .A3(new_n917), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n328), .A2(new_n334), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n919), .A2(new_n921), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n922), .A2(new_n923), .A3(new_n906), .ZN(G60));
  NAND2_X1  g738(.A1(new_n832), .A2(new_n889), .ZN(new_n925));
  NAND2_X1  g739(.A1(G478), .A2(G902), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT59), .Z(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n605), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n927), .B1(new_n603), .B2(new_n604), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n909), .B2(new_n910), .ZN(new_n931));
  INV_X1    g745(.A(new_n906), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n929), .A2(new_n933), .ZN(G63));
  NAND2_X1  g748(.A1(G217), .A2(G902), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT121), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT60), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n897), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n574), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n897), .A2(new_n629), .A3(new_n937), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n939), .A2(new_n932), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n939), .A2(KEYINPUT61), .A3(new_n932), .A4(new_n940), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(G66));
  AOI21_X1  g759(.A(new_n217), .B1(new_n351), .B2(G224), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n786), .A2(new_n799), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(new_n217), .ZN(new_n948));
  INV_X1    g762(.A(G898), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n900), .B1(new_n949), .B2(G953), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n948), .B(new_n950), .ZN(G69));
  XNOR2_X1  g765(.A(KEYINPUT122), .B(KEYINPUT123), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n512), .B(new_n952), .Z(new_n953));
  NAND2_X1  g767(.A1(new_n320), .A2(new_n321), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n804), .A2(KEYINPUT125), .A3(new_n738), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n804), .A2(new_n738), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT125), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n874), .A2(new_n810), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n768), .B2(new_n769), .ZN(new_n962));
  AOI22_X1  g776(.A1(new_n957), .A2(new_n960), .B1(new_n761), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n732), .B1(new_n865), .B2(new_n774), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n807), .B1(new_n964), .B2(new_n773), .ZN(new_n965));
  AOI21_X1  g779(.A(G953), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n217), .A2(G900), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT124), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n956), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n217), .B1(G227), .B2(G900), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n674), .A2(new_n539), .A3(new_n584), .A4(new_n796), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n971), .A2(new_n769), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n676), .A2(new_n808), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT62), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n676), .A2(KEYINPUT62), .A3(new_n808), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n771), .A2(new_n777), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n955), .B1(new_n978), .B2(G953), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n969), .A2(new_n970), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n970), .B1(new_n969), .B2(new_n979), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n980), .A2(new_n981), .ZN(G72));
  INV_X1    g796(.A(new_n947), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n963), .A2(new_n983), .A3(new_n965), .ZN(new_n984));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  AOI21_X1  g800(.A(new_n515), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n987), .A2(new_n906), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n771), .A2(new_n977), .A3(new_n777), .A4(new_n983), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n986), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT126), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n513), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n989), .A2(KEYINPUT126), .A3(new_n986), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n992), .A2(new_n474), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n528), .B1(new_n474), .B2(new_n513), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n996), .A2(new_n986), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n831), .A2(KEYINPUT127), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(KEYINPUT127), .B1(new_n831), .B2(new_n997), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n988), .B(new_n995), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(G57));
endmodule


