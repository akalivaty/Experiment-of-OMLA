//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n644,
    new_n645, new_n646, new_n649, new_n651, new_n652, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT64), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(KEYINPUT68), .A3(G137), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n466), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n466), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n473), .B(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT67), .B1(new_n467), .B2(new_n468), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n462), .A2(new_n479), .A3(new_n463), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n478), .A2(new_n480), .A3(G125), .ZN(new_n481));
  NAND2_X1  g056(.A1(G113), .A2(G2104), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n466), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n477), .A2(new_n483), .ZN(G160));
  NAND2_X1  g059(.A1(new_n464), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT72), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(new_n466), .B2(G112), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n462), .A2(new_n463), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT70), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n466), .B1(new_n462), .B2(new_n463), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  AND3_X1   g070(.A1(new_n495), .A2(KEYINPUT71), .A3(G124), .ZN(new_n496));
  AOI21_X1  g071(.A(KEYINPUT71), .B1(new_n495), .B2(G124), .ZN(new_n497));
  OAI221_X1 g072(.A(new_n485), .B1(new_n487), .B2(new_n488), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  XOR2_X1   g073(.A(new_n498), .B(KEYINPUT73), .Z(G162));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n478), .A2(new_n480), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n466), .A2(G114), .ZN(new_n505));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT74), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g082(.A1(G102), .A2(G2105), .ZN(new_n508));
  INV_X1    g083(.A(G114), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G2105), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT74), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n508), .A2(new_n510), .A3(new_n511), .A4(G2104), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  NOR3_X1   g088(.A1(new_n503), .A2(new_n500), .A3(G2105), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n492), .A2(G126), .B1(new_n489), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n504), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(G164));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT75), .B1(new_n519), .B2(KEYINPUT6), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT75), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(new_n522), .A3(G651), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n520), .A2(new_n523), .B1(KEYINPUT6), .B2(new_n519), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT76), .ZN(new_n525));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n526), .B2(KEYINPUT5), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT5), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(KEYINPUT76), .A3(G543), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n527), .A2(new_n529), .B1(KEYINPUT5), .B2(new_n526), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n524), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G50), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n518), .A2(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT77), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n530), .A2(G62), .ZN(new_n537));
  NAND2_X1  g112(.A1(G75), .A2(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n519), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n535), .A2(new_n536), .A3(new_n540), .ZN(new_n541));
  OAI21_X1  g116(.A(KEYINPUT77), .B1(new_n534), .B2(new_n539), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(G166));
  AND2_X1   g118(.A1(G63), .A2(G651), .ZN(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(KEYINPUT7), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n545), .A2(KEYINPUT7), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n530), .A2(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n524), .A2(new_n530), .A3(G89), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n524), .A2(G51), .A3(G543), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT78), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n548), .A2(new_n549), .A3(new_n550), .A4(KEYINPUT78), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(G168));
  INV_X1    g130(.A(G90), .ZN(new_n556));
  INV_X1    g131(.A(G52), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n556), .A2(new_n531), .B1(new_n532), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n530), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(new_n519), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n558), .A2(new_n560), .ZN(G171));
  INV_X1    g136(.A(G81), .ZN(new_n562));
  INV_X1    g137(.A(G43), .ZN(new_n563));
  OAI22_X1  g138(.A1(new_n562), .A2(new_n531), .B1(new_n532), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n530), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n565), .A2(new_n519), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT79), .ZN(G153));
  NAND4_X1  g145(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND4_X1  g148(.A1(G319), .A2(G483), .A3(G661), .A4(new_n573), .ZN(G188));
  AND2_X1   g149(.A1(new_n524), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G53), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(KEYINPUT80), .B2(KEYINPUT9), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n575), .B(new_n577), .C1(KEYINPUT80), .C2(KEYINPUT9), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT80), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT9), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n579), .B(new_n580), .C1(new_n532), .C2(new_n576), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n530), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G91), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n583), .A2(new_n519), .B1(new_n531), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G299));
  INV_X1    g162(.A(G171), .ZN(G301));
  INV_X1    g163(.A(G168), .ZN(G286));
  INV_X1    g164(.A(G166), .ZN(G303));
  AND2_X1   g165(.A1(new_n524), .A2(new_n530), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G87), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n575), .A2(G49), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G288));
  NAND2_X1  g170(.A1(new_n526), .A2(KEYINPUT5), .ZN(new_n596));
  AND3_X1   g171(.A1(new_n528), .A2(KEYINPUT76), .A3(G543), .ZN(new_n597));
  AOI21_X1  g172(.A(KEYINPUT76), .B1(new_n528), .B2(G543), .ZN(new_n598));
  OAI211_X1 g173(.A(G61), .B(new_n596), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n530), .A2(KEYINPUT81), .A3(G61), .ZN(new_n602));
  NAND2_X1  g177(.A1(G73), .A2(G543), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G651), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT82), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n604), .A2(KEYINPUT82), .A3(G651), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n524), .A2(new_n530), .A3(G86), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT83), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  AND3_X1   g186(.A1(new_n607), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n524), .A2(G48), .A3(G543), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(G305));
  NAND2_X1  g189(.A1(new_n530), .A2(G60), .ZN(new_n615));
  INV_X1    g190(.A(G72), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(new_n526), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT84), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n519), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n618), .B2(new_n617), .ZN(new_n620));
  AOI22_X1  g195(.A1(G47), .A2(new_n575), .B1(new_n591), .B2(G85), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(G290));
  NAND2_X1  g197(.A1(G301), .A2(G868), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n575), .A2(KEYINPUT86), .ZN(new_n624));
  INV_X1    g199(.A(G54), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT86), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n625), .B1(new_n532), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(KEYINPUT87), .B(G66), .Z(new_n629));
  AOI22_X1  g204(.A1(new_n530), .A2(new_n629), .B1(G79), .B2(G543), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n630), .A2(new_n519), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT85), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n591), .A2(new_n633), .A3(G92), .ZN(new_n634));
  INV_X1    g209(.A(G92), .ZN(new_n635));
  OAI21_X1  g210(.A(KEYINPUT85), .B1(new_n531), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(KEYINPUT10), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n634), .A2(KEYINPUT10), .A3(new_n636), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n623), .B1(new_n641), .B2(G868), .ZN(G284));
  OAI21_X1  g217(.A(new_n623), .B1(new_n641), .B2(G868), .ZN(G321));
  INV_X1    g218(.A(G868), .ZN(new_n644));
  NOR2_X1   g219(.A1(G286), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n586), .B(KEYINPUT88), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n645), .B1(new_n646), .B2(new_n644), .ZN(G297));
  XOR2_X1   g222(.A(G297), .B(KEYINPUT89), .Z(G280));
  INV_X1    g223(.A(G559), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n641), .B1(new_n649), .B2(G860), .ZN(G148));
  NAND2_X1  g225(.A1(new_n641), .A2(new_n649), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(G868), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(G868), .B2(new_n568), .ZN(G323));
  XNOR2_X1  g228(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g229(.A1(new_n478), .A2(new_n480), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(new_n475), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT12), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT13), .ZN(new_n658));
  INV_X1    g233(.A(G2100), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n495), .A2(G123), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n464), .A2(G135), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n466), .A2(G111), .ZN(new_n664));
  OAI21_X1  g239(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n662), .B(new_n663), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(G2096), .Z(new_n667));
  NAND3_X1  g242(.A1(new_n660), .A2(new_n661), .A3(new_n667), .ZN(G156));
  INV_X1    g243(.A(KEYINPUT14), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2427), .B(G2438), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2430), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT15), .B(G2435), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n669), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n673), .B1(new_n672), .B2(new_n671), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2451), .B(G2454), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT16), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1341), .B(G1348), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n674), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2443), .B(G2446), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n681), .A2(new_n682), .A3(G14), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT90), .ZN(G401));
  XOR2_X1   g259(.A(G2072), .B(G2078), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT91), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT17), .ZN(new_n687));
  XNOR2_X1  g262(.A(G2067), .B(G2678), .ZN(new_n688));
  XNOR2_X1  g263(.A(G2084), .B(G2090), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(new_n686), .B2(new_n688), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(new_n687), .B2(new_n688), .ZN(new_n692));
  INV_X1    g267(.A(new_n688), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n693), .A2(new_n689), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n686), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT18), .ZN(new_n696));
  NOR3_X1   g271(.A1(new_n690), .A2(new_n692), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G2096), .B(G2100), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(G227));
  XOR2_X1   g274(.A(G1971), .B(G1976), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT19), .ZN(new_n701));
  XOR2_X1   g276(.A(G1956), .B(G2474), .Z(new_n702));
  XOR2_X1   g277(.A(G1961), .B(G1966), .Z(new_n703));
  AND2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT92), .B(KEYINPUT20), .Z(new_n706));
  XOR2_X1   g281(.A(new_n705), .B(new_n706), .Z(new_n707));
  NOR2_X1   g282(.A1(new_n702), .A2(new_n703), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n701), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT93), .ZN(new_n710));
  NOR3_X1   g285(.A1(new_n701), .A2(new_n704), .A3(new_n708), .ZN(new_n711));
  NOR3_X1   g286(.A1(new_n707), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(G1991), .B(G1996), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(G1981), .B(G1986), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(G229));
  MUX2_X1   g294(.A(G6), .B(G305), .S(G16), .Z(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT32), .B(G1981), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  MUX2_X1   g297(.A(G23), .B(G288), .S(G16), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT33), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1976), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n720), .A2(new_n721), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G22), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G166), .B2(new_n727), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(G1971), .Z(new_n730));
  NAND4_X1  g305(.A1(new_n722), .A2(new_n725), .A3(new_n726), .A4(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(KEYINPUT34), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(KEYINPUT34), .ZN(new_n733));
  NOR2_X1   g308(.A1(G25), .A2(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n495), .A2(G119), .ZN(new_n735));
  OAI21_X1  g310(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n736));
  INV_X1    g311(.A(G107), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(G2105), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G131), .B2(new_n464), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n734), .B1(new_n741), .B2(G29), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT35), .B(G1991), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT94), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n742), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n727), .A2(G24), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(KEYINPUT95), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(KEYINPUT95), .ZN(new_n748));
  INV_X1    g323(.A(G290), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n747), .B(new_n748), .C1(new_n749), .C2(new_n727), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n745), .B(KEYINPUT96), .C1(G1986), .C2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G1986), .B2(new_n750), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n732), .A2(new_n733), .A3(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT36), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n475), .A2(G105), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT101), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n495), .A2(G129), .ZN(new_n760));
  NAND3_X1  g335(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT26), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  AOI22_X1  g339(.A1(G141), .A2(new_n464), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n759), .A2(new_n760), .A3(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT102), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  MUX2_X1   g345(.A(G32), .B(new_n770), .S(G29), .Z(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT27), .Z(new_n772));
  AND2_X1   g347(.A1(new_n772), .A2(G1996), .ZN(new_n773));
  NOR2_X1   g348(.A1(G16), .A2(G19), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n568), .B2(G16), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT97), .Z(new_n776));
  INV_X1    g351(.A(G1341), .ZN(new_n777));
  INV_X1    g352(.A(G2072), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT25), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n464), .A2(G139), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n655), .A2(G127), .ZN(new_n782));
  NAND2_X1  g357(.A1(G115), .A2(G2104), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n466), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT100), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n780), .B(new_n781), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(G29), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n789), .B2(G33), .ZN(new_n791));
  OAI22_X1  g366(.A1(new_n776), .A2(new_n777), .B1(new_n778), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n777), .B2(new_n776), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT24), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n789), .B1(new_n794), .B2(G34), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n794), .B2(G34), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G160), .B2(G29), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(G2084), .Z(new_n798));
  NAND2_X1  g373(.A1(new_n727), .A2(G5), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G171), .B2(new_n727), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n798), .B1(G1961), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT98), .B(KEYINPUT28), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n789), .A2(G26), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n495), .A2(G128), .ZN(new_n805));
  OAI21_X1  g380(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n806));
  INV_X1    g381(.A(G116), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(G2105), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G140), .B2(new_n464), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n805), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n804), .B1(new_n810), .B2(G29), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT99), .B(G2067), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT30), .B(G28), .ZN(new_n814));
  OR2_X1    g389(.A1(KEYINPUT31), .A2(G11), .ZN(new_n815));
  NAND2_X1  g390(.A1(KEYINPUT31), .A2(G11), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n814), .A2(new_n789), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n666), .B2(new_n789), .ZN(new_n818));
  NOR2_X1   g393(.A1(G164), .A2(new_n789), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G27), .B2(new_n789), .ZN(new_n820));
  INV_X1    g395(.A(G2078), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n818), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n800), .A2(G1961), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n813), .A2(new_n822), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(G4), .A2(G16), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(new_n641), .B2(G16), .ZN(new_n827));
  AOI211_X1 g402(.A(new_n801), .B(new_n825), .C1(G1348), .C2(new_n827), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n827), .A2(G1348), .ZN(new_n829));
  NOR2_X1   g404(.A1(G16), .A2(G21), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(G168), .B2(G16), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT103), .B(G1966), .Z(new_n832));
  XOR2_X1   g407(.A(new_n831), .B(new_n832), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n727), .A2(G20), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT23), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n586), .B2(new_n727), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G1956), .ZN(new_n837));
  AOI211_X1 g412(.A(new_n833), .B(new_n837), .C1(new_n778), .C2(new_n791), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n793), .A2(new_n828), .A3(new_n829), .A4(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n772), .A2(G1996), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n789), .A2(G35), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(G162), .B2(new_n789), .ZN(new_n842));
  XNOR2_X1  g417(.A(KEYINPUT29), .B(G2090), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NOR4_X1   g419(.A1(new_n773), .A2(new_n839), .A3(new_n840), .A4(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n755), .A2(new_n756), .A3(new_n845), .ZN(G150));
  INV_X1    g421(.A(G150), .ZN(G311));
  XNOR2_X1  g422(.A(KEYINPUT105), .B(G860), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n640), .A2(new_n649), .ZN(new_n850));
  XNOR2_X1  g425(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n575), .A2(G55), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n591), .A2(G93), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n853), .B(new_n854), .C1(new_n519), .C2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n567), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n852), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n849), .B1(new_n860), .B2(KEYINPUT39), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(KEYINPUT39), .B2(new_n860), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n856), .A2(new_n849), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT37), .Z(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(G145));
  XNOR2_X1  g440(.A(new_n770), .B(G164), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n786), .A2(new_n787), .A3(new_n810), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n810), .B1(new_n786), .B2(new_n787), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n495), .A2(G130), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT106), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n464), .A2(G142), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n875));
  INV_X1    g450(.A(G118), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n875), .B1(new_n876), .B2(G2105), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n868), .B(new_n869), .C1(new_n872), .C2(new_n878), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n872), .A2(new_n877), .A3(new_n874), .ZN(new_n880));
  INV_X1    g455(.A(new_n869), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n880), .B1(new_n881), .B2(new_n867), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n866), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n770), .B(new_n516), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n879), .A2(new_n882), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n740), .B(KEYINPUT107), .Z(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n657), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT108), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n883), .A2(new_n886), .A3(new_n889), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(G162), .A2(new_n666), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(G162), .A2(new_n666), .ZN(new_n897));
  OAI22_X1  g472(.A1(new_n896), .A2(new_n897), .B1(new_n483), .B2(new_n477), .ZN(new_n898));
  INV_X1    g473(.A(new_n897), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n899), .A2(G160), .A3(new_n895), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n894), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n901), .A2(new_n892), .A3(new_n891), .A4(new_n893), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g482(.A1(new_n856), .A2(new_n644), .ZN(new_n908));
  XNOR2_X1  g483(.A(G166), .B(G288), .ZN(new_n909));
  NAND2_X1  g484(.A1(G305), .A2(new_n749), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n612), .A2(new_n613), .A3(G290), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n909), .B1(new_n911), .B2(new_n910), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n914), .B(KEYINPUT42), .Z(new_n915));
  NAND2_X1  g490(.A1(new_n640), .A2(G299), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n638), .A2(new_n586), .A3(new_n639), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT41), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n916), .A2(new_n920), .A3(new_n917), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n921), .A3(KEYINPUT109), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n921), .A2(KEYINPUT109), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n651), .B(new_n858), .ZN(new_n925));
  MUX2_X1   g500(.A(new_n918), .B(new_n924), .S(new_n925), .Z(new_n926));
  XNOR2_X1  g501(.A(new_n915), .B(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n908), .B1(new_n927), .B2(new_n644), .ZN(G295));
  OAI21_X1  g503(.A(new_n908), .B1(new_n927), .B2(new_n644), .ZN(G331));
  INV_X1    g504(.A(KEYINPUT110), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n931));
  XNOR2_X1  g506(.A(G168), .B(G171), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n932), .A2(new_n857), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n857), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n922), .A2(new_n923), .A3(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n918), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n936), .A2(new_n938), .A3(new_n914), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n936), .A2(new_n938), .ZN(new_n941));
  INV_X1    g516(.A(new_n914), .ZN(new_n942));
  AOI21_X1  g517(.A(G37), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n931), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n919), .A2(new_n921), .B1(new_n933), .B2(new_n934), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n945), .A2(new_n937), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n904), .B1(new_n946), .B2(new_n914), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT43), .B1(new_n947), .B2(new_n939), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n930), .B1(new_n944), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n941), .A2(new_n942), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n936), .A2(new_n938), .A3(new_n914), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n950), .A2(new_n951), .A3(new_n904), .A4(new_n952), .ZN(new_n953));
  AND4_X1   g528(.A1(new_n930), .A2(new_n948), .A3(new_n953), .A4(KEYINPUT44), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n951), .B1(new_n943), .B2(new_n952), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n947), .A2(new_n939), .A3(KEYINPUT43), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI22_X1  g532(.A1(new_n949), .A2(new_n954), .B1(KEYINPUT44), .B2(new_n957), .ZN(G397));
  INV_X1    g533(.A(KEYINPUT51), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n553), .A2(G8), .A3(new_n554), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT123), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n960), .B(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT50), .ZN(new_n963));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n516), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n963), .B1(new_n516), .B2(new_n964), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n481), .A2(new_n482), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(G2105), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n968), .A2(G40), .A3(new_n476), .A4(new_n472), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n965), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  XOR2_X1   g545(.A(KEYINPUT118), .B(G2084), .Z(new_n971));
  INV_X1    g546(.A(G40), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n477), .A2(new_n483), .A3(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n516), .A2(new_n964), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n492), .A2(G126), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n489), .A2(new_n514), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n513), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(G1384), .B1(new_n980), .B2(new_n504), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n973), .B(new_n976), .C1(new_n981), .C2(KEYINPUT45), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n970), .A2(new_n971), .B1(new_n982), .B2(new_n832), .ZN(new_n983));
  INV_X1    g558(.A(G8), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n959), .B(new_n962), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT51), .B1(new_n983), .B2(new_n962), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n960), .B(KEYINPUT123), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n982), .A2(new_n832), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n966), .A2(new_n969), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n516), .A2(new_n963), .A3(new_n964), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(new_n990), .A3(new_n971), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n987), .B1(new_n992), .B2(G8), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n985), .B(KEYINPUT62), .C1(new_n986), .C2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT124), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n959), .B1(new_n992), .B2(new_n987), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n983), .A2(new_n984), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n997), .B1(new_n998), .B2(new_n987), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n999), .A2(KEYINPUT124), .A3(KEYINPUT62), .A4(new_n985), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1981), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n613), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n607), .A2(new_n608), .A3(new_n611), .A4(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n603), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(new_n599), .B2(new_n600), .ZN(new_n1008));
  AOI211_X1 g583(.A(new_n606), .B(new_n519), .C1(new_n1008), .C2(new_n602), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT82), .B1(new_n604), .B2(G651), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1011), .A2(KEYINPUT115), .A3(new_n611), .A4(new_n1003), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1006), .A2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT116), .B(G86), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n591), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1011), .A2(new_n613), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(G1981), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n1013), .A2(KEYINPUT49), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT49), .B1(new_n1013), .B2(new_n1017), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n502), .A2(new_n503), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n964), .B1(new_n1020), .B2(new_n979), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n969), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(new_n984), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n1018), .A2(new_n1019), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1976), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1023), .B1(new_n1026), .B2(G288), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT52), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT52), .B1(G288), .B2(new_n1026), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1028), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1021), .A2(KEYINPUT50), .ZN(new_n1032));
  INV_X1    g607(.A(G2090), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1032), .A2(new_n1033), .A3(new_n973), .A4(new_n990), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT114), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n989), .A2(new_n1036), .A3(new_n1033), .A4(new_n990), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1021), .A2(new_n974), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n516), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(new_n973), .A3(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g615(.A(KEYINPUT113), .B(G1971), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1035), .A2(new_n1037), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n541), .A2(G8), .A3(new_n542), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n541), .A2(KEYINPUT55), .A3(G8), .A4(new_n542), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1043), .A2(G8), .A3(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1032), .A2(new_n973), .A3(new_n990), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT117), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1032), .A2(new_n1052), .A3(new_n973), .A4(new_n990), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1033), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n984), .B1(new_n1054), .B2(new_n1042), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1049), .B1(new_n1055), .B2(new_n1048), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1025), .A2(new_n1031), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n1040), .B2(G2078), .ZN(new_n1059));
  INV_X1    g634(.A(G1961), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1050), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n821), .A2(KEYINPUT53), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n982), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(G171), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n985), .B1(new_n986), .B2(new_n993), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT62), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1001), .A2(new_n1057), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT125), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT125), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1001), .A2(new_n1057), .A3(new_n1073), .A4(new_n1070), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n998), .A2(G168), .ZN(new_n1076));
  NOR4_X1   g651(.A1(new_n1025), .A2(new_n1056), .A3(new_n1031), .A4(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT119), .B1(new_n1077), .B2(KEYINPUT63), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT63), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1019), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1013), .A2(KEYINPUT49), .A3(new_n1017), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(new_n1023), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1031), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1048), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1054), .A2(new_n1042), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1085), .B1(new_n1086), .B2(new_n984), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1083), .A2(new_n1084), .A3(new_n1049), .A4(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1079), .B(new_n1080), .C1(new_n1088), .C2(new_n1076), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1049), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1090), .A2(new_n1076), .A3(new_n1080), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1043), .A2(G8), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1085), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1091), .A2(new_n1083), .A3(new_n1084), .A4(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1078), .A2(new_n1089), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1083), .A2(new_n1090), .A3(new_n1084), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1097));
  NOR2_X1   g672(.A1(G288), .A2(G1976), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1097), .A2(new_n1098), .B1(new_n1006), .B2(new_n1012), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1096), .B1(new_n1099), .B2(new_n1024), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1040), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT56), .B(G2072), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT120), .B(G1956), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1101), .A2(new_n1102), .B1(new_n1050), .B2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n586), .B(KEYINPUT57), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G2067), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1022), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G1348), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1050), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n640), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1107), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT58), .B(G1341), .ZN(new_n1115));
  OAI22_X1  g690(.A1(new_n1040), .A2(G1996), .B1(new_n1022), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n568), .ZN(new_n1117));
  XOR2_X1   g692(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1118));
  XNOR2_X1  g693(.A(new_n1117), .B(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT61), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1106), .A2(new_n1120), .A3(new_n1113), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1120), .B1(new_n1106), .B2(new_n1113), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1119), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1111), .A2(new_n1109), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT60), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n641), .B1(new_n1126), .B2(KEYINPUT122), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1128), .B(new_n640), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1126), .A2(KEYINPUT122), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1130), .A2(new_n1131), .B1(new_n1125), .B2(new_n1124), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1114), .B1(new_n1123), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1066), .ZN(new_n1134));
  XNOR2_X1  g709(.A(G171), .B(KEYINPUT54), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1135), .B1(new_n1040), .B2(new_n1064), .ZN(new_n1136));
  OAI22_X1  g711(.A1(new_n1134), .A2(new_n1135), .B1(new_n1062), .B2(new_n1136), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1088), .A2(new_n1068), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1100), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1075), .A2(new_n1095), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n810), .A2(G2067), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n805), .A2(new_n1108), .A3(new_n809), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1143), .B1(new_n770), .B2(G1996), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1038), .A2(new_n969), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n1145), .B(KEYINPUT112), .Z(new_n1146));
  OR2_X1    g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1145), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1148), .A2(G1996), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n1149), .A2(new_n770), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n740), .B(new_n744), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1147), .B(new_n1150), .C1(new_n1146), .C2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g727(.A(G290), .B(G1986), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1152), .B1(new_n1145), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1140), .A2(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1149), .B(KEYINPUT46), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n770), .A2(new_n1143), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1156), .B1(new_n1146), .B2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(KEYINPUT47), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1148), .A2(G290), .A3(G1986), .ZN(new_n1160));
  XOR2_X1   g735(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1161));
  XNOR2_X1  g736(.A(new_n1160), .B(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1159), .B1(new_n1152), .B2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1147), .A2(new_n744), .A3(new_n741), .A4(new_n1150), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1146), .B1(new_n1164), .B2(new_n1142), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1165), .A2(KEYINPUT126), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1165), .A2(KEYINPUT126), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1163), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1155), .A2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g744(.A(G319), .ZN(new_n1171));
  NOR3_X1   g745(.A1(G401), .A2(new_n1171), .A3(G227), .ZN(new_n1172));
  AND2_X1   g746(.A1(new_n718), .A2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g747(.A(new_n906), .B(new_n1173), .C1(new_n955), .C2(new_n956), .ZN(G225));
  INV_X1    g748(.A(G225), .ZN(G308));
endmodule


