

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U551 ( .A1(G2105), .A2(G2104), .ZN(n866) );
  INV_X1 U552 ( .A(n713), .ZN(n697) );
  AND2_X2 U553 ( .A1(n525), .A2(G2104), .ZN(n860) );
  OR2_X1 U554 ( .A1(KEYINPUT33), .A2(n736), .ZN(n745) );
  NAND2_X1 U555 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U556 ( .A1(n745), .A2(n744), .ZN(n518) );
  AND2_X1 U557 ( .A1(n713), .A2(G1341), .ZN(n519) );
  AND2_X1 U558 ( .A1(n697), .A2(G1996), .ZN(n680) );
  OR2_X1 U559 ( .A1(n681), .A2(n519), .ZN(n682) );
  INV_X1 U560 ( .A(KEYINPUT99), .ZN(n720) );
  XNOR2_X1 U561 ( .A(n721), .B(n720), .ZN(n722) );
  NAND2_X1 U562 ( .A1(G160), .A2(G40), .ZN(n740) );
  NOR2_X1 U563 ( .A1(G543), .A2(G651), .ZN(n624) );
  NOR2_X1 U564 ( .A1(n529), .A2(n528), .ZN(G160) );
  INV_X1 U565 ( .A(G2105), .ZN(n525) );
  NAND2_X1 U566 ( .A1(G101), .A2(n860), .ZN(n520) );
  XOR2_X1 U567 ( .A(KEYINPUT23), .B(n520), .Z(n523) );
  NAND2_X1 U568 ( .A1(G113), .A2(n866), .ZN(n521) );
  XOR2_X1 U569 ( .A(KEYINPUT65), .B(n521), .Z(n522) );
  NAND2_X1 U570 ( .A1(n523), .A2(n522), .ZN(n529) );
  NOR2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  XOR2_X2 U572 ( .A(KEYINPUT17), .B(n524), .Z(n861) );
  NAND2_X1 U573 ( .A1(G137), .A2(n861), .ZN(n527) );
  NOR2_X1 U574 ( .A1(G2104), .A2(n525), .ZN(n864) );
  NAND2_X1 U575 ( .A1(G125), .A2(n864), .ZN(n526) );
  NAND2_X1 U576 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U577 ( .A(KEYINPUT66), .B(G651), .Z(n538) );
  NOR2_X1 U578 ( .A1(G543), .A2(n538), .ZN(n530) );
  XOR2_X1 U579 ( .A(KEYINPUT1), .B(n530), .Z(n638) );
  NAND2_X1 U580 ( .A1(G63), .A2(n638), .ZN(n533) );
  XOR2_X1 U581 ( .A(KEYINPUT0), .B(G543), .Z(n633) );
  NOR2_X1 U582 ( .A1(n633), .A2(G651), .ZN(n531) );
  XNOR2_X1 U583 ( .A(KEYINPUT64), .B(n531), .ZN(n634) );
  NAND2_X1 U584 ( .A1(G51), .A2(n634), .ZN(n532) );
  NAND2_X1 U585 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U586 ( .A(KEYINPUT6), .B(n534), .ZN(n543) );
  XOR2_X1 U587 ( .A(KEYINPUT4), .B(KEYINPUT70), .Z(n536) );
  NAND2_X1 U588 ( .A1(G89), .A2(n624), .ZN(n535) );
  XNOR2_X1 U589 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U590 ( .A(KEYINPUT69), .B(n537), .ZN(n540) );
  NOR2_X1 U591 ( .A1(n633), .A2(n538), .ZN(n627) );
  NAND2_X1 U592 ( .A1(n627), .A2(G76), .ZN(n539) );
  NAND2_X1 U593 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U594 ( .A(n541), .B(KEYINPUT5), .Z(n542) );
  NOR2_X1 U595 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U596 ( .A(KEYINPUT7), .B(n544), .Z(n545) );
  XOR2_X1 U597 ( .A(KEYINPUT71), .B(n545), .Z(G168) );
  XOR2_X1 U598 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U599 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U600 ( .A1(G65), .A2(n638), .ZN(n547) );
  NAND2_X1 U601 ( .A1(G53), .A2(n634), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n547), .A2(n546), .ZN(n551) );
  NAND2_X1 U603 ( .A1(G91), .A2(n624), .ZN(n549) );
  NAND2_X1 U604 ( .A1(G78), .A2(n627), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U606 ( .A1(n551), .A2(n550), .ZN(n691) );
  INV_X1 U607 ( .A(n691), .ZN(G299) );
  INV_X1 U608 ( .A(G57), .ZN(G237) );
  INV_X1 U609 ( .A(G132), .ZN(G219) );
  INV_X1 U610 ( .A(G82), .ZN(G220) );
  NAND2_X1 U611 ( .A1(G7), .A2(G661), .ZN(n552) );
  XNOR2_X1 U612 ( .A(n552), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U613 ( .A(G223), .ZN(n809) );
  NAND2_X1 U614 ( .A1(n809), .A2(G567), .ZN(n553) );
  XOR2_X1 U615 ( .A(KEYINPUT11), .B(n553), .Z(G234) );
  NAND2_X1 U616 ( .A1(n638), .A2(G56), .ZN(n554) );
  XOR2_X1 U617 ( .A(KEYINPUT14), .B(n554), .Z(n560) );
  NAND2_X1 U618 ( .A1(n624), .A2(G81), .ZN(n555) );
  XNOR2_X1 U619 ( .A(n555), .B(KEYINPUT12), .ZN(n557) );
  NAND2_X1 U620 ( .A1(G68), .A2(n627), .ZN(n556) );
  NAND2_X1 U621 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U622 ( .A(KEYINPUT13), .B(n558), .Z(n559) );
  NOR2_X1 U623 ( .A1(n560), .A2(n559), .ZN(n562) );
  NAND2_X1 U624 ( .A1(G43), .A2(n634), .ZN(n561) );
  NAND2_X1 U625 ( .A1(n562), .A2(n561), .ZN(n902) );
  INV_X1 U626 ( .A(G860), .ZN(n583) );
  OR2_X1 U627 ( .A1(n902), .A2(n583), .ZN(G153) );
  NAND2_X1 U628 ( .A1(G64), .A2(n638), .ZN(n564) );
  NAND2_X1 U629 ( .A1(G52), .A2(n634), .ZN(n563) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n569) );
  NAND2_X1 U631 ( .A1(G90), .A2(n624), .ZN(n566) );
  NAND2_X1 U632 ( .A1(G77), .A2(n627), .ZN(n565) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U634 ( .A(KEYINPUT9), .B(n567), .Z(n568) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(KEYINPUT68), .B(n570), .ZN(G171) );
  INV_X1 U637 ( .A(G171), .ZN(G301) );
  NAND2_X1 U638 ( .A1(G301), .A2(G868), .ZN(n579) );
  NAND2_X1 U639 ( .A1(n627), .A2(G79), .ZN(n572) );
  NAND2_X1 U640 ( .A1(G54), .A2(n634), .ZN(n571) );
  NAND2_X1 U641 ( .A1(n572), .A2(n571), .ZN(n576) );
  NAND2_X1 U642 ( .A1(G66), .A2(n638), .ZN(n574) );
  NAND2_X1 U643 ( .A1(G92), .A2(n624), .ZN(n573) );
  NAND2_X1 U644 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U645 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U646 ( .A(n577), .B(KEYINPUT15), .ZN(n913) );
  INV_X1 U647 ( .A(G868), .ZN(n580) );
  NAND2_X1 U648 ( .A1(n913), .A2(n580), .ZN(n578) );
  NAND2_X1 U649 ( .A1(n579), .A2(n578), .ZN(G284) );
  NOR2_X1 U650 ( .A1(G286), .A2(n580), .ZN(n582) );
  NOR2_X1 U651 ( .A1(G868), .A2(G299), .ZN(n581) );
  NOR2_X1 U652 ( .A1(n582), .A2(n581), .ZN(G297) );
  NAND2_X1 U653 ( .A1(G559), .A2(n583), .ZN(n584) );
  XNOR2_X1 U654 ( .A(KEYINPUT72), .B(n584), .ZN(n585) );
  INV_X1 U655 ( .A(n913), .ZN(n601) );
  NAND2_X1 U656 ( .A1(n585), .A2(n601), .ZN(n586) );
  XNOR2_X1 U657 ( .A(KEYINPUT16), .B(n586), .ZN(G148) );
  NOR2_X1 U658 ( .A1(G868), .A2(n902), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n601), .A2(G868), .ZN(n587) );
  NOR2_X1 U660 ( .A1(G559), .A2(n587), .ZN(n588) );
  NOR2_X1 U661 ( .A1(n589), .A2(n588), .ZN(G282) );
  XOR2_X1 U662 ( .A(KEYINPUT73), .B(KEYINPUT18), .Z(n591) );
  NAND2_X1 U663 ( .A1(G123), .A2(n864), .ZN(n590) );
  XNOR2_X1 U664 ( .A(n591), .B(n590), .ZN(n598) );
  NAND2_X1 U665 ( .A1(G135), .A2(n861), .ZN(n593) );
  NAND2_X1 U666 ( .A1(G111), .A2(n866), .ZN(n592) );
  NAND2_X1 U667 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n860), .A2(G99), .ZN(n594) );
  XOR2_X1 U669 ( .A(KEYINPUT74), .B(n594), .Z(n595) );
  NOR2_X1 U670 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n598), .A2(n597), .ZN(n994) );
  XOR2_X1 U672 ( .A(n994), .B(G2096), .Z(n600) );
  XNOR2_X1 U673 ( .A(G2100), .B(KEYINPUT75), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(G156) );
  NAND2_X1 U675 ( .A1(n601), .A2(G559), .ZN(n650) );
  XNOR2_X1 U676 ( .A(n902), .B(n650), .ZN(n602) );
  NOR2_X1 U677 ( .A1(n602), .A2(G860), .ZN(n610) );
  NAND2_X1 U678 ( .A1(G80), .A2(n627), .ZN(n603) );
  XNOR2_X1 U679 ( .A(n603), .B(KEYINPUT76), .ZN(n605) );
  NAND2_X1 U680 ( .A1(n638), .A2(G67), .ZN(n604) );
  NAND2_X1 U681 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U682 ( .A1(n624), .A2(G93), .ZN(n607) );
  NAND2_X1 U683 ( .A1(G55), .A2(n634), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U685 ( .A1(n609), .A2(n608), .ZN(n653) );
  XNOR2_X1 U686 ( .A(n610), .B(n653), .ZN(G145) );
  NAND2_X1 U687 ( .A1(G88), .A2(n624), .ZN(n612) );
  NAND2_X1 U688 ( .A1(G75), .A2(n627), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U690 ( .A1(G62), .A2(n638), .ZN(n614) );
  NAND2_X1 U691 ( .A1(G50), .A2(n634), .ZN(n613) );
  NAND2_X1 U692 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U693 ( .A1(n616), .A2(n615), .ZN(G166) );
  NAND2_X1 U694 ( .A1(G47), .A2(n634), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n638), .A2(G60), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U697 ( .A(KEYINPUT67), .B(n619), .ZN(n623) );
  NAND2_X1 U698 ( .A1(G85), .A2(n624), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G72), .A2(n627), .ZN(n620) );
  AND2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U701 ( .A1(n623), .A2(n622), .ZN(G290) );
  NAND2_X1 U702 ( .A1(G61), .A2(n638), .ZN(n626) );
  NAND2_X1 U703 ( .A1(G86), .A2(n624), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U705 ( .A1(n627), .A2(G73), .ZN(n628) );
  XOR2_X1 U706 ( .A(KEYINPUT2), .B(n628), .Z(n629) );
  NOR2_X1 U707 ( .A1(n630), .A2(n629), .ZN(n632) );
  NAND2_X1 U708 ( .A1(G48), .A2(n634), .ZN(n631) );
  NAND2_X1 U709 ( .A1(n632), .A2(n631), .ZN(G305) );
  NAND2_X1 U710 ( .A1(n633), .A2(G87), .ZN(n636) );
  NAND2_X1 U711 ( .A1(G49), .A2(n634), .ZN(n635) );
  NAND2_X1 U712 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U714 ( .A1(G651), .A2(G74), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n640), .A2(n639), .ZN(G288) );
  XNOR2_X1 U716 ( .A(G166), .B(G290), .ZN(n641) );
  XNOR2_X1 U717 ( .A(n641), .B(G305), .ZN(n647) );
  XOR2_X1 U718 ( .A(KEYINPUT19), .B(KEYINPUT78), .Z(n642) );
  XNOR2_X1 U719 ( .A(G288), .B(n642), .ZN(n643) );
  XNOR2_X1 U720 ( .A(KEYINPUT77), .B(n643), .ZN(n645) );
  XNOR2_X1 U721 ( .A(n902), .B(KEYINPUT79), .ZN(n644) );
  XNOR2_X1 U722 ( .A(n645), .B(n644), .ZN(n646) );
  XOR2_X1 U723 ( .A(n647), .B(n646), .Z(n649) );
  XNOR2_X1 U724 ( .A(n691), .B(n653), .ZN(n648) );
  XNOR2_X1 U725 ( .A(n649), .B(n648), .ZN(n880) );
  XNOR2_X1 U726 ( .A(n880), .B(KEYINPUT80), .ZN(n651) );
  XNOR2_X1 U727 ( .A(n651), .B(n650), .ZN(n652) );
  NAND2_X1 U728 ( .A1(n652), .A2(G868), .ZN(n655) );
  OR2_X1 U729 ( .A1(n653), .A2(G868), .ZN(n654) );
  NAND2_X1 U730 ( .A1(n655), .A2(n654), .ZN(G295) );
  NAND2_X1 U731 ( .A1(G2078), .A2(G2084), .ZN(n656) );
  XOR2_X1 U732 ( .A(KEYINPUT20), .B(n656), .Z(n657) );
  NAND2_X1 U733 ( .A1(G2090), .A2(n657), .ZN(n658) );
  XNOR2_X1 U734 ( .A(KEYINPUT21), .B(n658), .ZN(n659) );
  NAND2_X1 U735 ( .A1(n659), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U736 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U737 ( .A1(G220), .A2(G219), .ZN(n660) );
  XOR2_X1 U738 ( .A(KEYINPUT22), .B(n660), .Z(n661) );
  NOR2_X1 U739 ( .A1(G218), .A2(n661), .ZN(n662) );
  NAND2_X1 U740 ( .A1(G96), .A2(n662), .ZN(n815) );
  NAND2_X1 U741 ( .A1(n815), .A2(G2106), .ZN(n666) );
  NAND2_X1 U742 ( .A1(G69), .A2(G120), .ZN(n663) );
  NOR2_X1 U743 ( .A1(G237), .A2(n663), .ZN(n664) );
  NAND2_X1 U744 ( .A1(G108), .A2(n664), .ZN(n816) );
  NAND2_X1 U745 ( .A1(n816), .A2(G567), .ZN(n665) );
  NAND2_X1 U746 ( .A1(n666), .A2(n665), .ZN(n817) );
  NAND2_X1 U747 ( .A1(G483), .A2(G661), .ZN(n667) );
  NOR2_X1 U748 ( .A1(n817), .A2(n667), .ZN(n813) );
  NAND2_X1 U749 ( .A1(n813), .A2(G36), .ZN(G176) );
  NAND2_X1 U750 ( .A1(n861), .A2(G138), .ZN(n670) );
  NAND2_X1 U751 ( .A1(G102), .A2(n860), .ZN(n668) );
  XOR2_X1 U752 ( .A(KEYINPUT81), .B(n668), .Z(n669) );
  NAND2_X1 U753 ( .A1(n670), .A2(n669), .ZN(n674) );
  NAND2_X1 U754 ( .A1(G126), .A2(n864), .ZN(n672) );
  NAND2_X1 U755 ( .A1(G114), .A2(n866), .ZN(n671) );
  NAND2_X1 U756 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U757 ( .A1(n674), .A2(n673), .ZN(G164) );
  INV_X1 U758 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U759 ( .A(KEYINPUT93), .B(n740), .ZN(n675) );
  NOR2_X1 U760 ( .A1(G164), .A2(G1384), .ZN(n741) );
  NAND2_X2 U761 ( .A1(n675), .A2(n741), .ZN(n713) );
  NAND2_X1 U762 ( .A1(n697), .A2(G2072), .ZN(n676) );
  XNOR2_X1 U763 ( .A(n676), .B(KEYINPUT27), .ZN(n678) );
  AND2_X1 U764 ( .A1(G1956), .A2(n713), .ZN(n677) );
  NOR2_X1 U765 ( .A1(n678), .A2(n677), .ZN(n690) );
  NOR2_X1 U766 ( .A1(n691), .A2(n690), .ZN(n679) );
  XOR2_X1 U767 ( .A(n679), .B(KEYINPUT28), .Z(n695) );
  XNOR2_X1 U768 ( .A(n680), .B(KEYINPUT26), .ZN(n681) );
  NOR2_X1 U769 ( .A1(n902), .A2(n682), .ZN(n686) );
  NAND2_X1 U770 ( .A1(G1348), .A2(n713), .ZN(n684) );
  NAND2_X1 U771 ( .A1(G2067), .A2(n697), .ZN(n683) );
  NAND2_X1 U772 ( .A1(n684), .A2(n683), .ZN(n687) );
  NOR2_X1 U773 ( .A1(n913), .A2(n687), .ZN(n685) );
  OR2_X1 U774 ( .A1(n686), .A2(n685), .ZN(n689) );
  NAND2_X1 U775 ( .A1(n913), .A2(n687), .ZN(n688) );
  NAND2_X1 U776 ( .A1(n689), .A2(n688), .ZN(n693) );
  NAND2_X1 U777 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U778 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U779 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U780 ( .A(KEYINPUT29), .B(n696), .Z(n701) );
  XOR2_X1 U781 ( .A(G1961), .B(KEYINPUT95), .Z(n956) );
  NAND2_X1 U782 ( .A1(n956), .A2(n713), .ZN(n699) );
  XOR2_X1 U783 ( .A(G2078), .B(KEYINPUT25), .Z(n942) );
  NAND2_X1 U784 ( .A1(n697), .A2(n942), .ZN(n698) );
  NAND2_X1 U785 ( .A1(n699), .A2(n698), .ZN(n707) );
  OR2_X1 U786 ( .A1(n707), .A2(G301), .ZN(n700) );
  NAND2_X1 U787 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U788 ( .A(n702), .B(KEYINPUT96), .ZN(n712) );
  NAND2_X1 U789 ( .A1(G8), .A2(n713), .ZN(n753) );
  NOR2_X1 U790 ( .A1(G1966), .A2(n753), .ZN(n727) );
  NOR2_X1 U791 ( .A1(G2084), .A2(n713), .ZN(n724) );
  NOR2_X1 U792 ( .A1(n727), .A2(n724), .ZN(n703) );
  NAND2_X1 U793 ( .A1(G8), .A2(n703), .ZN(n704) );
  XNOR2_X1 U794 ( .A(KEYINPUT30), .B(n704), .ZN(n705) );
  NOR2_X1 U795 ( .A1(G168), .A2(n705), .ZN(n706) );
  XNOR2_X1 U796 ( .A(n706), .B(KEYINPUT97), .ZN(n709) );
  NAND2_X1 U797 ( .A1(G301), .A2(n707), .ZN(n708) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U799 ( .A(KEYINPUT31), .B(n710), .ZN(n711) );
  NAND2_X1 U800 ( .A1(n712), .A2(n711), .ZN(n728) );
  NAND2_X1 U801 ( .A1(n728), .A2(G286), .ZN(n719) );
  NOR2_X1 U802 ( .A1(G1971), .A2(n753), .ZN(n715) );
  NOR2_X1 U803 ( .A1(G2090), .A2(n713), .ZN(n714) );
  NOR2_X1 U804 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U805 ( .A(n716), .B(KEYINPUT98), .ZN(n717) );
  NAND2_X1 U806 ( .A1(n717), .A2(G303), .ZN(n718) );
  NAND2_X1 U807 ( .A1(n719), .A2(n718), .ZN(n721) );
  NAND2_X1 U808 ( .A1(n722), .A2(G8), .ZN(n723) );
  XNOR2_X1 U809 ( .A(n723), .B(KEYINPUT32), .ZN(n731) );
  NAND2_X1 U810 ( .A1(G8), .A2(n724), .ZN(n725) );
  XOR2_X1 U811 ( .A(KEYINPUT94), .B(n725), .Z(n726) );
  NOR2_X1 U812 ( .A1(n727), .A2(n726), .ZN(n729) );
  NAND2_X1 U813 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U814 ( .A1(n731), .A2(n730), .ZN(n748) );
  NOR2_X1 U815 ( .A1(G1976), .A2(G288), .ZN(n903) );
  NOR2_X1 U816 ( .A1(G1971), .A2(G303), .ZN(n919) );
  NOR2_X1 U817 ( .A1(n903), .A2(n919), .ZN(n732) );
  NAND2_X1 U818 ( .A1(n748), .A2(n732), .ZN(n735) );
  INV_X1 U819 ( .A(n753), .ZN(n733) );
  NAND2_X1 U820 ( .A1(G1976), .A2(G288), .ZN(n916) );
  AND2_X1 U821 ( .A1(n733), .A2(n916), .ZN(n734) );
  AND2_X1 U822 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U823 ( .A1(n903), .A2(KEYINPUT33), .ZN(n737) );
  NOR2_X1 U824 ( .A1(n737), .A2(n753), .ZN(n739) );
  XOR2_X1 U825 ( .A(G1981), .B(G305), .Z(n909) );
  INV_X1 U826 ( .A(n909), .ZN(n738) );
  NOR2_X1 U827 ( .A1(n739), .A2(n738), .ZN(n743) );
  XNOR2_X1 U828 ( .A(G1986), .B(G290), .ZN(n925) );
  NOR2_X1 U829 ( .A1(n741), .A2(n740), .ZN(n804) );
  NAND2_X1 U830 ( .A1(n925), .A2(n804), .ZN(n742) );
  XNOR2_X1 U831 ( .A(n742), .B(KEYINPUT82), .ZN(n756) );
  AND2_X1 U832 ( .A1(n743), .A2(n756), .ZN(n744) );
  NOR2_X1 U833 ( .A1(G2090), .A2(G303), .ZN(n746) );
  NAND2_X1 U834 ( .A1(G8), .A2(n746), .ZN(n747) );
  NAND2_X1 U835 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U836 ( .A(n749), .B(KEYINPUT100), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n750), .A2(n753), .ZN(n755) );
  NOR2_X1 U838 ( .A1(G1981), .A2(G305), .ZN(n751) );
  XOR2_X1 U839 ( .A(n751), .B(KEYINPUT24), .Z(n752) );
  OR2_X1 U840 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U841 ( .A1(n755), .A2(n754), .ZN(n757) );
  NAND2_X1 U842 ( .A1(n518), .A2(n758), .ZN(n795) );
  NAND2_X1 U843 ( .A1(G131), .A2(n861), .ZN(n759) );
  XNOR2_X1 U844 ( .A(n759), .B(KEYINPUT88), .ZN(n766) );
  NAND2_X1 U845 ( .A1(G95), .A2(n860), .ZN(n761) );
  NAND2_X1 U846 ( .A1(G119), .A2(n864), .ZN(n760) );
  NAND2_X1 U847 ( .A1(n761), .A2(n760), .ZN(n764) );
  NAND2_X1 U848 ( .A1(G107), .A2(n866), .ZN(n762) );
  XNOR2_X1 U849 ( .A(KEYINPUT87), .B(n762), .ZN(n763) );
  NOR2_X1 U850 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U851 ( .A1(n766), .A2(n765), .ZN(n857) );
  NAND2_X1 U852 ( .A1(G1991), .A2(n857), .ZN(n767) );
  XOR2_X1 U853 ( .A(KEYINPUT89), .B(n767), .Z(n778) );
  NAND2_X1 U854 ( .A1(G117), .A2(n866), .ZN(n768) );
  XOR2_X1 U855 ( .A(KEYINPUT90), .B(n768), .Z(n771) );
  NAND2_X1 U856 ( .A1(n860), .A2(G105), .ZN(n769) );
  XOR2_X1 U857 ( .A(KEYINPUT38), .B(n769), .Z(n770) );
  NOR2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n773) );
  NAND2_X1 U859 ( .A1(n864), .A2(G129), .ZN(n772) );
  NAND2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U861 ( .A(n774), .B(KEYINPUT91), .ZN(n776) );
  NAND2_X1 U862 ( .A1(G141), .A2(n861), .ZN(n775) );
  NAND2_X1 U863 ( .A1(n776), .A2(n775), .ZN(n856) );
  NAND2_X1 U864 ( .A1(G1996), .A2(n856), .ZN(n777) );
  NAND2_X1 U865 ( .A1(n778), .A2(n777), .ZN(n998) );
  NAND2_X1 U866 ( .A1(n998), .A2(n804), .ZN(n779) );
  XNOR2_X1 U867 ( .A(n779), .B(KEYINPUT92), .ZN(n793) );
  XNOR2_X1 U868 ( .A(KEYINPUT37), .B(G2067), .ZN(n802) );
  XNOR2_X1 U869 ( .A(KEYINPUT35), .B(KEYINPUT85), .ZN(n783) );
  NAND2_X1 U870 ( .A1(G128), .A2(n864), .ZN(n781) );
  NAND2_X1 U871 ( .A1(G116), .A2(n866), .ZN(n780) );
  NAND2_X1 U872 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U873 ( .A(n783), .B(n782), .ZN(n790) );
  XNOR2_X1 U874 ( .A(KEYINPUT83), .B(KEYINPUT84), .ZN(n784) );
  XNOR2_X1 U875 ( .A(n784), .B(KEYINPUT34), .ZN(n788) );
  NAND2_X1 U876 ( .A1(G104), .A2(n860), .ZN(n786) );
  NAND2_X1 U877 ( .A1(G140), .A2(n861), .ZN(n785) );
  NAND2_X1 U878 ( .A1(n786), .A2(n785), .ZN(n787) );
  XOR2_X1 U879 ( .A(n788), .B(n787), .Z(n789) );
  NOR2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U881 ( .A(KEYINPUT36), .B(n791), .ZN(n876) );
  NOR2_X1 U882 ( .A1(n802), .A2(n876), .ZN(n997) );
  NAND2_X1 U883 ( .A1(n804), .A2(n997), .ZN(n792) );
  XNOR2_X1 U884 ( .A(KEYINPUT86), .B(n792), .ZN(n800) );
  AND2_X1 U885 ( .A1(n793), .A2(n800), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n807) );
  NOR2_X1 U887 ( .A1(G1996), .A2(n856), .ZN(n1002) );
  NOR2_X1 U888 ( .A1(G1991), .A2(n857), .ZN(n993) );
  NOR2_X1 U889 ( .A1(G1986), .A2(G290), .ZN(n796) );
  NOR2_X1 U890 ( .A1(n993), .A2(n796), .ZN(n797) );
  NOR2_X1 U891 ( .A1(n998), .A2(n797), .ZN(n798) );
  NOR2_X1 U892 ( .A1(n1002), .A2(n798), .ZN(n799) );
  XNOR2_X1 U893 ( .A(n799), .B(KEYINPUT39), .ZN(n801) );
  NAND2_X1 U894 ( .A1(n801), .A2(n800), .ZN(n803) );
  NAND2_X1 U895 ( .A1(n802), .A2(n876), .ZN(n999) );
  NAND2_X1 U896 ( .A1(n803), .A2(n999), .ZN(n805) );
  NAND2_X1 U897 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U898 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U899 ( .A(n808), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U900 ( .A1(G2106), .A2(n809), .ZN(G217) );
  AND2_X1 U901 ( .A1(G15), .A2(G2), .ZN(n810) );
  NAND2_X1 U902 ( .A1(G661), .A2(n810), .ZN(G259) );
  NAND2_X1 U903 ( .A1(G3), .A2(G1), .ZN(n811) );
  XOR2_X1 U904 ( .A(KEYINPUT103), .B(n811), .Z(n812) );
  NAND2_X1 U905 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U906 ( .A(KEYINPUT104), .B(n814), .ZN(G188) );
  INV_X1 U908 ( .A(G120), .ZN(G236) );
  INV_X1 U909 ( .A(G96), .ZN(G221) );
  INV_X1 U910 ( .A(G69), .ZN(G235) );
  NOR2_X1 U911 ( .A1(n816), .A2(n815), .ZN(G325) );
  INV_X1 U912 ( .A(G325), .ZN(G261) );
  INV_X1 U913 ( .A(n817), .ZN(G319) );
  XOR2_X1 U914 ( .A(KEYINPUT41), .B(G1971), .Z(n819) );
  XNOR2_X1 U915 ( .A(G1966), .B(G1956), .ZN(n818) );
  XNOR2_X1 U916 ( .A(n819), .B(n818), .ZN(n820) );
  XOR2_X1 U917 ( .A(n820), .B(KEYINPUT107), .Z(n822) );
  XNOR2_X1 U918 ( .A(G1996), .B(G1991), .ZN(n821) );
  XNOR2_X1 U919 ( .A(n822), .B(n821), .ZN(n826) );
  XOR2_X1 U920 ( .A(G1976), .B(G1981), .Z(n824) );
  XNOR2_X1 U921 ( .A(G1986), .B(G1961), .ZN(n823) );
  XNOR2_X1 U922 ( .A(n824), .B(n823), .ZN(n825) );
  XOR2_X1 U923 ( .A(n826), .B(n825), .Z(n828) );
  XNOR2_X1 U924 ( .A(KEYINPUT106), .B(G2474), .ZN(n827) );
  XNOR2_X1 U925 ( .A(n828), .B(n827), .ZN(G229) );
  XOR2_X1 U926 ( .A(G2678), .B(G2084), .Z(n830) );
  XNOR2_X1 U927 ( .A(G2078), .B(G2072), .ZN(n829) );
  XNOR2_X1 U928 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U929 ( .A(n831), .B(G2100), .Z(n833) );
  XNOR2_X1 U930 ( .A(G2067), .B(G2090), .ZN(n832) );
  XNOR2_X1 U931 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U932 ( .A(G2096), .B(KEYINPUT105), .Z(n835) );
  XNOR2_X1 U933 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n834) );
  XNOR2_X1 U934 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U935 ( .A(n837), .B(n836), .Z(G227) );
  NAND2_X1 U936 ( .A1(n864), .A2(G124), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n838), .B(KEYINPUT44), .ZN(n840) );
  NAND2_X1 U938 ( .A1(G112), .A2(n866), .ZN(n839) );
  NAND2_X1 U939 ( .A1(n840), .A2(n839), .ZN(n844) );
  NAND2_X1 U940 ( .A1(G100), .A2(n860), .ZN(n842) );
  NAND2_X1 U941 ( .A1(G136), .A2(n861), .ZN(n841) );
  NAND2_X1 U942 ( .A1(n842), .A2(n841), .ZN(n843) );
  NOR2_X1 U943 ( .A1(n844), .A2(n843), .ZN(G162) );
  XOR2_X1 U944 ( .A(KEYINPUT110), .B(KEYINPUT48), .Z(n855) );
  NAND2_X1 U945 ( .A1(G130), .A2(n864), .ZN(n846) );
  NAND2_X1 U946 ( .A1(G118), .A2(n866), .ZN(n845) );
  NAND2_X1 U947 ( .A1(n846), .A2(n845), .ZN(n852) );
  NAND2_X1 U948 ( .A1(G106), .A2(n860), .ZN(n848) );
  NAND2_X1 U949 ( .A1(G142), .A2(n861), .ZN(n847) );
  NAND2_X1 U950 ( .A1(n848), .A2(n847), .ZN(n849) );
  XOR2_X1 U951 ( .A(KEYINPUT45), .B(n849), .Z(n850) );
  XNOR2_X1 U952 ( .A(KEYINPUT108), .B(n850), .ZN(n851) );
  NOR2_X1 U953 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n853), .B(KEYINPUT46), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n875) );
  XNOR2_X1 U956 ( .A(G160), .B(n856), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n994), .B(n859), .ZN(n873) );
  NAND2_X1 U959 ( .A1(G103), .A2(n860), .ZN(n863) );
  NAND2_X1 U960 ( .A1(G139), .A2(n861), .ZN(n862) );
  NAND2_X1 U961 ( .A1(n863), .A2(n862), .ZN(n871) );
  NAND2_X1 U962 ( .A1(n864), .A2(G127), .ZN(n865) );
  XOR2_X1 U963 ( .A(KEYINPUT109), .B(n865), .Z(n868) );
  NAND2_X1 U964 ( .A1(n866), .A2(G115), .ZN(n867) );
  NAND2_X1 U965 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U966 ( .A(KEYINPUT47), .B(n869), .Z(n870) );
  NOR2_X1 U967 ( .A1(n871), .A2(n870), .ZN(n987) );
  XNOR2_X1 U968 ( .A(G164), .B(n987), .ZN(n872) );
  XNOR2_X1 U969 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U970 ( .A(n875), .B(n874), .ZN(n878) );
  XNOR2_X1 U971 ( .A(n876), .B(G162), .ZN(n877) );
  XNOR2_X1 U972 ( .A(n878), .B(n877), .ZN(n879) );
  NOR2_X1 U973 ( .A1(G37), .A2(n879), .ZN(G395) );
  XOR2_X1 U974 ( .A(G286), .B(n880), .Z(n881) );
  XNOR2_X1 U975 ( .A(n913), .B(n881), .ZN(n882) );
  XOR2_X1 U976 ( .A(G171), .B(n882), .Z(n883) );
  NOR2_X1 U977 ( .A1(G37), .A2(n883), .ZN(n884) );
  XOR2_X1 U978 ( .A(KEYINPUT111), .B(n884), .Z(G397) );
  XNOR2_X1 U979 ( .A(G2451), .B(G2427), .ZN(n894) );
  XOR2_X1 U980 ( .A(G2430), .B(G2443), .Z(n886) );
  XNOR2_X1 U981 ( .A(G2435), .B(G2438), .ZN(n885) );
  XNOR2_X1 U982 ( .A(n886), .B(n885), .ZN(n890) );
  XOR2_X1 U983 ( .A(G2454), .B(KEYINPUT101), .Z(n888) );
  XNOR2_X1 U984 ( .A(G1341), .B(G1348), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U986 ( .A(n890), .B(n889), .Z(n892) );
  XNOR2_X1 U987 ( .A(G2446), .B(KEYINPUT102), .ZN(n891) );
  XNOR2_X1 U988 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U989 ( .A(n894), .B(n893), .ZN(n895) );
  NAND2_X1 U990 ( .A1(n895), .A2(G14), .ZN(n901) );
  NAND2_X1 U991 ( .A1(G319), .A2(n901), .ZN(n898) );
  NOR2_X1 U992 ( .A1(G229), .A2(G227), .ZN(n896) );
  XNOR2_X1 U993 ( .A(KEYINPUT49), .B(n896), .ZN(n897) );
  NOR2_X1 U994 ( .A1(n898), .A2(n897), .ZN(n900) );
  NOR2_X1 U995 ( .A1(G395), .A2(G397), .ZN(n899) );
  NAND2_X1 U996 ( .A1(n900), .A2(n899), .ZN(G225) );
  INV_X1 U997 ( .A(G225), .ZN(G308) );
  INV_X1 U998 ( .A(G108), .ZN(G238) );
  INV_X1 U999 ( .A(n901), .ZN(G401) );
  XNOR2_X1 U1000 ( .A(n902), .B(G1341), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(n903), .B(KEYINPUT122), .ZN(n904) );
  NOR2_X1 U1002 ( .A1(n905), .A2(n904), .ZN(n907) );
  NAND2_X1 U1003 ( .A1(G1971), .A2(G303), .ZN(n906) );
  NAND2_X1 U1004 ( .A1(n907), .A2(n906), .ZN(n923) );
  XNOR2_X1 U1005 ( .A(G1966), .B(G168), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n908), .B(KEYINPUT120), .ZN(n910) );
  NAND2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(n912) );
  XOR2_X1 U1008 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n921) );
  XNOR2_X1 U1010 ( .A(n913), .B(G1348), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(G299), .B(G1956), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(n917) );
  NAND2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1015 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1016 ( .A1(n923), .A2(n922), .ZN(n927) );
  XNOR2_X1 U1017 ( .A(G1961), .B(G301), .ZN(n924) );
  NOR2_X1 U1018 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1019 ( .A1(n927), .A2(n926), .ZN(n930) );
  XOR2_X1 U1020 ( .A(G16), .B(KEYINPUT56), .Z(n928) );
  XNOR2_X1 U1021 ( .A(KEYINPUT119), .B(n928), .ZN(n929) );
  NAND2_X1 U1022 ( .A1(n930), .A2(n929), .ZN(n985) );
  XOR2_X1 U1023 ( .A(KEYINPUT117), .B(G34), .Z(n932) );
  XNOR2_X1 U1024 ( .A(G2084), .B(KEYINPUT54), .ZN(n931) );
  XNOR2_X1 U1025 ( .A(n932), .B(n931), .ZN(n950) );
  XNOR2_X1 U1026 ( .A(G2090), .B(G35), .ZN(n933) );
  XNOR2_X1 U1027 ( .A(n933), .B(KEYINPUT114), .ZN(n947) );
  XNOR2_X1 U1028 ( .A(G2067), .B(G26), .ZN(n935) );
  XNOR2_X1 U1029 ( .A(G1991), .B(G25), .ZN(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n941) );
  XOR2_X1 U1031 ( .A(G2072), .B(G33), .Z(n936) );
  NAND2_X1 U1032 ( .A1(n936), .A2(G28), .ZN(n939) );
  XOR2_X1 U1033 ( .A(KEYINPUT115), .B(G1996), .Z(n937) );
  XNOR2_X1 U1034 ( .A(G32), .B(n937), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n944) );
  XNOR2_X1 U1037 ( .A(G27), .B(n942), .ZN(n943) );
  NOR2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1039 ( .A(n945), .B(KEYINPUT53), .ZN(n946) );
  NOR2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1041 ( .A(KEYINPUT116), .B(n948), .Z(n949) );
  NOR2_X1 U1042 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1043 ( .A(KEYINPUT55), .B(n951), .ZN(n953) );
  INV_X1 U1044 ( .A(G29), .ZN(n952) );
  NAND2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1046 ( .A1(n954), .A2(G11), .ZN(n955) );
  XNOR2_X1 U1047 ( .A(KEYINPUT118), .B(n955), .ZN(n983) );
  XOR2_X1 U1048 ( .A(n956), .B(G5), .Z(n967) );
  XNOR2_X1 U1049 ( .A(G1348), .B(KEYINPUT59), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(n957), .B(G4), .ZN(n961) );
  XNOR2_X1 U1051 ( .A(G1341), .B(G19), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(G1981), .B(G6), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n964) );
  XOR2_X1 U1055 ( .A(KEYINPUT123), .B(G1956), .Z(n962) );
  XNOR2_X1 U1056 ( .A(G20), .B(n962), .ZN(n963) );
  NOR2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(KEYINPUT60), .B(n965), .ZN(n966) );
  NAND2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n978) );
  XOR2_X1 U1060 ( .A(G1966), .B(G21), .Z(n976) );
  XOR2_X1 U1061 ( .A(G1971), .B(G22), .Z(n970) );
  XOR2_X1 U1062 ( .A(G23), .B(KEYINPUT124), .Z(n968) );
  XNOR2_X1 U1063 ( .A(n968), .B(G1976), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n973) );
  XOR2_X1 U1065 ( .A(KEYINPUT125), .B(G1986), .Z(n971) );
  XNOR2_X1 U1066 ( .A(G24), .B(n971), .ZN(n972) );
  NOR2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(n974), .B(KEYINPUT58), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1071 ( .A(KEYINPUT61), .B(n979), .Z(n980) );
  NOR2_X1 U1072 ( .A1(G16), .A2(n980), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(n981), .B(KEYINPUT126), .ZN(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(n986), .B(KEYINPUT127), .ZN(n1016) );
  XNOR2_X1 U1077 ( .A(G2072), .B(n987), .ZN(n990) );
  XOR2_X1 U1078 ( .A(G164), .B(G2078), .Z(n988) );
  XNOR2_X1 U1079 ( .A(KEYINPUT113), .B(n988), .ZN(n989) );
  NAND2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(n991), .B(KEYINPUT50), .ZN(n1010) );
  XOR2_X1 U1082 ( .A(G160), .B(G2084), .Z(n992) );
  NOR2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n995) );
  NAND2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n1008) );
  INV_X1 U1086 ( .A(n998), .ZN(n1000) );
  NAND2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1006) );
  XOR2_X1 U1088 ( .A(G2090), .B(G162), .Z(n1001) );
  NOR2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1090 ( .A(KEYINPUT112), .B(n1003), .Z(n1004) );
  XOR2_X1 U1091 ( .A(KEYINPUT51), .B(n1004), .Z(n1005) );
  NOR2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1094 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1095 ( .A(KEYINPUT52), .B(n1011), .ZN(n1013) );
  INV_X1 U1096 ( .A(KEYINPUT55), .ZN(n1012) );
  NAND2_X1 U1097 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1098 ( .A1(n1014), .A2(G29), .ZN(n1015) );
  NAND2_X1 U1099 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1100 ( .A(KEYINPUT62), .B(n1017), .Z(G311) );
  INV_X1 U1101 ( .A(G311), .ZN(G150) );
endmodule

