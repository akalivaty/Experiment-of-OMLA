//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n561, new_n563, new_n564, new_n565, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n616, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT64), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  XNOR2_X1  g032(.A(KEYINPUT3), .B(G2104), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n458), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n460), .A2(G101), .A3(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n463));
  OR2_X1    g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n463), .ZN(new_n465));
  OR2_X1    g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n464), .A2(new_n465), .B1(new_n468), .B2(G137), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n461), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(G160));
  AOI21_X1  g046(.A(new_n460), .B1(new_n466), .B2(new_n467), .ZN(new_n472));
  OR2_X1    g047(.A1(new_n472), .A2(KEYINPUT66), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(KEYINPUT66), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  MUX2_X1   g052(.A(G100), .B(G112), .S(G2105), .Z(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2104), .ZN(new_n479));
  XOR2_X1   g054(.A(new_n479), .B(KEYINPUT67), .Z(new_n480));
  AOI211_X1 g055(.A(new_n477), .B(new_n480), .C1(G136), .C2(new_n468), .ZN(G162));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n468), .A2(new_n482), .A3(G138), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n483), .B(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n486));
  AND2_X1   g061(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n487));
  NOR2_X1   g062(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n488));
  OAI211_X1 g063(.A(G138), .B(new_n460), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT68), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n458), .A2(new_n491), .A3(G138), .A4(new_n460), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n486), .B1(new_n493), .B2(KEYINPUT4), .ZN(new_n494));
  AOI211_X1 g069(.A(KEYINPUT69), .B(new_n482), .C1(new_n490), .C2(new_n492), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n485), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n472), .A2(G126), .ZN(new_n497));
  MUX2_X1   g072(.A(G102), .B(G114), .S(G2105), .Z(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G2104), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n496), .A2(KEYINPUT71), .A3(new_n501), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n509), .A2(new_n511), .B1(new_n508), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n513), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(KEYINPUT72), .A3(G651), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n515), .A2(new_n517), .B1(KEYINPUT6), .B2(new_n514), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(G543), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(G88), .A2(new_n520), .B1(new_n522), .B2(G50), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n512), .A2(KEYINPUT74), .A3(G62), .ZN(new_n524));
  NAND2_X1  g099(.A1(G75), .A2(G543), .ZN(new_n525));
  XOR2_X1   g100(.A(new_n525), .B(KEYINPUT75), .Z(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(KEYINPUT74), .B1(new_n512), .B2(G62), .ZN(new_n528));
  OAI21_X1  g103(.A(G651), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n523), .A2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NAND2_X1  g106(.A1(new_n520), .A2(G89), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n522), .A2(G51), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n512), .A2(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n532), .A2(new_n533), .A3(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n509), .A2(new_n511), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n508), .A2(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G64), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n541), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n514), .B1(new_n546), .B2(KEYINPUT76), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n547), .B1(KEYINPUT76), .B2(new_n546), .ZN(new_n548));
  AOI22_X1  g123(.A1(G90), .A2(new_n520), .B1(new_n522), .B2(G52), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  INV_X1    g127(.A(G43), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n519), .A2(new_n552), .B1(new_n521), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT77), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(new_n514), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  XOR2_X1   g137(.A(KEYINPUT78), .B(KEYINPUT8), .Z(new_n563));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n565), .ZN(G188));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n544), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n569), .B2(KEYINPUT79), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(KEYINPUT79), .B2(new_n569), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(KEYINPUT80), .ZN(new_n572));
  INV_X1    g147(.A(G53), .ZN(new_n573));
  OR3_X1    g148(.A1(new_n521), .A2(KEYINPUT9), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT9), .B1(new_n521), .B2(new_n573), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n574), .A2(new_n575), .B1(G91), .B2(new_n520), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n571), .A2(KEYINPUT80), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G299));
  NAND2_X1  g155(.A1(new_n520), .A2(G87), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n522), .A2(G49), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT81), .ZN(G288));
  NAND2_X1  g160(.A1(new_n512), .A2(G61), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT82), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n514), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n520), .A2(G86), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n522), .A2(G48), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G305));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n519), .A2(new_n594), .B1(new_n521), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n514), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g174(.A(new_n599), .B(KEYINPUT83), .Z(G290));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NOR2_X1   g176(.A1(G301), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n520), .A2(G92), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(KEYINPUT10), .Z(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n544), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G651), .B1(new_n522), .B2(G54), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n602), .B1(new_n610), .B2(new_n601), .ZN(G284));
  AOI21_X1  g186(.A(new_n602), .B1(new_n610), .B2(new_n601), .ZN(G321));
  NOR2_X1   g187(.A1(G286), .A2(new_n601), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(new_n579), .B2(new_n601), .ZN(G297));
  AOI21_X1  g189(.A(new_n613), .B1(new_n579), .B2(new_n601), .ZN(G280));
  XNOR2_X1  g190(.A(KEYINPUT84), .B(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n610), .B1(G860), .B2(new_n616), .ZN(G148));
  NAND2_X1  g192(.A1(new_n610), .A2(new_n616), .ZN(new_n618));
  MUX2_X1   g193(.A(new_n558), .B(new_n618), .S(G868), .Z(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n468), .A2(G2104), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT12), .Z(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT13), .Z(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n624), .A2(G2100), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(G2100), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n468), .A2(G135), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  AND2_X1   g203(.A1(new_n628), .A2(KEYINPUT85), .ZN(new_n629));
  OAI22_X1  g204(.A1(new_n628), .A2(KEYINPUT85), .B1(G111), .B2(new_n460), .ZN(new_n630));
  INV_X1    g205(.A(G123), .ZN(new_n631));
  OAI221_X1 g206(.A(new_n627), .B1(new_n629), .B2(new_n630), .C1(new_n475), .C2(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(G2096), .Z(new_n633));
  NAND3_X1  g208(.A1(new_n625), .A2(new_n626), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT86), .ZN(G156));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT89), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2427), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT88), .B(G2438), .Z(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT90), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT87), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2451), .B(G2454), .Z(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT91), .ZN(new_n653));
  INV_X1    g228(.A(G14), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n654), .B1(new_n650), .B2(new_n651), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT17), .Z(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n660), .B2(new_n658), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT92), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n663), .A2(new_n660), .A3(new_n658), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT18), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n664), .A2(new_n660), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n669), .B1(new_n659), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT93), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G2096), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2100), .ZN(G227));
  XOR2_X1   g250(.A(G1971), .B(G1976), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT20), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  OR3_X1    g259(.A1(new_n677), .A2(new_n680), .A3(new_n683), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(new_n691), .ZN(G229));
  NOR2_X1   g267(.A1(G29), .A2(G35), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(G162), .B2(G29), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT29), .Z(new_n695));
  INV_X1    g270(.A(G2090), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G21), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G168), .B2(new_n698), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n700), .A2(G1966), .ZN(new_n701));
  OR2_X1    g276(.A1(KEYINPUT30), .A2(G28), .ZN(new_n702));
  NAND2_X1  g277(.A1(KEYINPUT30), .A2(G28), .ZN(new_n703));
  AOI21_X1  g278(.A(G29), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT31), .B(G11), .Z(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  INV_X1    g282(.A(G34), .ZN(new_n708));
  AOI21_X1  g283(.A(G29), .B1(new_n708), .B2(KEYINPUT24), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n709), .A2(KEYINPUT99), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(KEYINPUT99), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(KEYINPUT24), .B2(new_n708), .ZN(new_n712));
  OAI22_X1  g287(.A1(new_n470), .A2(new_n707), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G2084), .ZN(new_n714));
  OAI221_X1 g289(.A(new_n706), .B1(new_n713), .B2(new_n714), .C1(new_n707), .C2(new_n632), .ZN(new_n715));
  AOI211_X1 g290(.A(new_n701), .B(new_n715), .C1(new_n714), .C2(new_n713), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n707), .A2(G32), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT100), .B(KEYINPUT26), .ZN(new_n718));
  NAND3_X1  g293(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n468), .A2(G141), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n718), .A2(new_n719), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n460), .A2(G105), .A3(G2104), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n720), .A2(new_n721), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n476), .B2(G129), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n717), .B1(new_n725), .B2(new_n707), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT27), .B(G1996), .Z(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT101), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n726), .B(new_n728), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT25), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n468), .A2(G139), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n458), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n731), .B(new_n732), .C1(new_n733), .C2(new_n460), .ZN(new_n734));
  MUX2_X1   g309(.A(G33), .B(new_n734), .S(G29), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G2072), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n729), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n707), .A2(G26), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT28), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n476), .A2(G128), .ZN(new_n740));
  MUX2_X1   g315(.A(G104), .B(G116), .S(G2105), .Z(new_n741));
  AOI22_X1  g316(.A1(G140), .A2(new_n468), .B1(new_n741), .B2(G2104), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n739), .B1(new_n743), .B2(G29), .ZN(new_n744));
  INV_X1    g319(.A(G2067), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G1966), .B2(new_n700), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n697), .A2(new_n716), .A3(new_n737), .A4(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n695), .A2(new_n696), .ZN(new_n749));
  NOR2_X1   g324(.A1(G4), .A2(G16), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n610), .B2(G16), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1348), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n748), .A2(new_n749), .A3(new_n752), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT102), .B(KEYINPUT23), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n698), .A2(G20), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n579), .B2(new_n698), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT103), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G1956), .ZN(new_n759));
  NOR2_X1   g334(.A1(G16), .A2(G19), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n559), .B2(G16), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(G1341), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n698), .A2(G5), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G171), .B2(new_n698), .ZN(new_n764));
  INV_X1    g339(.A(G1961), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n753), .A2(new_n759), .A3(new_n762), .A4(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n758), .A2(G1956), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n707), .A2(G27), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G164), .B2(new_n707), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2078), .ZN(new_n771));
  NOR3_X1   g346(.A1(new_n767), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  MUX2_X1   g347(.A(G6), .B(G305), .S(G16), .Z(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT95), .Z(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT32), .B(G1981), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  MUX2_X1   g352(.A(G23), .B(new_n584), .S(G16), .Z(new_n778));
  XOR2_X1   g353(.A(KEYINPUT33), .B(G1976), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT97), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT96), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n778), .B(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G16), .A2(G22), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G166), .B2(G16), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n782), .B1(G1971), .B2(new_n784), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(G1971), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n774), .A2(new_n776), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n777), .A2(new_n785), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n788), .A2(KEYINPUT34), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n476), .A2(G119), .ZN(new_n790));
  MUX2_X1   g365(.A(G95), .B(G107), .S(G2105), .Z(new_n791));
  AOI22_X1  g366(.A1(G131), .A2(new_n468), .B1(new_n791), .B2(G2104), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  MUX2_X1   g368(.A(G25), .B(new_n793), .S(G29), .Z(new_n794));
  XOR2_X1   g369(.A(KEYINPUT35), .B(G1991), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(G1986), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n698), .A2(G24), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n798), .A2(KEYINPUT94), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n798), .A2(KEYINPUT94), .ZN(new_n800));
  AOI211_X1 g375(.A(new_n799), .B(new_n800), .C1(G290), .C2(G16), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n796), .B1(new_n797), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n797), .B2(new_n801), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n788), .B2(KEYINPUT34), .ZN(new_n804));
  OAI22_X1  g379(.A1(new_n789), .A2(new_n804), .B1(KEYINPUT98), .B2(KEYINPUT36), .ZN(new_n805));
  AND2_X1   g380(.A1(KEYINPUT98), .A2(KEYINPUT36), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n772), .A2(new_n807), .A3(new_n808), .ZN(G150));
  INV_X1    g384(.A(G150), .ZN(G311));
  NAND2_X1  g385(.A1(new_n610), .A2(G559), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  AOI22_X1  g388(.A1(G93), .A2(new_n520), .B1(new_n522), .B2(G55), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n514), .B2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT105), .ZN(new_n817));
  MUX2_X1   g392(.A(new_n816), .B(new_n817), .S(new_n558), .Z(new_n818));
  XOR2_X1   g393(.A(new_n813), .B(new_n818), .Z(new_n819));
  INV_X1    g394(.A(KEYINPUT39), .ZN(new_n820));
  AOI21_X1  g395(.A(G860), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n820), .B2(new_n819), .ZN(new_n822));
  INV_X1    g397(.A(new_n817), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G860), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT37), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n822), .A2(new_n825), .ZN(G145));
  XNOR2_X1  g401(.A(new_n793), .B(new_n622), .ZN(new_n827));
  MUX2_X1   g402(.A(G106), .B(G118), .S(G2105), .Z(new_n828));
  AOI22_X1  g403(.A1(G142), .A2(new_n468), .B1(new_n828), .B2(G2104), .ZN(new_n829));
  INV_X1    g404(.A(G130), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n475), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n827), .B(new_n831), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n500), .B(KEYINPUT107), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n496), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n743), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n832), .B(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n725), .B(new_n734), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n632), .B(new_n470), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT106), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(G162), .Z(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(G37), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n843), .B2(new_n839), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g421(.A1(new_n823), .A2(G868), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n818), .B(new_n618), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n579), .B(new_n610), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(KEYINPUT41), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n850), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(G290), .B(new_n584), .ZN(new_n853));
  XOR2_X1   g428(.A(G303), .B(G305), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT42), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n855), .B1(KEYINPUT108), .B2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n852), .B(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n856), .A2(KEYINPUT108), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n858), .B(new_n859), .Z(new_n860));
  AOI21_X1  g435(.A(new_n847), .B1(new_n860), .B2(G868), .ZN(G295));
  AOI21_X1  g436(.A(new_n847), .B1(new_n860), .B2(G868), .ZN(G331));
  INV_X1    g437(.A(KEYINPUT44), .ZN(new_n863));
  XNOR2_X1  g438(.A(G301), .B(G168), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n818), .B(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n851), .A2(new_n865), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n865), .A2(new_n849), .ZN(new_n867));
  AOI21_X1  g442(.A(KEYINPUT109), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(new_n855), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(G37), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n868), .B2(new_n855), .ZN(new_n872));
  OAI21_X1  g447(.A(KEYINPUT43), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n866), .A2(new_n867), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT109), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n855), .ZN(new_n877));
  AOI21_X1  g452(.A(G37), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n879), .A3(new_n869), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n863), .B1(new_n873), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT110), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n873), .A2(new_n880), .A3(new_n863), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n884), .ZN(new_n886));
  OAI21_X1  g461(.A(KEYINPUT110), .B1(new_n886), .B2(new_n881), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(G397));
  XNOR2_X1  g463(.A(KEYINPUT111), .B(G1384), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n834), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT112), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n889), .B1(new_n496), .B2(new_n833), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT112), .ZN(new_n895));
  AOI21_X1  g470(.A(KEYINPUT45), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  XOR2_X1   g471(.A(KEYINPUT113), .B(G40), .Z(new_n897));
  NOR2_X1   g472(.A1(new_n470), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n743), .B(new_n745), .ZN(new_n900));
  OR3_X1    g475(.A1(new_n899), .A2(KEYINPUT115), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(KEYINPUT115), .B1(new_n899), .B2(new_n900), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n725), .B(G1996), .Z(new_n903));
  NAND3_X1  g478(.A1(new_n896), .A2(new_n903), .A3(new_n898), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n793), .B(new_n795), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n905), .B1(new_n899), .B2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(G290), .B(new_n797), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n899), .A2(new_n908), .ZN(new_n909));
  XOR2_X1   g484(.A(new_n909), .B(KEYINPUT114), .Z(new_n910));
  NOR2_X1   g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(G1384), .B1(new_n496), .B2(new_n833), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n898), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G8), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(KEYINPUT117), .B(G86), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n592), .B1(new_n519), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(G1981), .B1(new_n918), .B2(new_n589), .ZN(new_n919));
  INV_X1    g494(.A(G1981), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n590), .A2(new_n591), .A3(new_n592), .A4(new_n920), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n919), .A2(KEYINPUT49), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT49), .B1(new_n919), .B2(new_n921), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI211_X1 g499(.A(G1976), .B(G288), .C1(new_n916), .C2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n921), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n916), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(G8), .A3(new_n913), .ZN(new_n928));
  INV_X1    g503(.A(G1976), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT52), .B1(G288), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n584), .A2(new_n929), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT116), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n930), .A2(new_n932), .A3(G8), .A4(new_n913), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n928), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT52), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n935), .B1(new_n916), .B2(new_n932), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(G303), .A2(G8), .ZN(new_n939));
  XOR2_X1   g514(.A(new_n939), .B(KEYINPUT55), .Z(new_n940));
  INV_X1    g515(.A(G1384), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n504), .A2(new_n941), .A3(new_n505), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT50), .ZN(new_n943));
  INV_X1    g518(.A(new_n898), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT50), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n944), .B1(new_n912), .B2(new_n945), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n943), .A2(new_n696), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n942), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n944), .B1(new_n894), .B2(KEYINPUT45), .ZN(new_n950));
  AOI21_X1  g525(.A(G1971), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI211_X1 g526(.A(G8), .B(new_n940), .C1(new_n947), .C2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n927), .B1(new_n938), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT119), .ZN(new_n954));
  XNOR2_X1  g529(.A(KEYINPUT118), .B(KEYINPUT63), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n912), .A2(KEYINPUT50), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n496), .A2(KEYINPUT71), .A3(new_n501), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT71), .B1(new_n496), .B2(new_n501), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n957), .A2(new_n958), .A3(G1384), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n956), .B1(new_n959), .B2(KEYINPUT50), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n960), .A2(new_n696), .A3(new_n898), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n950), .B1(new_n959), .B2(KEYINPUT45), .ZN(new_n962));
  INV_X1    g537(.A(G1971), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n915), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n952), .B(new_n937), .C1(new_n965), .C2(new_n940), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n943), .A2(new_n714), .A3(new_n946), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n942), .A2(KEYINPUT45), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n912), .A2(new_n948), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n944), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n967), .B1(new_n971), .B2(G1966), .ZN(new_n972));
  NOR2_X1   g547(.A1(G286), .A2(new_n915), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n954), .B(new_n955), .C1(new_n966), .C2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n940), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n943), .A2(new_n696), .A3(new_n946), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n964), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT120), .B1(new_n978), .B2(G8), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT120), .ZN(new_n980));
  AOI211_X1 g555(.A(new_n980), .B(new_n915), .C1(new_n964), .C2(new_n977), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n976), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n952), .A2(new_n937), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n972), .A2(KEYINPUT63), .A3(new_n973), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n975), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n955), .B1(new_n966), .B2(new_n974), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT119), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n953), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n946), .B1(new_n959), .B2(new_n945), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT122), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1348), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n943), .A2(KEYINPUT122), .A3(new_n946), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n914), .A2(new_n745), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n609), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g573(.A(KEYINPUT121), .B(KEYINPUT57), .Z(new_n999));
  XNOR2_X1  g574(.A(new_n579), .B(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n898), .B1(new_n891), .B2(new_n948), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1001), .B1(new_n948), .B2(new_n942), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT56), .B(G2072), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n960), .A2(new_n898), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n1000), .B(new_n1004), .C1(new_n1005), .C2(G1956), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n998), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1000), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1009));
  AOI21_X1  g584(.A(G1956), .B1(new_n960), .B2(new_n898), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1008), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n996), .A2(new_n609), .A3(new_n997), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT60), .B1(new_n1013), .B2(new_n998), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1011), .A2(new_n1006), .A3(KEYINPUT61), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT58), .B(G1341), .ZN(new_n1016));
  OAI22_X1  g591(.A1(new_n962), .A2(G1996), .B1(new_n914), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT123), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT59), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1017), .A2(new_n559), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1020), .B1(new_n1017), .B2(new_n559), .ZN(new_n1022));
  OAI22_X1  g597(.A1(new_n1021), .A2(new_n1022), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n609), .A2(KEYINPUT60), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n996), .A2(new_n997), .A3(new_n1024), .ZN(new_n1025));
  AND4_X1   g600(.A1(new_n1014), .A2(new_n1015), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT61), .B1(new_n1011), .B2(new_n1006), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT124), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1012), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n993), .A2(new_n765), .A3(new_n995), .ZN(new_n1031));
  INV_X1    g606(.A(G2078), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n971), .A2(KEYINPUT53), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n962), .B2(G2078), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1031), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G171), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT125), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT126), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G160), .A2(G40), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1040), .B1(new_n896), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n894), .A2(KEYINPUT112), .ZN(new_n1043));
  AOI211_X1 g618(.A(new_n892), .B(new_n889), .C1(new_n496), .C2(new_n833), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n948), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1045), .A2(KEYINPUT126), .A3(G40), .A4(G160), .ZN(new_n1046));
  AOI211_X1 g621(.A(new_n1034), .B(G2078), .C1(new_n894), .C2(KEYINPUT45), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1042), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1048), .A2(new_n1031), .A3(new_n1035), .ZN(new_n1049));
  OR2_X1    g624(.A1(new_n1049), .A2(G171), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1036), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1039), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1049), .A2(G171), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1031), .A2(new_n1033), .A3(G301), .A4(new_n1035), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(KEYINPUT54), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1966), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n969), .B1(KEYINPUT45), .B2(new_n942), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1058), .B1(new_n1059), .B2(new_n944), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1060), .A2(G168), .A3(new_n967), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G8), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT51), .ZN(new_n1063));
  AOI21_X1  g638(.A(G168), .B1(new_n1060), .B2(new_n967), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT51), .ZN(new_n1065));
  OAI211_X1 g640(.A(G8), .B(new_n1061), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n966), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1057), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1054), .A2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n990), .B(KEYINPUT127), .C1(new_n1030), .C2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n966), .B1(new_n1039), .B2(new_n1051), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1067), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1073), .A2(KEYINPUT62), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1073), .A2(KEYINPUT62), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1072), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1071), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1012), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1079));
  AOI211_X1 g654(.A(KEYINPUT124), .B(KEYINPUT61), .C1(new_n1011), .C2(new_n1006), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1014), .A2(new_n1015), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1078), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1083), .A2(new_n1054), .A3(new_n1069), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT127), .B1(new_n1084), .B2(new_n990), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n911), .B1(new_n1077), .B2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n899), .A2(G1996), .ZN(new_n1087));
  XNOR2_X1  g662(.A(new_n1087), .B(KEYINPUT46), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n899), .B1(new_n725), .B2(new_n900), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n1090), .B(KEYINPUT47), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n905), .A2(new_n790), .A3(new_n792), .A4(new_n795), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n835), .A2(new_n745), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n899), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n899), .A2(G1986), .A3(G290), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1095), .B(KEYINPUT48), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n907), .A2(new_n1096), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1091), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1086), .A2(new_n1098), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g674(.A1(new_n873), .A2(new_n880), .ZN(new_n1101));
  INV_X1    g675(.A(new_n1101), .ZN(new_n1102));
  INV_X1    g676(.A(G319), .ZN(new_n1103));
  NOR3_X1   g677(.A1(G227), .A2(new_n1103), .A3(G229), .ZN(new_n1104));
  NAND3_X1  g678(.A1(new_n656), .A2(new_n845), .A3(new_n1104), .ZN(new_n1105));
  NOR2_X1   g679(.A1(new_n1102), .A2(new_n1105), .ZN(G308));
  INV_X1    g680(.A(G308), .ZN(G225));
endmodule


