//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n613, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT67), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n466), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT68), .B1(new_n471), .B2(new_n467), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AND2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n478), .A2(new_n479), .A3(G2105), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n470), .B1(new_n472), .B2(new_n480), .ZN(G160));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(new_n463), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n467), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n488));
  INV_X1    g063(.A(G136), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n486), .B(new_n488), .C1(new_n489), .C2(new_n468), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  OAI211_X1 g066(.A(G138), .B(new_n467), .C1(new_n474), .C2(new_n475), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n466), .A2(new_n494), .A3(G138), .A4(new_n467), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT69), .A2(G114), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n499), .A2(G2105), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(G126), .A2(new_n485), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  XNOR2_X1  g081(.A(KEYINPUT5), .B(G543), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n509), .A2(G88), .B1(G50), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n507), .A2(G62), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n514), .B1(KEYINPUT70), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n518), .A2(KEYINPUT70), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(G166));
  AND2_X1   g096(.A1(G63), .A2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n507), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT71), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n507), .A2(new_n525), .A3(new_n522), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n513), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(KEYINPUT73), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(KEYINPUT73), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT7), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n532), .A2(new_n536), .A3(new_n533), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n535), .A2(new_n537), .B1(G89), .B2(new_n509), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n530), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n528), .B1(new_n527), .B2(new_n529), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(G168));
  NAND2_X1  g116(.A1(new_n507), .A2(G64), .ZN(new_n542));
  NAND2_X1  g117(.A1(G77), .A2(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n515), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n544), .A2(KEYINPUT74), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n544), .A2(KEYINPUT74), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n513), .A2(G52), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n507), .A2(new_n508), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR3_X1   g125(.A1(new_n545), .A2(new_n546), .A3(new_n550), .ZN(G171));
  NAND2_X1  g126(.A1(new_n513), .A2(G43), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n553), .B2(new_n549), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n515), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(new_n513), .A2(G53), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n549), .A2(KEYINPUT75), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n507), .A2(new_n508), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(G91), .A3(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n569), .A2(new_n515), .ZN(new_n570));
  AND3_X1   g145(.A1(new_n564), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G299));
  INV_X1    g147(.A(G171), .ZN(G301));
  INV_X1    g148(.A(G168), .ZN(G286));
  INV_X1    g149(.A(G166), .ZN(G303));
  NAND3_X1  g150(.A1(new_n565), .A2(G87), .A3(new_n567), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n507), .A2(G74), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(G49), .B2(new_n513), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(G288));
  NAND2_X1  g154(.A1(new_n507), .A2(G61), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(G48), .B2(new_n513), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n565), .A2(G86), .A3(new_n567), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(new_n513), .A2(G47), .ZN(new_n586));
  INV_X1    g161(.A(G85), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n587), .B2(new_n549), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n515), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n565), .A2(G92), .A3(new_n567), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(KEYINPUT76), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT76), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n565), .A2(new_n596), .A3(G92), .A4(new_n567), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n595), .A2(KEYINPUT10), .A3(new_n597), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(new_n507), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(G651), .B1(G54), .B2(new_n513), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n600), .A2(new_n601), .A3(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n593), .B1(new_n608), .B2(G868), .ZN(G284));
  OAI21_X1  g184(.A(new_n593), .B1(new_n608), .B2(G868), .ZN(G321));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NOR2_X1   g186(.A1(G168), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n613), .B(KEYINPUT77), .C1(G868), .C2(new_n571), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(KEYINPUT77), .B2(new_n613), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT78), .ZN(G297));
  XNOR2_X1  g191(.A(new_n615), .B(KEYINPUT79), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n608), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n608), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n485), .A2(G123), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n467), .A2(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  INV_X1    g201(.A(G135), .ZN(new_n627));
  OAI221_X1 g202(.A(new_n624), .B1(new_n625), .B2(new_n626), .C1(new_n627), .C2(new_n468), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT81), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2096), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT80), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G2100), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n466), .A2(new_n464), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT13), .Z(new_n635));
  NOR2_X1   g210(.A1(new_n631), .A2(G2100), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n630), .B(new_n637), .C1(new_n635), .C2(new_n632), .ZN(G156));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2430), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT82), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(new_n640), .B2(new_n641), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n649), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(new_n653), .A3(G14), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(G401));
  INV_X1    g230(.A(KEYINPUT18), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(KEYINPUT17), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n656), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2100), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n659), .B2(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2096), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n663), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  AND2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT20), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n671), .A2(new_n672), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n670), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n670), .B2(new_n676), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G1981), .ZN(new_n680));
  INV_X1    g255(.A(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT83), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n682), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G229));
  XOR2_X1   g263(.A(KEYINPUT88), .B(G16), .Z(new_n689));
  INV_X1    g264(.A(G20), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT23), .Z(new_n692));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n692), .B1(new_n571), .B2(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT98), .B(G1956), .Z(new_n695));
  XOR2_X1   g270(.A(new_n694), .B(new_n695), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(G21), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G168), .B2(new_n693), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n698), .A2(G1966), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT96), .ZN(new_n700));
  INV_X1    g275(.A(new_n468), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G139), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT93), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT25), .Z(new_n705));
  AOI22_X1  g280(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n703), .B(new_n705), .C1(new_n467), .C2(new_n706), .ZN(new_n707));
  MUX2_X1   g282(.A(G33), .B(new_n707), .S(G29), .Z(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(G2072), .Z(new_n709));
  INV_X1    g284(.A(KEYINPUT24), .ZN(new_n710));
  INV_X1    g285(.A(G34), .ZN(new_n711));
  AOI21_X1  g286(.A(G29), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n710), .B2(new_n711), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(G160), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G2084), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(G32), .ZN(new_n717));
  NAND3_X1  g292(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT26), .Z(new_n719));
  NAND2_X1  g294(.A1(new_n485), .A2(G129), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n464), .A2(G105), .ZN(new_n722));
  INV_X1    g297(.A(G141), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n468), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n717), .B1(new_n725), .B2(new_n714), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT27), .B(G1996), .Z(new_n727));
  OAI211_X1 g302(.A(new_n709), .B(new_n716), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n700), .B1(new_n728), .B2(KEYINPUT94), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n693), .A2(G5), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G171), .B2(new_n693), .ZN(new_n731));
  INV_X1    g306(.A(G1961), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(G29), .A2(G35), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G162), .B2(G29), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G2090), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n735), .B(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT31), .B(G11), .Z(new_n739));
  INV_X1    g314(.A(KEYINPUT30), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n714), .B1(new_n740), .B2(G28), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(KEYINPUT95), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n742), .A2(KEYINPUT95), .B1(new_n740), .B2(G28), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n739), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n628), .B2(new_n714), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n726), .B2(new_n727), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n738), .B(new_n747), .C1(G2084), .C2(new_n715), .ZN(new_n748));
  NOR2_X1   g323(.A1(G164), .A2(new_n714), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G27), .B2(new_n714), .ZN(new_n750));
  INV_X1    g325(.A(G2078), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n689), .A2(G19), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n557), .B2(new_n689), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(G1341), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n714), .A2(G26), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT28), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n701), .A2(G140), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n485), .A2(G128), .ZN(new_n759));
  OR2_X1    g334(.A1(G104), .A2(G2105), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n760), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n757), .B1(new_n763), .B2(new_n714), .ZN(new_n764));
  INV_X1    g339(.A(G2067), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n750), .A2(new_n751), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n752), .A2(new_n755), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n748), .B(new_n768), .C1(G1966), .C2(new_n698), .ZN(new_n769));
  AND4_X1   g344(.A1(new_n696), .A2(new_n729), .A3(new_n733), .A4(new_n769), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n576), .A2(new_n578), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(new_n693), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n693), .B2(G23), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT33), .B(G1976), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n693), .A2(G6), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G305), .B2(G16), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT32), .B(G1981), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT90), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n775), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n689), .A2(G22), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G166), .B2(new_n689), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(G1971), .Z(new_n783));
  NOR2_X1   g358(.A1(new_n777), .A2(new_n779), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n773), .B2(new_n774), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n780), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n786), .A2(KEYINPUT34), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(KEYINPUT34), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n714), .A2(G25), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT84), .Z(new_n790));
  AOI22_X1  g365(.A1(new_n701), .A2(G131), .B1(G119), .B2(new_n485), .ZN(new_n791));
  INV_X1    g366(.A(G95), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(new_n467), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT85), .ZN(new_n794));
  OAI21_X1  g369(.A(G2104), .B1(new_n467), .B2(G107), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT86), .Z(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n790), .B1(new_n798), .B2(G29), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT35), .B(G1991), .Z(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT87), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n799), .B(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n689), .A2(G24), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n591), .B(KEYINPUT89), .Z(new_n804));
  AOI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(new_n689), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(new_n681), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n787), .A2(new_n788), .A3(new_n802), .A4(new_n806), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT91), .B(KEYINPUT36), .Z(new_n808));
  OR2_X1    g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n608), .A2(G16), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G4), .B2(G16), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT92), .B(G1348), .ZN(new_n812));
  OAI22_X1  g387(.A1(new_n728), .A2(KEYINPUT94), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n811), .B2(new_n812), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n807), .A2(new_n808), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n770), .A2(new_n809), .A3(new_n814), .A4(new_n815), .ZN(G150));
  INV_X1    g391(.A(G150), .ZN(G311));
  NAND2_X1  g392(.A1(new_n608), .A2(G559), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT38), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n513), .A2(G55), .ZN(new_n820));
  INV_X1    g395(.A(G93), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(new_n549), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(KEYINPUT99), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT99), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n820), .B(new_n824), .C1(new_n821), .C2(new_n549), .ZN(new_n825));
  NAND2_X1  g400(.A1(G80), .A2(G543), .ZN(new_n826));
  INV_X1    g401(.A(G67), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n603), .B2(new_n827), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n823), .A2(new_n825), .B1(G651), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n557), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n819), .B(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n832), .A2(KEYINPUT39), .ZN(new_n833));
  INV_X1    g408(.A(G860), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(KEYINPUT39), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n829), .A2(new_n834), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT37), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(G145));
  OR2_X1    g414(.A1(G102), .A2(G2105), .ZN(new_n840));
  OAI21_X1  g415(.A(G2105), .B1(KEYINPUT69), .B2(G114), .ZN(new_n841));
  AND2_X1   g416(.A1(KEYINPUT69), .A2(G114), .ZN(new_n842));
  OAI211_X1 g417(.A(G2104), .B(new_n840), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  OAI211_X1 g418(.A(G126), .B(G2105), .C1(new_n474), .C2(new_n475), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(KEYINPUT100), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n843), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n846), .A2(new_n496), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n762), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n707), .B(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n725), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n796), .B(new_n634), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT101), .ZN(new_n855));
  INV_X1    g430(.A(G118), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n854), .A2(new_n855), .B1(new_n856), .B2(G2105), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n855), .B2(new_n854), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n485), .A2(G130), .ZN(new_n859));
  INV_X1    g434(.A(G142), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n858), .B(new_n859), .C1(new_n860), .C2(new_n468), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n853), .B(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n852), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT102), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n852), .A2(new_n862), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(G162), .B(new_n628), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(G160), .ZN(new_n868));
  OR3_X1    g443(.A1(new_n852), .A2(new_n864), .A3(new_n862), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  XOR2_X1   g445(.A(KEYINPUT103), .B(G37), .Z(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n868), .B1(new_n852), .B2(new_n862), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n872), .B1(new_n863), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g451(.A(new_n829), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n611), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n620), .B(new_n831), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n607), .A2(new_n571), .ZN(new_n880));
  NAND4_X1  g455(.A1(G299), .A2(new_n601), .A3(new_n600), .A4(new_n606), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT41), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n607), .A2(new_n886), .A3(new_n571), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n881), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n886), .B1(new_n607), .B2(new_n571), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n885), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT105), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n892), .B(new_n885), .C1(new_n888), .C2(new_n889), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(new_n882), .B2(new_n885), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n880), .A2(KEYINPUT106), .A3(KEYINPUT41), .A4(new_n881), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n891), .A2(new_n893), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n884), .B1(new_n898), .B2(new_n879), .ZN(new_n899));
  XNOR2_X1  g474(.A(G166), .B(G290), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n771), .B(G305), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n900), .B(new_n901), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n902), .B(KEYINPUT42), .Z(new_n903));
  XNOR2_X1  g478(.A(new_n899), .B(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n878), .B1(new_n904), .B2(new_n611), .ZN(G295));
  OAI21_X1  g480(.A(new_n878), .B1(new_n904), .B2(new_n611), .ZN(G331));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n888), .A2(new_n885), .A3(new_n889), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT109), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n910), .B1(new_n539), .B2(new_n540), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n527), .A2(new_n529), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT72), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n913), .A2(KEYINPUT107), .A3(new_n530), .A4(new_n538), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(G301), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(G168), .A2(KEYINPUT107), .A3(G171), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n831), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  INV_X1    g493(.A(new_n831), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI22_X1  g495(.A1(new_n908), .A2(new_n909), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n909), .B1(new_n882), .B2(new_n885), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n880), .A2(KEYINPUT104), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n923), .A2(KEYINPUT41), .A3(new_n881), .A4(new_n887), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n831), .A2(new_n915), .A3(new_n916), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n877), .A2(new_n830), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n829), .A2(new_n557), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n915), .A2(new_n916), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n926), .B1(new_n929), .B2(KEYINPUT108), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n920), .A2(new_n931), .A3(new_n917), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n921), .A2(new_n925), .B1(new_n882), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT110), .B1(new_n934), .B2(new_n902), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n926), .A2(new_n929), .A3(KEYINPUT108), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n918), .A2(new_n919), .A3(new_n931), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n882), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n925), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n920), .A2(new_n917), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(new_n924), .B2(KEYINPUT109), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n938), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n943));
  INV_X1    g518(.A(new_n902), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n935), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n940), .A2(new_n883), .ZN(new_n948));
  INV_X1    g523(.A(new_n933), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n948), .B1(new_n898), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n872), .B1(new_n950), .B2(new_n902), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n946), .A2(new_n947), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(G37), .B1(new_n950), .B2(new_n902), .ZN(new_n953));
  AOI22_X1  g528(.A1(new_n890), .A2(KEYINPUT105), .B1(new_n895), .B2(new_n896), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n933), .B1(new_n954), .B2(new_n893), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n944), .B1(new_n955), .B2(new_n948), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n947), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n907), .B1(new_n952), .B2(new_n957), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n925), .B(new_n940), .C1(KEYINPUT109), .C2(new_n924), .ZN(new_n959));
  AOI211_X1 g534(.A(KEYINPUT110), .B(new_n902), .C1(new_n959), .C2(new_n938), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n943), .B1(new_n942), .B2(new_n944), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n950), .A2(new_n902), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n871), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT43), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G37), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n956), .A2(new_n963), .A3(new_n947), .A4(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n953), .A2(KEYINPUT111), .A3(new_n947), .A4(new_n956), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n965), .A2(new_n969), .A3(KEYINPUT44), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n958), .A2(new_n971), .ZN(G397));
  INV_X1    g547(.A(KEYINPUT123), .ZN(new_n973));
  INV_X1    g548(.A(G1384), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n849), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G40), .ZN(new_n978));
  AOI211_X1 g553(.A(new_n978), .B(new_n470), .C1(new_n472), .C2(new_n480), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n505), .A2(new_n974), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n977), .B(new_n979), .C1(new_n976), .C2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G1966), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n980), .A2(KEYINPUT50), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT50), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n849), .A2(new_n985), .A3(new_n974), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n984), .A2(new_n979), .A3(new_n986), .ZN(new_n987));
  OR2_X1    g562(.A1(new_n987), .A2(G2084), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n983), .A2(new_n988), .A3(G168), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(G8), .ZN(new_n990));
  AND2_X1   g565(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n989), .A2(G8), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G8), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(new_n983), .B2(new_n988), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(G286), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n992), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n771), .A2(G1976), .ZN(new_n1000));
  INV_X1    g575(.A(new_n470), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n471), .A2(KEYINPUT68), .A3(new_n467), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n479), .B1(new_n478), .B2(G2105), .ZN(new_n1003));
  OAI211_X1 g578(.A(G40), .B(new_n1001), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1000), .B(G8), .C1(new_n1004), .C2(new_n975), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT52), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n504), .A2(new_n847), .B1(new_n493), .B2(new_n495), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1384), .B1(new_n1007), .B2(new_n846), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n979), .ZN(new_n1009));
  INV_X1    g584(.A(G1976), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT52), .B1(G288), .B2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1009), .A2(G8), .A3(new_n1011), .A4(new_n1000), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1006), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1981), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n583), .A2(new_n584), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT115), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n583), .A2(new_n584), .A3(new_n1017), .A4(new_n1014), .ZN(new_n1018));
  INV_X1    g593(.A(G86), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n583), .B1(new_n1019), .B2(new_n549), .ZN(new_n1020));
  AOI22_X1  g595(.A1(new_n1016), .A2(new_n1018), .B1(G1981), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT49), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1009), .A2(G8), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1020), .A2(G1981), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT49), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1023), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1013), .B1(new_n1022), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n980), .A2(new_n976), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n849), .A2(KEYINPUT45), .A3(new_n974), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(new_n979), .A3(new_n1031), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT113), .B(G1971), .Z(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G2090), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n984), .A2(new_n979), .A3(new_n986), .A4(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT114), .ZN(new_n1039));
  NOR2_X1   g614(.A1(G166), .A2(new_n996), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n1040), .B(KEYINPUT55), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1035), .A2(new_n1042), .A3(new_n1037), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1039), .A2(new_n1041), .A3(G8), .A4(new_n1043), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1029), .A2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(KEYINPUT117), .B(new_n979), .C1(new_n1008), .C2(new_n985), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n985), .B1(new_n849), .B2(new_n974), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1047), .B1(new_n1048), .B2(new_n1004), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n505), .A2(new_n985), .A3(new_n974), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1046), .A2(new_n1049), .A3(new_n1036), .A4(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n996), .B1(new_n1051), .B2(new_n1035), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1052), .A2(new_n1041), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1032), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n751), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1055), .A2(new_n1056), .B1(new_n732), .B2(new_n987), .ZN(new_n1057));
  OR3_X1    g632(.A1(new_n981), .A2(new_n1056), .A3(G2078), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  XOR2_X1   g634(.A(G171), .B(KEYINPUT54), .Z(new_n1060));
  NOR3_X1   g635(.A1(new_n1056), .A2(new_n978), .A3(G2078), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1001), .B(new_n1061), .C1(new_n467), .C2(new_n471), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(new_n975), .B2(new_n976), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1060), .B1(new_n1031), .B2(new_n1063), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1059), .A2(new_n1060), .B1(new_n1064), .B2(new_n1057), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n999), .A2(new_n1045), .A3(new_n1053), .A4(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT56), .B(G2072), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1054), .A2(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n571), .B(KEYINPUT57), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1046), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1072));
  INV_X1    g647(.A(G1956), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1072), .A2(KEYINPUT119), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT119), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1071), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1054), .A2(new_n1067), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1078), .B1(new_n1081), .B2(new_n1074), .ZN(new_n1082));
  OAI211_X1 g657(.A(KEYINPUT61), .B(new_n1077), .C1(new_n1082), .C2(new_n1069), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n975), .A2(new_n1004), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1085), .B(G1341), .ZN(new_n1086));
  OAI22_X1  g661(.A1(new_n1032), .A2(G1996), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n557), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(new_n1089), .A3(KEYINPUT59), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(KEYINPUT59), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1087), .A2(new_n557), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G1348), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n987), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1084), .A2(new_n765), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1095), .A2(new_n607), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n607), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT60), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT60), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n608), .A2(new_n1100), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1093), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1068), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1069), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1081), .A2(new_n1074), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1103), .A2(new_n1104), .B1(new_n1105), .B2(new_n1071), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1083), .B(new_n1102), .C1(new_n1106), .C2(KEYINPUT61), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1082), .A2(new_n1069), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1077), .B1(new_n1108), .B2(new_n1098), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1066), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT118), .B(KEYINPUT63), .Z(new_n1111));
  OAI211_X1 g686(.A(new_n1029), .B(new_n1044), .C1(new_n1041), .C2(new_n1052), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n997), .A2(G168), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1039), .A2(G8), .A3(new_n1043), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1041), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n997), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1045), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1114), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n771), .A2(new_n1010), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1121), .B1(new_n1028), .B2(new_n1022), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1024), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT116), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT116), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1084), .A2(new_n996), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1021), .B2(KEYINPUT49), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1125), .B(new_n1024), .C1(new_n1129), .C2(new_n1121), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1124), .A2(new_n1130), .A3(new_n1127), .ZN(new_n1131));
  OR3_X1    g706(.A1(new_n1044), .A2(new_n1129), .A3(new_n1013), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1120), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n973), .B1(new_n1110), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1133), .B1(new_n1114), .B2(new_n1119), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1070), .B1(new_n1081), .B2(new_n1074), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1098), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1093), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1138), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1142), .B1(new_n1144), .B2(new_n1139), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1143), .B1(new_n1108), .B2(new_n1138), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1141), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1137), .B(KEYINPUT123), .C1(new_n1147), .C2(new_n1066), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n999), .A2(KEYINPUT62), .ZN(new_n1149));
  AOI21_X1  g724(.A(G301), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1045), .A2(new_n1150), .A3(new_n1053), .ZN(new_n1151));
  OR3_X1    g726(.A1(new_n1149), .A2(new_n1151), .A3(KEYINPUT124), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n999), .A2(KEYINPUT62), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT124), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1136), .A2(new_n1148), .A3(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n977), .A2(new_n1004), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n796), .B(new_n800), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(G1996), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT112), .ZN(new_n1163));
  INV_X1    g738(.A(new_n725), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n762), .B(new_n765), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1166), .B1(G1996), .B2(new_n1164), .ZN(new_n1167));
  OAI22_X1  g742(.A1(new_n1163), .A2(new_n1164), .B1(new_n1158), .B2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n591), .B(new_n681), .ZN(new_n1169));
  AOI211_X1 g744(.A(new_n1160), .B(new_n1168), .C1(new_n1157), .C2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1156), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n797), .A2(new_n800), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n762), .A2(G2067), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1158), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(KEYINPUT125), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1177), .A2(KEYINPUT126), .A3(new_n1178), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1157), .B1(new_n1166), .B2(new_n1164), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n1163), .A2(KEYINPUT46), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1163), .A2(KEYINPUT46), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  OR2_X1    g761(.A1(new_n1186), .A2(KEYINPUT47), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(KEYINPUT47), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1168), .A2(new_n1160), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1157), .A2(new_n681), .A3(new_n591), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(KEYINPUT48), .ZN(new_n1191));
  AOI22_X1  g766(.A1(new_n1187), .A2(new_n1188), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1181), .A2(new_n1182), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1171), .A2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g769(.A1(new_n952), .A2(new_n957), .ZN(new_n1196));
  NOR2_X1   g770(.A1(new_n461), .A2(G227), .ZN(new_n1197));
  NAND4_X1  g771(.A1(new_n687), .A2(new_n654), .A3(new_n875), .A4(new_n1197), .ZN(new_n1198));
  NOR2_X1   g772(.A1(new_n1196), .A2(new_n1198), .ZN(G308));
  AND3_X1   g773(.A1(new_n687), .A2(new_n654), .A3(new_n1197), .ZN(new_n1200));
  OAI211_X1 g774(.A(new_n1200), .B(new_n875), .C1(new_n957), .C2(new_n952), .ZN(G225));
endmodule


