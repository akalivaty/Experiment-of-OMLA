//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1273,
    new_n1274, new_n1275, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342;
  NOR2_X1   g0000(.A1(G50), .A2(G58), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  INV_X1    g0009(.A(KEYINPUT65), .ZN(new_n210));
  OR2_X1    g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G50), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n217), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  INV_X1    g0025(.A(G68), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n219), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n211), .A2(new_n225), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(new_n210), .B2(new_n209), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G226), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G68), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT67), .ZN(new_n250));
  XOR2_X1   g0050(.A(G50), .B(G58), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n248), .B(new_n252), .ZN(G351));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n230), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n219), .A2(KEYINPUT8), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT8), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G58), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n231), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n260), .A2(new_n262), .B1(G150), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n231), .B1(new_n201), .B2(new_n226), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n256), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n231), .A2(G1), .ZN(new_n268));
  OAI21_X1  g0068(.A(KEYINPUT70), .B1(new_n268), .B2(new_n213), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G13), .A3(G20), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(G20), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT70), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(new_n273), .A3(G50), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n269), .A2(new_n256), .A3(new_n271), .A4(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n271), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n213), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(KEYINPUT71), .B1(new_n267), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT8), .B(G58), .ZN(new_n280));
  INV_X1    g0080(.A(G150), .ZN(new_n281));
  INV_X1    g0081(.A(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n231), .A2(new_n282), .ZN(new_n283));
  OAI22_X1  g0083(.A1(new_n280), .A2(new_n261), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n255), .B1(new_n284), .B2(new_n265), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT71), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n285), .A2(new_n286), .A3(new_n277), .A4(new_n275), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n279), .A2(KEYINPUT9), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT72), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n279), .A2(KEYINPUT72), .A3(new_n287), .A4(KEYINPUT9), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(KEYINPUT9), .B1(new_n279), .B2(new_n287), .ZN(new_n293));
  INV_X1    g0093(.A(G41), .ZN(new_n294));
  INV_X1    g0094(.A(G45), .ZN(new_n295));
  AOI21_X1  g0095(.A(G1), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G41), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n297), .A2(G1), .A3(G13), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n296), .A2(new_n298), .A3(G274), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n270), .B1(G41), .B2(G45), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(G226), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT3), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n282), .ZN(new_n304));
  NAND2_X1  g0104(.A1(KEYINPUT3), .A2(G33), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AND2_X1   g0106(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n307));
  NOR2_X1   g0107(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n306), .A2(new_n309), .A3(G222), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n306), .A2(G223), .A3(G1698), .ZN(new_n311));
  AND2_X1   g0111(.A1(KEYINPUT3), .A2(G33), .ZN(new_n312));
  NOR2_X1   g0112(.A1(KEYINPUT3), .A2(G33), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G77), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n310), .A2(new_n311), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n302), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G190), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n293), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(G200), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n292), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT10), .ZN(new_n325));
  INV_X1    g0125(.A(G200), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT73), .B1(new_n318), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT10), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT73), .ZN(new_n329));
  INV_X1    g0129(.A(G1698), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n304), .B2(new_n305), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n331), .A2(G223), .B1(new_n314), .B2(G77), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n298), .B1(new_n332), .B2(new_n310), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n329), .B(G200), .C1(new_n333), .C2(new_n302), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n327), .A2(new_n328), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AND4_X1   g0136(.A1(KEYINPUT74), .A2(new_n292), .A3(new_n322), .A4(new_n336), .ZN(new_n337));
  NOR3_X1   g0137(.A1(new_n335), .A2(new_n293), .A3(new_n321), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT74), .B1(new_n338), .B2(new_n292), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n325), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NOR3_X1   g0141(.A1(new_n307), .A2(new_n308), .A3(new_n214), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n220), .A2(new_n330), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n306), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G33), .A2(G97), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT75), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n298), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n317), .A2(new_n296), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G238), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n299), .ZN(new_n351));
  OAI21_X1  g0151(.A(KEYINPUT13), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT69), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n330), .ZN(new_n354));
  NAND2_X1  g0154(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(G226), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n343), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n314), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n317), .B1(new_n358), .B2(new_n346), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n298), .A2(G274), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n349), .A2(G238), .B1(new_n360), .B2(new_n296), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT13), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n359), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n352), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G190), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n352), .A2(KEYINPUT76), .A3(new_n363), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT76), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n359), .A2(new_n361), .A3(new_n367), .A4(new_n362), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n366), .A2(G200), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n276), .A2(new_n226), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n370), .B(KEYINPUT12), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n263), .A2(G50), .B1(G20), .B2(new_n226), .ZN(new_n372));
  INV_X1    g0172(.A(G77), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n372), .B1(new_n373), .B2(new_n261), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n374), .A2(KEYINPUT11), .A3(new_n255), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n276), .A2(new_n255), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n376), .A2(G68), .A3(new_n272), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n371), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT11), .B1(new_n374), .B2(new_n255), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n365), .A2(new_n369), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n366), .A2(G169), .A3(new_n368), .ZN(new_n383));
  NAND2_X1  g0183(.A1(KEYINPUT77), .A2(KEYINPUT14), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n384), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n366), .A2(new_n368), .A3(G169), .A4(new_n386), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n385), .A2(new_n387), .B1(G179), .B2(new_n364), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n382), .B1(new_n388), .B2(new_n381), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT16), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G58), .A2(G68), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n231), .B1(new_n227), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n263), .A2(G159), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT78), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n391), .ZN(new_n396));
  NOR2_X1   g0196(.A1(G58), .A2(G68), .ZN(new_n397));
  OAI21_X1  g0197(.A(G20), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT78), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(new_n399), .A3(new_n393), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT7), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n306), .B2(G20), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n314), .A2(KEYINPUT7), .A3(new_n231), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n226), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n390), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT7), .B1(new_n314), .B2(new_n231), .ZN(new_n407));
  NOR4_X1   g0207(.A1(new_n312), .A2(new_n313), .A3(new_n402), .A4(G20), .ZN(new_n408));
  OAI21_X1  g0208(.A(G68), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n409), .A2(KEYINPUT16), .A3(new_n400), .A4(new_n395), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n406), .A2(new_n255), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n376), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n260), .A2(new_n272), .ZN(new_n413));
  OAI22_X1  g0213(.A1(new_n412), .A2(new_n413), .B1(new_n271), .B2(new_n260), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT18), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n298), .A2(G232), .A3(new_n300), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n299), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g0219(.A(G226), .B(G1698), .C1(new_n312), .C2(new_n313), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G87), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n354), .B(new_n355), .C1(new_n312), .C2(new_n313), .ZN(new_n422));
  INV_X1    g0222(.A(G223), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n420), .B(new_n421), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n419), .B1(new_n424), .B2(new_n317), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(G169), .ZN(new_n426));
  AOI211_X1 g0226(.A(G179), .B(new_n419), .C1(new_n424), .C2(new_n317), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n416), .A2(new_n417), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n417), .B1(new_n416), .B2(new_n428), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  XOR2_X1   g0231(.A(KEYINPUT80), .B(KEYINPUT17), .Z(new_n432));
  NAND2_X1  g0232(.A1(new_n424), .A2(new_n317), .ZN(new_n433));
  INV_X1    g0233(.A(new_n419), .ZN(new_n434));
  AND4_X1   g0234(.A1(KEYINPUT79), .A2(new_n433), .A3(new_n320), .A4(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n425), .A2(new_n320), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT79), .B1(new_n425), .B2(G200), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n432), .B1(new_n438), .B2(new_n416), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(new_n436), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n425), .A2(KEYINPUT79), .A3(new_n320), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n409), .A2(new_n400), .A3(new_n395), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n256), .B1(new_n443), .B2(new_n390), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n414), .B1(new_n444), .B2(new_n410), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT80), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT17), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n442), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n439), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n431), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n349), .A2(G244), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n299), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n331), .A2(G238), .ZN(new_n453));
  INV_X1    g0253(.A(G107), .ZN(new_n454));
  OAI221_X1 g0254(.A(new_n453), .B1(new_n454), .B2(new_n306), .C1(new_n220), .C2(new_n422), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n452), .B1(new_n455), .B2(new_n317), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n260), .A2(new_n263), .B1(G20), .B2(G77), .ZN(new_n457));
  XNOR2_X1  g0257(.A(KEYINPUT15), .B(G87), .ZN(new_n458));
  OR2_X1    g0258(.A1(new_n458), .A2(new_n261), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n256), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n376), .A2(G77), .A3(new_n272), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(G77), .B2(new_n271), .ZN(new_n462));
  OAI22_X1  g0262(.A1(new_n456), .A2(G169), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G179), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n456), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n456), .A2(G190), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n462), .A2(new_n460), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n468), .B(new_n469), .C1(new_n326), .C2(new_n456), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n319), .A2(G179), .ZN(new_n471));
  OAI22_X1  g0271(.A1(new_n318), .A2(G169), .B1(new_n267), .B2(new_n278), .ZN(new_n472));
  OR2_X1    g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n467), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  NOR4_X1   g0274(.A1(new_n341), .A2(new_n389), .A3(new_n450), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n270), .A2(G33), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n376), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT25), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(new_n271), .B2(G107), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n271), .A2(new_n478), .A3(G107), .ZN(new_n481));
  OAI22_X1  g0281(.A1(new_n477), .A2(new_n454), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n231), .B(G87), .C1(new_n312), .C2(new_n313), .ZN(new_n483));
  AND2_X1   g0283(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n484));
  NOR2_X1   g0284(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n306), .A2(new_n231), .A3(G87), .A4(new_n484), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT86), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n489), .B(KEYINPUT23), .C1(new_n231), .C2(G107), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n231), .A2(G33), .A3(G116), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT23), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(new_n454), .A3(G20), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n490), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT23), .B1(new_n231), .B2(G107), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT86), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n487), .A2(new_n488), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT87), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT24), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n500), .A2(new_n255), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n497), .A2(new_n498), .ZN(new_n502));
  AND4_X1   g0302(.A1(new_n496), .A2(new_n490), .A3(new_n491), .A4(new_n493), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n503), .A2(KEYINPUT87), .A3(new_n488), .A4(new_n487), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n504), .A3(KEYINPUT24), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n482), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g0306(.A(KEYINPUT5), .B(G41), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n295), .A2(G1), .ZN(new_n508));
  INV_X1    g0308(.A(new_n230), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n297), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G264), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n507), .A2(new_n298), .A3(G274), .A4(new_n508), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g0315(.A(G257), .B(G1698), .C1(new_n312), .C2(new_n313), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G33), .A2(G294), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n516), .B(new_n517), .C1(new_n422), .C2(new_n216), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT88), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n306), .A2(new_n309), .A3(G250), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n521), .A2(KEYINPUT88), .A3(new_n516), .A4(new_n517), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n298), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n515), .B1(new_n523), .B2(KEYINPUT89), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT89), .ZN(new_n525));
  AOI211_X1 g0325(.A(new_n525), .B(new_n298), .C1(new_n520), .C2(new_n522), .ZN(new_n526));
  OAI21_X1  g0326(.A(G169), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n523), .A2(new_n512), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n528), .A2(G179), .A3(new_n513), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n506), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n482), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n502), .A2(new_n504), .A3(KEYINPUT24), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n500), .A2(new_n255), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n520), .A2(new_n522), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n317), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n525), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n523), .A2(KEYINPUT89), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n537), .A2(new_n320), .A3(new_n538), .A4(new_n515), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n536), .A2(new_n513), .A3(new_n511), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n326), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n534), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n530), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT81), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n544), .A2(KEYINPUT4), .ZN(new_n545));
  INV_X1    g0345(.A(G244), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n422), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G283), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n331), .B2(G250), .ZN(new_n550));
  INV_X1    g0350(.A(new_n545), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n306), .A2(new_n309), .A3(new_n551), .A4(G244), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n547), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT82), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT82), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n547), .A2(new_n550), .A3(new_n552), .A4(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n317), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n514), .B1(G257), .B2(new_n510), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n464), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT6), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n560), .A2(new_n221), .A3(G107), .ZN(new_n561));
  XNOR2_X1  g0361(.A(G97), .B(G107), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n561), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  OAI22_X1  g0363(.A1(new_n563), .A2(new_n231), .B1(new_n373), .B2(new_n283), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n454), .B1(new_n403), .B2(new_n404), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n255), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n276), .A2(new_n221), .ZN(new_n567));
  INV_X1    g0367(.A(new_n477), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G97), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n558), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n298), .B1(new_n553), .B2(KEYINPUT82), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n571), .B1(new_n572), .B2(new_n556), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n559), .B(new_n570), .C1(G169), .C2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n557), .A2(G190), .A3(new_n558), .ZN(new_n575));
  INV_X1    g0375(.A(new_n570), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n575), .B(new_n576), .C1(new_n326), .C2(new_n573), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(G264), .B(G1698), .C1(new_n312), .C2(new_n313), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n304), .A2(G303), .A3(new_n305), .ZN(new_n580));
  OAI21_X1  g0380(.A(G257), .B1(new_n312), .B2(new_n313), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n354), .A2(new_n355), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n317), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n270), .A2(G45), .ZN(new_n585));
  NOR2_X1   g0385(.A1(KEYINPUT5), .A2(G41), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(KEYINPUT5), .A2(G41), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n585), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n510), .A2(G270), .B1(new_n360), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(G116), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n276), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n256), .A2(G116), .A3(new_n271), .A4(new_n476), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n254), .A2(new_n230), .B1(G20), .B2(new_n592), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n548), .B(new_n231), .C1(G33), .C2(new_n221), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n595), .A2(KEYINPUT20), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT20), .B1(new_n595), .B2(new_n596), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n593), .B(new_n594), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n591), .A2(KEYINPUT21), .A3(G169), .A4(new_n599), .ZN(new_n600));
  AND2_X1   g0400(.A1(KEYINPUT5), .A2(G41), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n508), .B1(new_n601), .B2(new_n586), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(G270), .A3(new_n298), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n513), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n317), .B2(new_n583), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(G179), .A3(new_n599), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n600), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(G169), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n584), .B2(new_n590), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT21), .B1(new_n609), .B2(new_n599), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NOR3_X1   g0411(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n345), .A2(KEYINPUT75), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n345), .A2(KEYINPUT75), .ZN(new_n614));
  OAI21_X1  g0414(.A(KEYINPUT19), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n612), .B1(new_n615), .B2(new_n231), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT19), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n261), .B2(new_n221), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT83), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n306), .A2(new_n231), .A3(G68), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT83), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n621), .B(new_n617), .C1(new_n261), .C2(new_n221), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n619), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n255), .B1(new_n616), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n458), .A2(new_n276), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n477), .A2(new_n458), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n508), .A2(new_n216), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n298), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n298), .A2(G274), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n629), .B1(new_n630), .B2(new_n585), .ZN(new_n631));
  OAI211_X1 g0431(.A(G244), .B(G1698), .C1(new_n312), .C2(new_n313), .ZN(new_n632));
  NAND2_X1  g0432(.A1(G33), .A2(G116), .ZN(new_n633));
  INV_X1    g0433(.A(G238), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n632), .B(new_n633), .C1(new_n422), .C2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n631), .B1(new_n317), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n464), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n627), .B(new_n637), .C1(G169), .C2(new_n636), .ZN(new_n638));
  AOI21_X1  g0438(.A(G20), .B1(new_n304), .B2(new_n305), .ZN(new_n639));
  AOI22_X1  g0439(.A1(G68), .A2(new_n639), .B1(new_n618), .B2(KEYINPUT83), .ZN(new_n640));
  AOI21_X1  g0440(.A(G20), .B1(new_n346), .B2(KEYINPUT19), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n640), .B(new_n622), .C1(new_n641), .C2(new_n612), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n642), .A2(new_n255), .B1(new_n276), .B2(new_n458), .ZN(new_n643));
  INV_X1    g0443(.A(new_n631), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n635), .A2(new_n317), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(G200), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n644), .A2(new_n645), .A3(G190), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n568), .A2(G87), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n643), .A2(new_n647), .A3(new_n648), .A4(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT84), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n326), .B1(new_n584), .B2(new_n590), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n651), .B1(new_n652), .B2(new_n599), .ZN(new_n653));
  INV_X1    g0453(.A(new_n599), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n654), .B(KEYINPUT84), .C1(new_n605), .C2(new_n326), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n605), .A2(G190), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n653), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n611), .A2(new_n638), .A3(new_n650), .A4(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n578), .A2(new_n658), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n475), .A2(new_n543), .A3(new_n659), .ZN(G372));
  INV_X1    g0460(.A(new_n611), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n530), .A2(new_n661), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n635), .A2(KEYINPUT90), .A3(new_n317), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT90), .B1(new_n635), .B2(new_n317), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n644), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n608), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT91), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n627), .A2(new_n637), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT91), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n665), .A2(new_n670), .A3(new_n608), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n667), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n648), .A2(new_n624), .A3(new_n625), .A4(new_n649), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(G200), .B2(new_n665), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NOR4_X1   g0476(.A1(new_n662), .A2(new_n676), .A3(new_n578), .A4(new_n542), .ZN(new_n677));
  INV_X1    g0477(.A(new_n574), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT26), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n678), .A2(new_n679), .A3(new_n672), .A4(new_n675), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n638), .A2(new_n650), .ZN(new_n681));
  OAI21_X1  g0481(.A(KEYINPUT26), .B1(new_n574), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n680), .A2(new_n672), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n475), .B1(new_n677), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n473), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT92), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n340), .A2(new_n686), .ZN(new_n687));
  OAI211_X1 g0487(.A(KEYINPUT92), .B(new_n325), .C1(new_n337), .C2(new_n339), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n388), .A2(new_n381), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n382), .A2(new_n466), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n449), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n431), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n685), .B1(new_n689), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n684), .A2(new_n694), .ZN(G369));
  NAND3_X1  g0495(.A1(new_n270), .A2(new_n231), .A3(G13), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G213), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G343), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n534), .A2(new_n701), .ZN(new_n702));
  AOI22_X1  g0502(.A1(new_n543), .A2(new_n702), .B1(new_n530), .B2(new_n701), .ZN(new_n703));
  INV_X1    g0503(.A(new_n701), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n654), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n661), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n611), .A2(new_n657), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n706), .B1(new_n707), .B2(new_n705), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n703), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n611), .A2(new_n701), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n713), .A2(new_n530), .A3(new_n542), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n530), .B2(new_n704), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n711), .A2(new_n715), .ZN(G399));
  INV_X1    g0516(.A(new_n207), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(G41), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n612), .A2(new_n592), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(G1), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n228), .B2(new_n719), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT28), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT94), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n680), .A2(new_n672), .A3(new_n682), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n578), .A2(new_n542), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n527), .A2(new_n529), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n611), .B1(new_n727), .B2(new_n506), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n668), .B1(KEYINPUT91), .B2(new_n666), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n674), .B1(new_n729), .B2(new_n671), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n726), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n701), .B1(new_n725), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n724), .B1(new_n732), .B2(KEYINPUT29), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n704), .B1(new_n677), .B2(new_n683), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT29), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(KEYINPUT94), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n679), .B1(new_n730), .B2(new_n678), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n638), .A2(new_n650), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n570), .B1(new_n573), .B2(G169), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n738), .A2(new_n740), .A3(new_n679), .A4(new_n559), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n672), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n737), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n701), .B1(new_n743), .B2(new_n731), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(KEYINPUT29), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n733), .A2(new_n736), .A3(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n659), .A2(new_n543), .A3(new_n704), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT30), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n584), .A2(new_n590), .A3(G179), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n536), .A2(new_n511), .A3(new_n749), .A4(new_n636), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n557), .A2(new_n558), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n748), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n646), .A2(new_n591), .A3(new_n464), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n573), .A2(new_n753), .A3(KEYINPUT30), .A4(new_n528), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n665), .A2(KEYINPUT93), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT93), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n756), .B(new_n644), .C1(new_n663), .C2(new_n664), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n755), .A2(new_n751), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n540), .A2(new_n464), .A3(new_n591), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n752), .B(new_n754), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(new_n701), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT31), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n760), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n747), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n765), .A2(G330), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n746), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n723), .B1(new_n769), .B2(G1), .ZN(G364));
  XNOR2_X1  g0570(.A(new_n709), .B(KEYINPUT95), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n231), .A2(G13), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT96), .Z(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G45), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G1), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n718), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n772), .B(new_n778), .C1(G330), .C2(new_n708), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n207), .A2(G355), .A3(new_n306), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(G116), .B2(new_n207), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n252), .A2(G45), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n306), .B(new_n717), .C1(new_n295), .C2(new_n229), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G13), .A2(G33), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n230), .B1(G20), .B2(new_n608), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n777), .B1(new_n784), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n231), .A2(G190), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n464), .A2(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G311), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G179), .A2(G200), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n231), .B1(new_n796), .B2(G190), .ZN(new_n797));
  INV_X1    g0597(.A(G294), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n794), .A2(new_n795), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n320), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n799), .B1(G326), .B2(new_n801), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT100), .Z(new_n803));
  XNOR2_X1  g0603(.A(KEYINPUT33), .B(G317), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n804), .A2(KEYINPUT101), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n800), .A2(G190), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(KEYINPUT101), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n231), .A2(new_n320), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n793), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n792), .A2(new_n796), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G322), .A2(new_n811), .B1(new_n813), .B2(G329), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n326), .A2(G179), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n792), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n306), .B1(new_n817), .B2(G283), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n809), .A2(new_n815), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n820), .A2(KEYINPUT98), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(KEYINPUT98), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n819), .B1(G303), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n803), .A2(new_n808), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n797), .A2(new_n221), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n806), .B2(G68), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT99), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n817), .A2(G107), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n830), .B(new_n306), .C1(new_n373), .C2(new_n794), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n810), .B(KEYINPUT97), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n831), .B1(G58), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(G159), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n812), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT32), .ZN(new_n836));
  INV_X1    g0636(.A(new_n801), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n835), .A2(new_n836), .B1(new_n213), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(new_n836), .B2(new_n835), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n824), .A2(G87), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n829), .A2(new_n833), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n826), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n791), .B1(new_n788), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n787), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n708), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n779), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(G396));
  NAND2_X1  g0647(.A1(new_n466), .A2(new_n704), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n470), .B1(new_n469), .B2(new_n704), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n849), .B1(new_n467), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n734), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n704), .B(new_n851), .C1(new_n677), .C2(new_n683), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n855), .A2(new_n767), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT103), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n777), .B1(new_n855), .B2(new_n767), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n788), .A2(new_n785), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n778), .B1(new_n373), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n788), .ZN(new_n862));
  AOI22_X1  g0662(.A1(G294), .A2(new_n811), .B1(new_n817), .B2(G87), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n863), .B1(new_n795), .B2(new_n812), .C1(new_n823), .C2(new_n454), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n314), .B1(new_n794), .B2(new_n592), .ZN(new_n865));
  INV_X1    g0665(.A(new_n806), .ZN(new_n866));
  INV_X1    g0666(.A(G283), .ZN(new_n867));
  INV_X1    g0667(.A(G303), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n866), .A2(new_n867), .B1(new_n837), .B2(new_n868), .ZN(new_n869));
  NOR4_X1   g0669(.A1(new_n864), .A2(new_n827), .A3(new_n865), .A4(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n794), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n871), .A2(G159), .B1(G137), .B2(new_n801), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n281), .B2(new_n866), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(G143), .B2(new_n832), .ZN(new_n874));
  XOR2_X1   g0674(.A(new_n874), .B(KEYINPUT34), .Z(new_n875));
  OAI21_X1  g0675(.A(new_n306), .B1(new_n816), .B2(new_n226), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(G132), .B2(new_n813), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n877), .B1(new_n219), .B2(new_n797), .C1(new_n213), .C2(new_n823), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n878), .B(KEYINPUT102), .Z(new_n879));
  AOI21_X1  g0679(.A(new_n870), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  OAI221_X1 g0680(.A(new_n861), .B1(new_n862), .B2(new_n880), .C1(new_n851), .C2(new_n786), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n859), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(G384));
  INV_X1    g0683(.A(new_n563), .ZN(new_n884));
  OR2_X1    g0684(.A1(new_n884), .A2(KEYINPUT35), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(KEYINPUT35), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n885), .A2(G116), .A3(new_n232), .A4(new_n886), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT36), .Z(new_n888));
  NAND3_X1  g0688(.A1(new_n229), .A2(G77), .A3(new_n391), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n213), .A2(G68), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n270), .B(G13), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT40), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n445), .A2(new_n699), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n450), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n442), .A2(new_n445), .ZN(new_n896));
  INV_X1    g0696(.A(new_n699), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n416), .B1(new_n428), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n896), .A2(new_n898), .A3(KEYINPUT37), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT37), .B1(new_n896), .B2(new_n898), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n895), .A2(KEYINPUT38), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT106), .ZN(new_n904));
  INV_X1    g0704(.A(new_n894), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n431), .B2(new_n449), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n896), .A2(new_n898), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT37), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n899), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT106), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT38), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n904), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n908), .B1(new_n898), .B2(KEYINPUT105), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(new_n907), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n895), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT38), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n893), .B1(new_n914), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n765), .A2(new_n851), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n385), .A2(new_n387), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n364), .A2(G179), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(new_n923), .A3(new_n382), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT104), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n380), .A2(new_n701), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n382), .B(new_n926), .C1(new_n388), .C2(new_n381), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n925), .B1(new_n924), .B2(new_n927), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n921), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n918), .B1(new_n906), .B2(new_n910), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n903), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n924), .A2(new_n927), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT104), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(new_n929), .A3(new_n928), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n935), .A2(new_n938), .A3(new_n765), .A4(new_n851), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n920), .A2(new_n933), .B1(new_n893), .B2(new_n939), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n475), .A2(new_n765), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n942), .A2(G330), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n903), .A2(new_n934), .A3(KEYINPUT39), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n690), .A2(new_n704), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n904), .A2(new_n913), .B1(new_n918), .B2(new_n917), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n945), .B(new_n947), .C1(new_n948), .C2(KEYINPUT39), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n431), .A2(new_n897), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n932), .B1(new_n854), .B2(new_n848), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n950), .B1(new_n951), .B2(new_n935), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n733), .A2(new_n736), .A3(new_n475), .A4(new_n745), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n694), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n953), .B(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n944), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n270), .B2(new_n774), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n944), .A2(new_n956), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n892), .B1(new_n958), .B2(new_n959), .ZN(G367));
  INV_X1    g0760(.A(KEYINPUT42), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n574), .A2(new_n704), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT109), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n574), .B(new_n577), .C1(new_n576), .C2(new_n704), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n543), .A2(new_n712), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n961), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n964), .A2(new_n965), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(KEYINPUT42), .A3(new_n714), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n704), .B1(new_n643), .B2(new_n649), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT107), .Z(new_n973));
  OR2_X1    g0773(.A1(new_n973), .A2(new_n672), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n730), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT108), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n976), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n530), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(new_n964), .B2(new_n965), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n704), .B1(new_n983), .B2(new_n678), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n971), .A2(new_n981), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(KEYINPUT110), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT110), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n971), .A2(new_n987), .A3(new_n981), .A4(new_n984), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n980), .B2(new_n976), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n971), .B2(new_n984), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n989), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT111), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n711), .A2(new_n966), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n989), .A2(KEYINPUT111), .A3(new_n993), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(KEYINPUT111), .B1(new_n989), .B2(new_n993), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n995), .B(new_n992), .C1(new_n986), .C2(new_n988), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n1000), .A2(new_n1001), .B1(new_n711), .B2(new_n966), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n776), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT45), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n967), .B1(new_n982), .B2(new_n701), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1004), .B1(new_n966), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n715), .A2(new_n969), .A3(KEYINPUT45), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n966), .A2(KEYINPUT44), .A3(new_n1005), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT44), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n715), .B2(new_n969), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  AND3_X1   g0812(.A1(new_n1008), .A2(new_n711), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n711), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n714), .B1(new_n703), .B2(new_n713), .ZN(new_n1016));
  MUX2_X1   g0816(.A(new_n771), .B(new_n709), .S(new_n1016), .Z(new_n1017));
  AOI21_X1  g0817(.A(new_n768), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n718), .B(KEYINPUT41), .Z(new_n1019));
  OAI21_X1  g0819(.A(new_n1003), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n999), .A2(new_n1002), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n789), .B1(new_n207), .B2(new_n458), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n717), .A2(new_n306), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1022), .B1(new_n1023), .B2(new_n243), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n824), .A2(G58), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n306), .B1(new_n810), .B2(new_n281), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n797), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1026), .B1(G68), .B2(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n806), .A2(G159), .B1(new_n801), .B2(G143), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n213), .A2(new_n794), .B1(new_n816), .B2(new_n373), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G137), .B2(new_n813), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1025), .A2(new_n1028), .A3(new_n1029), .A4(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n823), .A2(new_n592), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT46), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n866), .A2(new_n798), .B1(new_n837), .B2(new_n795), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(G107), .B2(new_n1027), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n832), .A2(G303), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n306), .B1(new_n813), .B2(G317), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n816), .A2(new_n221), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G283), .B2(new_n871), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .A4(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1032), .B1(new_n1034), .B2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT47), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n778), .B(new_n1024), .C1(new_n1043), .C2(new_n788), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n976), .B2(new_n844), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1021), .A2(new_n1045), .ZN(G387));
  NAND2_X1  g0846(.A1(new_n703), .A2(new_n787), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n240), .A2(G45), .A3(new_n314), .ZN(new_n1048));
  OAI21_X1  g0848(.A(KEYINPUT50), .B1(new_n280), .B2(G50), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1049), .B(new_n295), .C1(new_n226), .C2(new_n373), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n280), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n314), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n720), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n717), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n789), .B1(new_n207), .B2(new_n454), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n777), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n797), .A2(new_n458), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G50), .B2(new_n811), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT112), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n834), .A2(new_n837), .B1(new_n866), .B2(new_n280), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n794), .A2(new_n226), .B1(new_n812), .B2(new_n281), .ZN(new_n1061));
  NOR4_X1   g0861(.A1(new_n1060), .A2(new_n1061), .A3(new_n314), .A4(new_n1039), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1059), .B(new_n1062), .C1(new_n373), .C2(new_n823), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n823), .A2(new_n798), .B1(new_n867), .B2(new_n797), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n871), .A2(G303), .B1(G311), .B2(new_n806), .ZN(new_n1065));
  INV_X1    g0865(.A(G322), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1065), .B1(new_n1066), .B2(new_n837), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(G317), .B2(new_n832), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1064), .B1(new_n1068), .B2(KEYINPUT48), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT113), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(KEYINPUT48), .B2(new_n1068), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT49), .Z(new_n1072));
  AOI21_X1  g0872(.A(new_n306), .B1(new_n813), .B2(G326), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n592), .B2(new_n816), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1063), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1056), .B1(new_n1075), .B2(new_n788), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1047), .A2(new_n1076), .B1(new_n1017), .B2(new_n776), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n769), .A2(new_n1017), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n718), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n769), .A2(new_n1017), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1077), .B1(new_n1079), .B2(new_n1080), .ZN(G393));
  OAI22_X1  g0881(.A1(new_n823), .A2(new_n867), .B1(new_n1066), .B2(new_n812), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1082), .A2(KEYINPUT115), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(KEYINPUT115), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1083), .A2(new_n314), .A3(new_n830), .A4(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT116), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n811), .A2(G311), .B1(G317), .B2(new_n801), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G294), .A2(new_n871), .B1(new_n1027), .B2(G116), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n868), .B2(new_n866), .ZN(new_n1093));
  NOR4_X1   g0893(.A1(new_n1086), .A2(new_n1090), .A3(new_n1091), .A4(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n794), .A2(new_n280), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n306), .B1(new_n816), .B2(new_n215), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(G143), .C2(new_n813), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1027), .A2(G77), .B1(G50), .B2(new_n806), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1097), .B(new_n1098), .C1(new_n226), .C2(new_n823), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n811), .A2(G159), .B1(G150), .B2(new_n801), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT51), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n788), .B1(new_n1094), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n248), .A2(new_n1023), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n790), .B1(new_n717), .B2(G97), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n778), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1103), .B(new_n1106), .C1(new_n969), .C2(new_n844), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1015), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n718), .B1(new_n1108), .B2(new_n1078), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1015), .B1(new_n769), .B2(new_n1017), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1107), .B1(new_n1003), .B2(new_n1108), .C1(new_n1109), .C2(new_n1110), .ZN(G390));
  AOI21_X1  g0911(.A(new_n778), .B1(new_n280), .B2(new_n860), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n823), .A2(new_n281), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT53), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n813), .A2(G125), .ZN(new_n1115));
  INV_X1    g0915(.A(G132), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT54), .B(G143), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n1115), .B1(new_n1116), .B2(new_n810), .C1(new_n794), .C2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(G128), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n306), .B1(new_n816), .B2(new_n213), .C1(new_n837), .C2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n806), .A2(G137), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n834), .B2(new_n797), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n1118), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n314), .B1(new_n816), .B2(new_n226), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n866), .A2(new_n454), .B1(new_n837), .B2(new_n867), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1124), .B(new_n1125), .C1(G77), .C2(new_n1027), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(G116), .A2(new_n811), .B1(new_n871), .B2(G97), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n798), .B2(new_n812), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G87), .B2(new_n824), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1114), .A2(new_n1123), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1112), .B1(new_n1130), .B2(new_n862), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n945), .B1(new_n948), .B2(KEYINPUT39), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1131), .B1(new_n1132), .B2(new_n785), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n912), .B1(new_n911), .B2(KEYINPUT38), .ZN(new_n1134));
  NOR4_X1   g0934(.A1(new_n906), .A2(new_n910), .A3(KEYINPUT106), .A4(new_n918), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n919), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n850), .A2(new_n467), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n849), .B1(new_n744), .B2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1136), .B(new_n946), .C1(new_n1138), .C2(new_n932), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n945), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT39), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1140), .B1(new_n1136), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n951), .A2(new_n947), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1139), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n765), .A2(G330), .A3(new_n851), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1145), .A2(new_n932), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1145), .A2(new_n932), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1139), .B(new_n1148), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1147), .A2(new_n776), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(KEYINPUT118), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT118), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1147), .A2(new_n1152), .A3(new_n776), .A4(new_n1149), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1133), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n849), .B1(new_n732), .B2(new_n851), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1145), .A2(new_n932), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1157), .B1(new_n1159), .B2(new_n1146), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1148), .A2(new_n1138), .A3(new_n1158), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n766), .A2(new_n475), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n954), .A2(new_n694), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n719), .B1(new_n1155), .B2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n954), .A2(new_n694), .A3(new_n1163), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1168), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1169));
  AOI21_X1  g0969(.A(KEYINPUT117), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1149), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n946), .B1(new_n1156), .B2(new_n932), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1132), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1148), .B1(new_n1173), .B2(new_n1139), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1165), .B1(new_n1171), .B2(new_n1174), .ZN(new_n1175));
  AND4_X1   g0975(.A1(KEYINPUT117), .A2(new_n1175), .A3(new_n718), .A4(new_n1169), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1154), .B1(new_n1170), .B2(new_n1176), .ZN(G378));
  NAND3_X1  g0977(.A1(new_n687), .A2(new_n473), .A3(new_n688), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(KEYINPUT122), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT122), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n687), .A2(new_n1180), .A3(new_n473), .A4(new_n688), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n699), .B1(new_n279), .B2(new_n287), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT55), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1183), .B(new_n1184), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1179), .A2(new_n1181), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1185), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n940), .B2(G330), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1136), .A2(new_n933), .A3(KEYINPUT40), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n939), .A2(new_n893), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(G330), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1185), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1179), .A2(new_n1181), .A3(new_n1185), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1192), .A2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n953), .B1(new_n1189), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT123), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n940), .A2(G330), .A3(new_n1188), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n953), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1192), .A2(new_n1197), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1199), .A2(new_n1200), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1169), .A2(new_n1164), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .A4(KEYINPUT123), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT57), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1209), .B1(new_n1169), .B2(new_n1164), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1199), .A2(new_n1204), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n719), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1205), .A2(new_n776), .A3(new_n1207), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n860), .A2(new_n213), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n777), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(G137), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n810), .A2(new_n1119), .B1(new_n794), .B2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G132), .B2(new_n806), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1027), .A2(G150), .B1(G125), .B2(new_n801), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(new_n823), .C2(new_n1117), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n282), .B(new_n294), .C1(new_n816), .C2(new_n834), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G124), .B2(new_n813), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1227), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n837), .A2(new_n592), .B1(new_n797), .B2(new_n226), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT119), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n823), .A2(new_n373), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n813), .A2(G283), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1232), .B1(new_n219), .B2(new_n816), .C1(new_n458), .C2(new_n794), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n306), .A2(G41), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n454), .B2(new_n810), .C1(new_n866), .C2(new_n221), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(new_n1230), .A2(new_n1231), .A3(new_n1233), .A4(new_n1235), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1236), .A2(KEYINPUT58), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(KEYINPUT58), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1234), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1239), .B(new_n213), .C1(G33), .C2(G41), .ZN(new_n1240));
  AND4_X1   g1040(.A1(new_n1228), .A2(new_n1237), .A3(new_n1238), .A4(new_n1240), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1217), .B1(new_n862), .B2(new_n1241), .C1(new_n1188), .C2(new_n786), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1215), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1214), .A2(new_n1243), .ZN(G375));
  NAND2_X1  g1044(.A1(new_n1162), .A2(new_n776), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n794), .A2(new_n281), .B1(new_n812), .B2(new_n1119), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n314), .B(new_n1246), .C1(G58), .C2(new_n817), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n824), .A2(G159), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n1116), .A2(new_n837), .B1(new_n866), .B2(new_n1117), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(G50), .B2(new_n1027), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n832), .A2(G137), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1247), .A2(new_n1248), .A3(new_n1250), .A4(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n824), .A2(G97), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n306), .B(new_n1057), .C1(G77), .C2(new_n817), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n806), .A2(G116), .B1(new_n801), .B2(G294), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n810), .A2(new_n867), .B1(new_n794), .B2(new_n454), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(G303), .B2(new_n813), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .A4(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n862), .B1(new_n1252), .B2(new_n1258), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n778), .B(new_n1259), .C1(new_n226), .C2(new_n860), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n938), .B2(new_n786), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1245), .A2(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1168), .A2(new_n1019), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1167), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1262), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(G381));
  NOR4_X1   g1066(.A1(G390), .A2(G384), .A3(G396), .A4(G393), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1265), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1154), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  OR4_X1    g1071(.A1(G387), .A2(new_n1268), .A3(G375), .A4(new_n1271), .ZN(G407));
  INV_X1    g1072(.A(G213), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1273), .A2(G343), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1270), .A2(new_n1274), .ZN(new_n1275));
  OAI211_X1 g1075(.A(G407), .B(G213), .C1(G375), .C2(new_n1275), .ZN(G409));
  NAND3_X1  g1076(.A1(new_n1214), .A2(G378), .A3(new_n1243), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1212), .A2(new_n776), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1242), .B(new_n1278), .C1(new_n1208), .C2(new_n1019), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1270), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1277), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1274), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1165), .A2(KEYINPUT60), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1264), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n719), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1165), .A2(KEYINPUT60), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1264), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1262), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1288), .A2(G384), .ZN(new_n1289));
  AOI211_X1 g1089(.A(new_n1262), .B(new_n882), .C1(new_n1285), .C2(new_n1287), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1281), .A2(KEYINPUT63), .A3(new_n1282), .A4(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT125), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1274), .B1(new_n1277), .B2(new_n1280), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT125), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1294), .A2(new_n1295), .A3(KEYINPUT63), .A4(new_n1291), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1293), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1274), .A2(G2897), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1300), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n718), .B1(new_n1286), .B2(new_n1264), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1302), .B1(new_n1264), .B2(new_n1286), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n882), .B1(new_n1303), .B2(new_n1262), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1288), .A2(G384), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1304), .A2(new_n1305), .A3(new_n1299), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1301), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1298), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(G390), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT124), .B1(G387), .B2(new_n1310), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(G393), .B(new_n846), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1021), .A2(G390), .A3(new_n1045), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(G390), .B1(new_n1021), .B2(new_n1045), .ZN(new_n1316));
  OAI22_X1  g1116(.A1(new_n1311), .A2(new_n1313), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT61), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1316), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1319), .A2(KEYINPUT124), .A3(new_n1312), .A4(new_n1314), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1317), .A2(new_n1318), .A3(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1281), .A2(new_n1282), .A3(new_n1291), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n1309), .B(new_n1321), .C1(new_n1323), .C2(KEYINPUT63), .ZN(new_n1324));
  XOR2_X1   g1124(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1325));
  OAI21_X1  g1125(.A(new_n1325), .B1(new_n1294), .B2(new_n1307), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT62), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1322), .A2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1294), .A2(KEYINPUT62), .A3(new_n1291), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1326), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1317), .A2(new_n1320), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT127), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1317), .A2(KEYINPUT127), .A3(new_n1320), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  OAI22_X1  g1135(.A1(new_n1297), .A2(new_n1324), .B1(new_n1330), .B2(new_n1335), .ZN(G405));
  NAND2_X1  g1136(.A1(G375), .A2(new_n1270), .ZN(new_n1337));
  OAI211_X1 g1137(.A(new_n1337), .B(new_n1277), .C1(new_n1289), .C2(new_n1290), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1271), .B1(new_n1214), .B2(new_n1243), .ZN(new_n1339));
  AND3_X1   g1139(.A1(new_n1214), .A2(G378), .A3(new_n1243), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1291), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1338), .A2(new_n1341), .ZN(new_n1342));
  XNOR2_X1  g1142(.A(new_n1342), .B(new_n1331), .ZN(G402));
endmodule


