//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n540, new_n542, new_n543, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n609, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT66), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT67), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n460), .A2(G137), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n462), .B(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n466), .A2(G2105), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n472), .A2(G2105), .B1(G101), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n464), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  OAI21_X1  g051(.A(G2104), .B1(new_n461), .B2(G112), .ZN(new_n477));
  INV_X1    g052(.A(G100), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(new_n461), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT69), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n470), .A2(new_n461), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n470), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  NAND4_X1  g061(.A1(new_n467), .A2(new_n469), .A3(KEYINPUT4), .A4(G138), .ZN(new_n487));
  NAND2_X1  g062(.A1(G102), .A2(G2104), .ZN(new_n488));
  AOI21_X1  g063(.A(G2105), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(G114), .A2(G2104), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(new_n460), .B2(G126), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT4), .B1(new_n492), .B2(new_n461), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n460), .A2(G138), .A3(new_n461), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n489), .B1(new_n493), .B2(new_n494), .ZN(G164));
  INV_X1    g070(.A(KEYINPUT6), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT70), .B1(new_n496), .B2(G651), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n498));
  INV_X1    g073(.A(G651), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT6), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n497), .A2(new_n500), .B1(new_n496), .B2(G651), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n501), .A2(G88), .B1(G62), .B2(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n504), .A2(new_n510), .ZN(G166));
  XNOR2_X1  g086(.A(KEYINPUT71), .B(G89), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n501), .A2(new_n512), .B1(G63), .B2(G651), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n513), .A2(new_n509), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n501), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G51), .ZN(new_n517));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT7), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n514), .A2(new_n517), .A3(new_n519), .ZN(G286));
  INV_X1    g095(.A(G286), .ZN(G168));
  AND2_X1   g096(.A1(new_n506), .A2(new_n508), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n523), .A2(new_n499), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n501), .A2(new_n522), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G90), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n516), .A2(G52), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n524), .A2(new_n527), .A3(new_n528), .ZN(G301));
  INV_X1    g104(.A(G301), .ZN(G171));
  INV_X1    g105(.A(G43), .ZN(new_n531));
  INV_X1    g106(.A(G81), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n531), .A2(new_n515), .B1(new_n525), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT72), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n499), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G860), .ZN(G153));
  AND3_X1   g114(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G36), .ZN(G176));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT8), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n540), .A2(new_n543), .ZN(G188));
  NAND2_X1  g119(.A1(new_n522), .A2(KEYINPUT75), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT75), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n509), .A2(new_n546), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT76), .B(G65), .Z(new_n548));
  NAND3_X1  g123(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(G78), .A2(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n551), .A2(G651), .B1(G91), .B2(new_n526), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT9), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(KEYINPUT73), .ZN(new_n554));
  INV_X1    g129(.A(G53), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n515), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT74), .ZN(new_n557));
  INV_X1    g132(.A(new_n554), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n501), .A2(G53), .A3(G543), .A4(new_n558), .ZN(new_n559));
  AND3_X1   g134(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n557), .B1(new_n556), .B2(new_n559), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n552), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g139(.A(KEYINPUT77), .B(new_n552), .C1(new_n560), .C2(new_n561), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G299));
  OR2_X1    g142(.A1(new_n504), .A2(new_n510), .ZN(G303));
  NAND2_X1  g143(.A1(new_n516), .A2(G49), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n526), .A2(G87), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT78), .ZN(new_n574));
  AND3_X1   g149(.A1(new_n506), .A2(new_n508), .A3(G61), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n501), .A2(G86), .A3(new_n522), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n501), .A2(G48), .A3(G543), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G305));
  INV_X1    g154(.A(G47), .ZN(new_n580));
  INV_X1    g155(.A(G85), .ZN(new_n581));
  OAI22_X1  g156(.A1(new_n580), .A2(new_n515), .B1(new_n525), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n582), .B(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(G72), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G60), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n509), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G651), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  AND3_X1   g165(.A1(new_n545), .A2(G66), .A3(new_n547), .ZN(new_n591));
  INV_X1    g166(.A(G79), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n503), .ZN(new_n593));
  OAI21_X1  g168(.A(KEYINPUT80), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n545), .A2(G66), .A3(new_n547), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n596));
  OAI211_X1 g171(.A(new_n595), .B(new_n596), .C1(new_n592), .C2(new_n503), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n594), .A2(G651), .A3(new_n597), .ZN(new_n598));
  AND3_X1   g173(.A1(new_n501), .A2(G92), .A3(new_n522), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT10), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n516), .A2(G54), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n598), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n590), .B1(new_n603), .B2(G868), .ZN(G284));
  OAI21_X1  g179(.A(new_n590), .B1(new_n603), .B2(G868), .ZN(G321));
  NAND2_X1  g180(.A1(G286), .A2(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n566), .B2(G868), .ZN(G280));
  XNOR2_X1  g182(.A(G280), .B(KEYINPUT81), .ZN(G297));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n603), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n603), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n538), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT82), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n460), .A2(new_n473), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(G2100), .Z(new_n619));
  NAND2_X1  g194(.A1(new_n481), .A2(G123), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n483), .A2(G135), .ZN(new_n621));
  NOR2_X1   g196(.A1(G99), .A2(G2105), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(new_n461), .B2(G111), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n620), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2096), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n619), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT83), .ZN(G156));
  XNOR2_X1  g202(.A(G1341), .B(G1348), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT15), .B(G2435), .Z(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT87), .B(KEYINPUT88), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT86), .B(G2438), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(KEYINPUT14), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT85), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2451), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2454), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n637), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n642), .A2(new_n644), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n629), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n642), .A2(new_n644), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n649), .A2(new_n628), .A3(new_n645), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n648), .A2(G14), .A3(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n653), .B1(new_n657), .B2(KEYINPUT18), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2096), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2100), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n657), .A2(KEYINPUT17), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n655), .A2(new_n656), .ZN(new_n662));
  AOI21_X1  g237(.A(KEYINPUT18), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n660), .B(new_n663), .Z(G227));
  XNOR2_X1  g239(.A(G1971), .B(G1976), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n670), .A2(KEYINPUT89), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(KEYINPUT89), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n667), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT20), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n668), .A2(new_n669), .ZN(new_n675));
  AOI22_X1  g250(.A1(new_n673), .A2(new_n674), .B1(new_n667), .B2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n675), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n677), .A2(new_n666), .A3(new_n670), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n676), .B(new_n678), .C1(new_n674), .C2(new_n673), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT21), .B(G1986), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT22), .B(G1981), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G229));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n686), .A2(G4), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n602), .B2(G16), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT92), .B(G1348), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n691), .A2(G35), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(new_n485), .B2(G29), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT29), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI211_X1 g270(.A(KEYINPUT29), .B(new_n692), .C1(new_n485), .C2(G29), .ZN(new_n696));
  OAI21_X1  g271(.A(G2090), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT99), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI211_X1 g274(.A(KEYINPUT99), .B(G2090), .C1(new_n695), .C2(new_n696), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(G16), .A2(G21), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G286), .B2(new_n686), .ZN(new_n703));
  INV_X1    g278(.A(G1966), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT97), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n690), .A2(new_n701), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(G171), .A2(G16), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G5), .B2(G16), .ZN(new_n710));
  INV_X1    g285(.A(G1961), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n691), .A2(G27), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G164), .B2(new_n691), .ZN(new_n714));
  MUX2_X1   g289(.A(new_n713), .B(new_n714), .S(KEYINPUT98), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G2078), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n686), .A2(G20), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT23), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n566), .B2(new_n686), .ZN(new_n719));
  INV_X1    g294(.A(G1956), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n708), .A2(new_n712), .A3(new_n716), .A4(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G19), .ZN(new_n723));
  OAI21_X1  g298(.A(KEYINPUT93), .B1(new_n723), .B2(G16), .ZN(new_n724));
  OR3_X1    g299(.A1(new_n723), .A2(KEYINPUT93), .A3(G16), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n724), .B(new_n725), .C1(new_n538), .C2(new_n686), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G1341), .ZN(new_n727));
  NOR3_X1   g302(.A1(new_n695), .A2(new_n696), .A3(G2090), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT28), .ZN(new_n729));
  INV_X1    g304(.A(G26), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(G29), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n730), .A2(G29), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n481), .A2(G128), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n483), .A2(G140), .ZN(new_n734));
  NOR2_X1   g309(.A1(G104), .A2(G2105), .ZN(new_n735));
  OAI21_X1  g310(.A(G2104), .B1(new_n461), .B2(G116), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n733), .B(new_n734), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n732), .B1(new_n737), .B2(G29), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n731), .B1(new_n738), .B2(new_n729), .ZN(new_n739));
  INV_X1    g314(.A(G2067), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  AOI22_X1  g316(.A1(G129), .A2(new_n481), .B1(new_n483), .B2(G141), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n473), .A2(G105), .ZN(new_n743));
  NAND3_X1  g318(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT26), .Z(new_n745));
  NAND3_X1  g320(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  MUX2_X1   g321(.A(G32), .B(new_n746), .S(G29), .Z(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT27), .B(G1996), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT95), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n747), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n741), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT94), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G29), .B2(G33), .ZN(new_n753));
  OR3_X1    g328(.A1(new_n752), .A2(G29), .A3(G33), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n473), .A2(G103), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT25), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n483), .A2(G139), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n757), .B(new_n758), .C1(new_n461), .C2(new_n759), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n753), .B(new_n754), .C1(new_n760), .C2(new_n691), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G2072), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT30), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(G28), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(G28), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n764), .A2(new_n765), .A3(new_n691), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n762), .B(new_n766), .C1(new_n715), .C2(G2078), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n751), .A2(new_n767), .ZN(new_n768));
  OR2_X1    g343(.A1(KEYINPUT24), .A2(G34), .ZN(new_n769));
  NAND2_X1  g344(.A1(KEYINPUT24), .A2(G34), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n769), .A2(new_n691), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G160), .B2(new_n691), .ZN(new_n772));
  INV_X1    g347(.A(G2084), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n768), .B(new_n774), .C1(new_n691), .C2(new_n624), .ZN(new_n775));
  NOR4_X1   g350(.A1(new_n722), .A2(new_n727), .A3(new_n728), .A4(new_n775), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n703), .A2(new_n704), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT96), .Z(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT31), .B(G11), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n710), .A2(new_n711), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n776), .A2(new_n778), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n686), .A2(G22), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G166), .B2(new_n686), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(G1971), .Z(new_n784));
  NOR2_X1   g359(.A1(G16), .A2(G23), .ZN(new_n785));
  AND3_X1   g360(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT33), .B(G1976), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n686), .A2(G6), .ZN(new_n790));
  INV_X1    g365(.A(G305), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(new_n686), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT32), .B(G1981), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n784), .A2(new_n789), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT91), .B(KEYINPUT34), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n686), .A2(G24), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n582), .A2(new_n583), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n582), .A2(new_n583), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n799), .A2(new_n800), .B1(G651), .B2(new_n587), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n798), .B1(new_n801), .B2(new_n686), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT90), .B(G1986), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n691), .A2(G25), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n481), .A2(G119), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n483), .A2(G131), .ZN(new_n807));
  OR2_X1    g382(.A1(G95), .A2(G2105), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n808), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n806), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n805), .B1(new_n811), .B2(new_n691), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT35), .B(G1991), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n812), .B(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n797), .A2(new_n804), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT36), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n781), .A2(new_n818), .ZN(G311));
  AND3_X1   g394(.A1(new_n776), .A2(new_n779), .A3(new_n780), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n820), .A2(KEYINPUT100), .A3(new_n817), .A4(new_n778), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT100), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n781), .B2(new_n818), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n823), .ZN(G150));
  NAND2_X1  g399(.A1(G80), .A2(G543), .ZN(new_n825));
  INV_X1    g400(.A(G67), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n509), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT101), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(G651), .ZN(new_n829));
  AOI22_X1  g404(.A1(G55), .A2(new_n516), .B1(new_n526), .B2(G93), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT102), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G860), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT37), .Z(new_n835));
  NAND2_X1  g410(.A1(new_n538), .A2(new_n831), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n833), .B2(new_n538), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n602), .A2(new_n609), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n835), .B1(new_n841), .B2(G860), .ZN(G145));
  NAND3_X1  g417(.A1(new_n467), .A2(new_n469), .A3(G126), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n461), .B1(new_n843), .B2(new_n490), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT4), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n494), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n489), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n737), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(new_n746), .Z(new_n850));
  AND2_X1   g425(.A1(new_n850), .A2(new_n760), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n760), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n481), .A2(G130), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n483), .A2(G142), .ZN(new_n854));
  NOR2_X1   g429(.A1(G106), .A2(G2105), .ZN(new_n855));
  OAI21_X1  g430(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n853), .B(new_n854), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n617), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n858), .A2(new_n811), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n811), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT103), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n861), .A2(new_n862), .ZN(new_n865));
  OAI22_X1  g440(.A1(new_n851), .A2(new_n852), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n475), .B(new_n624), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n850), .A2(new_n760), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n850), .A2(new_n760), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n869), .A2(new_n863), .A3(new_n870), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n866), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n868), .B1(new_n866), .B2(new_n871), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n485), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n866), .A2(new_n871), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n867), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n866), .A2(new_n871), .A3(new_n868), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n876), .A2(G162), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(G37), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n874), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g456(.A1(G303), .A2(new_n786), .ZN(new_n882));
  NAND2_X1  g457(.A1(G166), .A2(G288), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n801), .ZN(new_n885));
  NAND3_X1  g460(.A1(G290), .A2(new_n883), .A3(new_n882), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(G305), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(new_n886), .A3(new_n791), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT42), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n892), .A2(KEYINPUT106), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(KEYINPUT106), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(new_n894), .B2(new_n891), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n556), .A2(new_n559), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT74), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT77), .B1(new_n900), .B2(new_n552), .ZN(new_n901));
  INV_X1    g476(.A(new_n565), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n602), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n603), .A2(new_n564), .A3(new_n565), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n905), .A2(KEYINPUT104), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(KEYINPUT104), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n837), .B(new_n611), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n903), .A2(KEYINPUT41), .A3(new_n904), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n903), .A2(KEYINPUT105), .A3(new_n904), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n566), .A2(new_n913), .A3(new_n602), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT41), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n912), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n909), .A2(new_n911), .A3(new_n916), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n896), .A2(new_n910), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n896), .B1(new_n910), .B2(new_n917), .ZN(new_n919));
  OAI21_X1  g494(.A(G868), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n833), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n920), .B1(G868), .B2(new_n921), .ZN(G295));
  OAI21_X1  g497(.A(new_n920), .B1(G868), .B2(new_n921), .ZN(G331));
  NAND2_X1  g498(.A1(new_n912), .A2(new_n914), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT41), .ZN(new_n925));
  XNOR2_X1  g500(.A(G286), .B(G301), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n836), .B(new_n926), .C1(new_n538), .C2(new_n833), .ZN(new_n927));
  INV_X1    g502(.A(new_n926), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n829), .A2(new_n830), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n832), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n831), .A2(KEYINPUT102), .ZN(new_n931));
  AOI22_X1  g506(.A1(new_n930), .A2(new_n931), .B1(new_n536), .B2(new_n534), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n537), .A2(new_n929), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n928), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n927), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n905), .A2(new_n915), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n925), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n888), .A2(KEYINPUT107), .A3(new_n889), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT107), .B1(new_n888), .B2(new_n889), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n906), .A2(new_n907), .A3(new_n927), .A4(new_n934), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n937), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n916), .A2(new_n935), .A3(new_n911), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n927), .A2(new_n934), .A3(new_n903), .A4(new_n904), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n890), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n942), .A2(new_n946), .A3(new_n947), .A4(new_n879), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT108), .ZN(new_n949));
  AOI21_X1  g524(.A(G37), .B1(new_n945), .B2(new_n890), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n940), .A2(new_n944), .A3(new_n943), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n950), .A2(new_n954), .A3(new_n947), .A4(new_n942), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n949), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n950), .A2(KEYINPUT43), .A3(new_n942), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT43), .B1(new_n950), .B2(new_n951), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT44), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n958), .A2(new_n961), .ZN(G397));
  NAND3_X1  g537(.A1(new_n464), .A2(G40), .A3(new_n474), .ZN(new_n963));
  AOI21_X1  g538(.A(G1384), .B1(new_n846), .B2(new_n847), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n963), .A2(new_n964), .A3(KEYINPUT45), .ZN(new_n965));
  OR2_X1    g540(.A1(G290), .A2(G1986), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n810), .A2(new_n813), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n811), .A2(new_n814), .ZN(new_n968));
  INV_X1    g543(.A(G1996), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n746), .B(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n737), .B(new_n740), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n966), .A2(new_n967), .A3(new_n968), .A4(new_n973), .ZN(new_n974));
  AND2_X1   g549(.A1(G290), .A2(G1986), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n965), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n978));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n978), .B1(new_n848), .B2(new_n979), .ZN(new_n980));
  AOI211_X1 g555(.A(KEYINPUT111), .B(G1384), .C1(new_n846), .C2(new_n847), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n977), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n964), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n963), .B1(new_n983), .B2(KEYINPUT50), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n982), .A2(new_n773), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT119), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT111), .B1(G164), .B2(G1384), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n848), .A2(new_n978), .A3(new_n979), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n963), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n964), .A2(KEYINPUT45), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n704), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT119), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n982), .A2(new_n995), .A3(new_n984), .A4(new_n773), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n986), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(G8), .ZN(new_n998));
  NAND2_X1  g573(.A1(G286), .A2(G8), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT122), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n999), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT122), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n998), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n1001), .B(G8), .C1(new_n997), .C2(G286), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n997), .A2(new_n1003), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT62), .ZN(new_n1009));
  XOR2_X1   g584(.A(KEYINPUT112), .B(G1981), .Z(new_n1010));
  NAND4_X1  g585(.A1(new_n576), .A2(new_n577), .A3(new_n578), .A4(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT49), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT115), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT113), .B(G86), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n501), .A2(new_n522), .A3(new_n1016), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n578), .A2(new_n1017), .A3(KEYINPUT114), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT114), .B1(new_n578), .B2(new_n1017), .ZN(new_n1019));
  INV_X1    g594(.A(new_n576), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1981), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1015), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1012), .A2(KEYINPUT115), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G8), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n987), .A2(new_n989), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1027), .B1(new_n1028), .B2(new_n991), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1024), .B(new_n1015), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1026), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1026), .A2(new_n1029), .A3(KEYINPUT116), .A4(new_n1030), .ZN(new_n1034));
  INV_X1    g609(.A(G1976), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1029), .B1(new_n1035), .B2(G288), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1033), .A2(new_n1034), .B1(new_n1036), .B2(KEYINPUT52), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n964), .A2(new_n977), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n991), .B(new_n1038), .C1(new_n1028), .C2(new_n977), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1039), .A2(G2090), .ZN(new_n1040));
  XOR2_X1   g615(.A(KEYINPUT110), .B(G1971), .Z(new_n1041));
  NOR3_X1   g616(.A1(G164), .A2(new_n988), .A3(G1384), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT109), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n963), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1043), .B1(new_n964), .B2(KEYINPUT45), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n992), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1041), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(G8), .B1(new_n1040), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(G303), .A2(G8), .ZN(new_n1049));
  XOR2_X1   g624(.A(new_n1049), .B(KEYINPUT55), .Z(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n982), .A2(new_n984), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(G2090), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1050), .B(G8), .C1(new_n1054), .C2(new_n1047), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n786), .A2(G1976), .ZN(new_n1056));
  OR3_X1    g631(.A1(new_n1036), .A2(KEYINPUT52), .A3(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1037), .A2(new_n1052), .A3(new_n1055), .A4(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G2078), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1044), .A2(new_n1060), .A3(new_n1046), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1053), .A2(new_n711), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1062), .A2(G2078), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n990), .A2(new_n991), .A3(new_n992), .A4(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(G171), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT62), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1005), .A2(new_n1070), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1009), .A2(new_n1059), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT126), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1068), .B1(new_n1008), .B2(KEYINPUT62), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT126), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1074), .A2(new_n1075), .A3(new_n1059), .A4(new_n1071), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(KEYINPUT120), .A2(KEYINPUT63), .ZN(new_n1078));
  OR2_X1    g653(.A1(KEYINPUT120), .A2(KEYINPUT63), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n998), .A2(G286), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1078), .B(new_n1079), .C1(new_n1058), .C2(new_n1081), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1037), .A2(new_n1057), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT63), .ZN(new_n1084));
  OAI21_X1  g659(.A(G8), .B1(new_n1054), .B2(new_n1047), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n1085), .B2(new_n1051), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1083), .A2(new_n1055), .A3(new_n1080), .A4(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1082), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1055), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1011), .B(KEYINPUT117), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1091));
  NOR2_X1   g666(.A1(G288), .A2(G1976), .ZN(new_n1092));
  XOR2_X1   g667(.A(new_n1092), .B(KEYINPUT118), .Z(new_n1093));
  OAI21_X1  g668(.A(new_n1090), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1089), .A2(new_n1083), .B1(new_n1094), .B2(new_n1029), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT56), .B(G2072), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1044), .A2(new_n1046), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT121), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1039), .A2(new_n720), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT57), .B1(new_n556), .B2(new_n559), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n562), .A2(KEYINPUT57), .B1(new_n552), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1044), .A2(new_n1102), .A3(new_n1046), .A4(new_n1096), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1098), .A2(new_n1099), .A3(new_n1101), .A4(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT61), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1028), .A2(new_n991), .ZN(new_n1106));
  XOR2_X1   g681(.A(KEYINPUT58), .B(G1341), .Z(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1044), .A2(new_n969), .A3(new_n1046), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n537), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1110), .B(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1028), .A2(new_n740), .A3(new_n991), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1053), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1113), .B1(new_n1114), .B2(G1348), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n602), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n603), .B(new_n1113), .C1(new_n1114), .C2(G1348), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(new_n1117), .A3(KEYINPUT60), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n1117), .A2(KEYINPUT60), .ZN(new_n1119));
  AND4_X1   g694(.A1(new_n1105), .A2(new_n1112), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1115), .A2(new_n603), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1098), .A2(new_n1099), .A3(new_n1103), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1121), .B1(new_n1122), .B2(new_n1101), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1123), .A2(new_n1104), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1059), .B1(new_n1120), .B2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1104), .A2(KEYINPUT61), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT53), .B1(new_n1127), .B2(KEYINPUT125), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1061), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1127), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1130), .A2(KEYINPUT125), .A3(KEYINPUT53), .A4(new_n1060), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1064), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1053), .A2(KEYINPUT124), .A3(new_n711), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1129), .A2(new_n1131), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(G171), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1067), .A2(G171), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT54), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1126), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1068), .B1(new_n1135), .B2(G171), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT123), .B(KEYINPUT54), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1140), .A2(new_n1143), .A3(new_n1008), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1088), .B(new_n1095), .C1(new_n1125), .C2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n976), .B1(new_n1077), .B2(new_n1145), .ZN(new_n1146));
  OAI22_X1  g721(.A1(new_n972), .A2(new_n968), .B1(G2067), .B2(new_n737), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1147), .A2(new_n965), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT46), .ZN(new_n1149));
  INV_X1    g724(.A(new_n965), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1149), .B1(new_n1150), .B2(G1996), .ZN(new_n1151));
  INV_X1    g726(.A(new_n971), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n965), .B1(new_n1152), .B2(new_n746), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n965), .A2(KEYINPUT46), .A3(new_n969), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1151), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  XOR2_X1   g730(.A(new_n1155), .B(KEYINPUT47), .Z(new_n1156));
  NOR2_X1   g731(.A1(new_n966), .A2(new_n1150), .ZN(new_n1157));
  XOR2_X1   g732(.A(new_n1157), .B(KEYINPUT48), .Z(new_n1158));
  NAND3_X1  g733(.A1(new_n973), .A2(new_n967), .A3(new_n968), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n965), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT127), .ZN(new_n1161));
  AOI211_X1 g736(.A(new_n1148), .B(new_n1156), .C1(new_n1158), .C2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1146), .A2(new_n1162), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g738(.A(G227), .ZN(new_n1165));
  AND2_X1   g739(.A1(new_n651), .A2(new_n1165), .ZN(new_n1166));
  AND2_X1   g740(.A1(new_n880), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g741(.A(G319), .ZN(new_n1168));
  NOR2_X1   g742(.A1(G229), .A2(new_n1168), .ZN(new_n1169));
  AND3_X1   g743(.A1(new_n1167), .A2(new_n956), .A3(new_n1169), .ZN(G308));
  NAND3_X1  g744(.A1(new_n1167), .A2(new_n956), .A3(new_n1169), .ZN(G225));
endmodule


