//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 0 0 1 0 1 0 0 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023;
  INV_X1    g000(.A(KEYINPUT17), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n203), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n204));
  XOR2_X1   g003(.A(KEYINPUT14), .B(G29gat), .Z(new_n205));
  OAI21_X1  g004(.A(new_n204), .B1(new_n205), .B2(G36gat), .ZN(new_n206));
  XOR2_X1   g005(.A(KEYINPUT89), .B(G43gat), .Z(new_n207));
  INV_X1    g006(.A(G50gat), .ZN(new_n208));
  AND2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G43gat), .A2(G50gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT15), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n206), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G43gat), .A2(G50gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n211), .B1(new_n215), .B2(new_n210), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n206), .A2(new_n216), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n202), .B1(new_n220), .B2(KEYINPUT90), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT90), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n218), .A2(new_n222), .A3(KEYINPUT17), .A4(new_n219), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G15gat), .B(G22gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT16), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(G1gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(KEYINPUT91), .A3(G8gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n225), .A2(G1gat), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(G8gat), .B1(new_n227), .B2(KEYINPUT92), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(KEYINPUT92), .B2(new_n227), .ZN(new_n232));
  NAND2_X1  g031(.A1(KEYINPUT91), .A2(G8gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n224), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n235), .A2(new_n220), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G229gat), .A2(G233gat), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n236), .A2(KEYINPUT18), .A3(new_n238), .A4(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n235), .B(new_n220), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n239), .B(KEYINPUT13), .Z(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n236), .A2(new_n238), .A3(new_n239), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT18), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT93), .ZN(new_n248));
  XNOR2_X1  g047(.A(G113gat), .B(G141gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(G197gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT11), .B(G169gat), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n250), .B(new_n251), .Z(new_n252));
  XOR2_X1   g051(.A(new_n252), .B(KEYINPUT12), .Z(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n244), .B(new_n247), .C1(new_n248), .C2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n240), .A2(new_n248), .A3(new_n243), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n243), .ZN(new_n257));
  INV_X1    g056(.A(new_n235), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n258), .B1(new_n221), .B2(new_n223), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n259), .A2(new_n237), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT18), .B1(new_n260), .B2(new_n239), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n256), .B(new_n253), .C1(new_n257), .C2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT36), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT67), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT27), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n267), .A2(G183gat), .ZN(new_n268));
  INV_X1    g067(.A(G183gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n269), .A2(KEYINPUT27), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n266), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(KEYINPUT27), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n267), .A2(G183gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n272), .A2(new_n273), .A3(KEYINPUT67), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT28), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(G190gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n271), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G190gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n272), .A2(new_n273), .A3(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n275), .B1(new_n279), .B2(KEYINPUT66), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT66), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT27), .B(G183gat), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n281), .B1(new_n282), .B2(new_n278), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n277), .B1(new_n280), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT26), .ZN(new_n287));
  NAND2_X1  g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n285), .A2(KEYINPUT26), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n284), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT25), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT23), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n296), .B1(new_n285), .B2(KEYINPUT65), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT65), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n298), .B(KEYINPUT23), .C1(G169gat), .C2(G176gat), .ZN(new_n299));
  AND2_X1   g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT24), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(G183gat), .A3(G190gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n290), .A2(KEYINPUT24), .ZN(new_n303));
  NOR2_X1   g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n288), .B(new_n302), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n295), .B1(new_n300), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n288), .B1(new_n290), .B2(KEYINPUT24), .ZN(new_n307));
  INV_X1    g106(.A(new_n303), .ZN(new_n308));
  INV_X1    g107(.A(new_n304), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n297), .A2(new_n299), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(KEYINPUT25), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n294), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G120gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G113gat), .ZN(new_n316));
  INV_X1    g115(.A(G113gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G120gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320));
  XNOR2_X1  g119(.A(G127gat), .B(G134gat), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n319), .B(new_n320), .C1(new_n321), .C2(KEYINPUT68), .ZN(new_n322));
  INV_X1    g121(.A(G127gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G134gat), .ZN(new_n324));
  INV_X1    g123(.A(G134gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G127gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n320), .A2(KEYINPUT68), .ZN(new_n328));
  XNOR2_X1  g127(.A(G113gat), .B(G120gat), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n327), .B(new_n328), .C1(new_n329), .C2(KEYINPUT1), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n322), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G227gat), .A2(G233gat), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n333), .B(KEYINPUT64), .Z(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n284), .A2(new_n293), .B1(new_n306), .B2(new_n312), .ZN(new_n336));
  INV_X1    g135(.A(new_n331), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n332), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT34), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT34), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n332), .A2(new_n338), .A3(new_n341), .A4(new_n335), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(KEYINPUT69), .B(G71gat), .Z(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(G99gat), .ZN(new_n345));
  XOR2_X1   g144(.A(G15gat), .B(G43gat), .Z(new_n346));
  XOR2_X1   g145(.A(new_n345), .B(new_n346), .Z(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n314), .A2(new_n331), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n336), .A2(new_n337), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n334), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT33), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n348), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n343), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n335), .B1(new_n332), .B2(new_n338), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n347), .B1(new_n355), .B2(KEYINPUT33), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n356), .A2(new_n340), .A3(new_n342), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n351), .A2(KEYINPUT32), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n354), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n359), .B1(new_n354), .B2(new_n357), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n265), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n354), .A2(new_n357), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n358), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n354), .A2(new_n357), .A3(new_n359), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(KEYINPUT36), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT31), .B(G50gat), .ZN(new_n369));
  INV_X1    g168(.A(G106gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G155gat), .A2(G162gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT2), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT74), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n373), .A2(KEYINPUT74), .A3(KEYINPUT2), .ZN(new_n377));
  AND2_X1   g176(.A1(G141gat), .A2(G148gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(G141gat), .A2(G148gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n376), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G155gat), .B(G162gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT75), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n385), .B1(new_n373), .B2(KEYINPUT2), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n373), .A2(new_n385), .A3(KEYINPUT2), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n387), .A2(new_n380), .A3(new_n382), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT3), .ZN(new_n391));
  AND2_X1   g190(.A1(G211gat), .A2(G218gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(G211gat), .A2(G218gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(G197gat), .A2(G204gat), .ZN(new_n395));
  NOR2_X1   g194(.A1(G197gat), .A2(G204gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G211gat), .B(G218gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(G197gat), .B(G204gat), .ZN(new_n401));
  INV_X1    g200(.A(new_n398), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT29), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT79), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n391), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI211_X1 g205(.A(KEYINPUT79), .B(KEYINPUT29), .C1(new_n399), .C2(new_n403), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n390), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT80), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT80), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n410), .B(new_n390), .C1(new_n406), .C2(new_n407), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n399), .A2(new_n403), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n384), .A2(new_n391), .A3(new_n389), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT29), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n409), .A2(new_n411), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(G228gat), .A2(G233gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G22gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n390), .A2(new_n404), .ZN(new_n421));
  XNOR2_X1  g220(.A(G141gat), .B(G148gat), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT74), .B1(new_n373), .B2(KEYINPUT2), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n382), .B1(new_n424), .B2(new_n377), .ZN(new_n425));
  INV_X1    g224(.A(G141gat), .ZN(new_n426));
  INV_X1    g225(.A(G148gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(G141gat), .A2(G148gat), .ZN(new_n429));
  INV_X1    g228(.A(new_n373), .ZN(new_n430));
  NOR2_X1   g229(.A1(G155gat), .A2(G162gat), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n428), .B(new_n429), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n388), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n432), .A2(new_n433), .A3(new_n386), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT3), .B1(new_n425), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n418), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n421), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT81), .B1(new_n413), .B2(new_n414), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n438), .A2(new_n412), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n413), .A2(KEYINPUT81), .A3(new_n414), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n419), .A2(new_n420), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n415), .B1(new_n408), .B2(KEYINPUT80), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n436), .B1(new_n444), .B2(new_n411), .ZN(new_n445));
  OAI21_X1  g244(.A(G22gat), .B1(new_n445), .B2(new_n441), .ZN(new_n446));
  INV_X1    g245(.A(G78gat), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n443), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n447), .B1(new_n443), .B2(new_n446), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n372), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n443), .A2(new_n446), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(G78gat), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n443), .A2(new_n446), .A3(new_n447), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(new_n453), .A3(new_n371), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n435), .A2(new_n331), .A3(new_n413), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n384), .A2(new_n389), .A3(new_n322), .A4(new_n330), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT4), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(G225gat), .A2(G233gat), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n337), .A2(KEYINPUT4), .A3(new_n384), .A4(new_n389), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n456), .A2(new_n459), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT77), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT5), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n331), .B1(new_n425), .B2(new_n434), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT76), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n457), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n460), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n390), .A2(KEYINPUT76), .A3(new_n331), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n465), .A2(KEYINPUT5), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(KEYINPUT5), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(new_n462), .A3(new_n464), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G1gat), .B(G29gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(KEYINPUT0), .ZN(new_n477));
  XNOR2_X1  g276(.A(G57gat), .B(G85gat), .ZN(new_n478));
  XOR2_X1   g277(.A(new_n477), .B(new_n478), .Z(new_n479));
  NAND2_X1  g278(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481));
  INV_X1    g280(.A(new_n479), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n472), .A2(new_n482), .A3(new_n474), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT78), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n483), .A2(new_n481), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT78), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n480), .A2(new_n488), .A3(new_n481), .A4(new_n483), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G8gat), .B(G36gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(G64gat), .B(G92gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n493), .B(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(G226gat), .ZN(new_n496));
  INV_X1    g295(.A(G233gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(new_n336), .B2(KEYINPUT29), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n314), .A2(new_n498), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(new_n412), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT70), .B1(new_n336), .B2(new_n499), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT70), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n300), .A2(new_n295), .A3(new_n305), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT25), .B1(new_n310), .B2(new_n311), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n279), .A2(KEYINPUT66), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n282), .A2(new_n281), .A3(new_n278), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(new_n509), .A3(new_n275), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n292), .B1(new_n510), .B2(new_n277), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n504), .B(new_n498), .C1(new_n507), .C2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n414), .B1(new_n507), .B2(new_n511), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n503), .A2(new_n512), .B1(new_n499), .B2(new_n513), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n495), .B(new_n502), .C1(new_n514), .C2(new_n412), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT30), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n503), .A2(new_n512), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n412), .B1(new_n518), .B2(new_n500), .ZN(new_n519));
  INV_X1    g318(.A(new_n502), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT71), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT71), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n522), .B(new_n502), .C1(new_n514), .C2(new_n412), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n495), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n517), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n490), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n368), .B1(new_n455), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n515), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT37), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n529), .B(new_n502), .C1(new_n514), .C2(new_n412), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n495), .A2(KEYINPUT38), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT86), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n500), .A2(new_n501), .ZN(new_n534));
  INV_X1    g333(.A(new_n412), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n518), .A2(new_n412), .A3(new_n500), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n514), .A2(new_n533), .A3(new_n412), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(KEYINPUT37), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n528), .B1(new_n532), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n483), .A2(KEYINPUT85), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT85), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n472), .A2(new_n474), .A3(new_n543), .A4(new_n482), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n542), .A2(new_n480), .A3(new_n481), .A4(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n541), .A2(new_n545), .A3(new_n487), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT87), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n541), .A2(new_n545), .A3(KEYINPUT87), .A4(new_n487), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT38), .ZN(new_n551));
  INV_X1    g350(.A(new_n530), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n521), .A2(new_n523), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n495), .B1(new_n553), .B2(KEYINPUT37), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n552), .B1(new_n554), .B2(KEYINPUT88), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT88), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n529), .B1(new_n521), .B2(new_n523), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n556), .B1(new_n557), .B2(new_n495), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n551), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n550), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n450), .A2(new_n454), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n542), .A2(new_n544), .ZN(new_n562));
  INV_X1    g361(.A(new_n524), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n515), .B(KEYINPUT30), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT39), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n456), .A2(new_n459), .A3(new_n461), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT82), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n567), .A2(new_n568), .A3(new_n469), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n568), .B1(new_n567), .B2(new_n469), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n566), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n479), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n570), .A2(new_n571), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n468), .A2(new_n470), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n566), .B1(new_n575), .B2(new_n460), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n573), .A2(KEYINPUT83), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT83), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n572), .A2(new_n578), .A3(new_n479), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT84), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT40), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n565), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n469), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT82), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT39), .B1(new_n584), .B2(new_n569), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT83), .B1(new_n585), .B2(new_n482), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n574), .A2(new_n576), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n579), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT84), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n588), .A2(new_n589), .A3(new_n581), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n561), .B1(new_n582), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n527), .B1(new_n560), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n360), .A2(new_n361), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(new_n450), .A3(new_n454), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT35), .B1(new_n526), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT35), .B1(new_n545), .B2(new_n487), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n561), .A2(new_n525), .A3(new_n593), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n264), .B1(new_n592), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n490), .ZN(new_n600));
  XOR2_X1   g399(.A(G134gat), .B(G162gat), .Z(new_n601));
  AND2_X1   g400(.A1(G232gat), .A2(G233gat), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n602), .A2(KEYINPUT41), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n601), .B(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n604), .B(KEYINPUT103), .Z(new_n605));
  INV_X1    g404(.A(KEYINPUT8), .ZN(new_n606));
  NAND2_X1  g405(.A1(G99gat), .A2(G106gat), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT100), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n609), .B1(new_n608), .B2(new_n607), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n611));
  NAND3_X1  g410(.A1(KEYINPUT99), .A2(G85gat), .A3(G92gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g412(.A1(KEYINPUT99), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n610), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  OR2_X1    g414(.A1(G99gat), .A2(G106gat), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(new_n607), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n607), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n610), .A2(new_n618), .A3(new_n613), .A4(new_n614), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT101), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n224), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT102), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT101), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n620), .B(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n220), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n602), .A2(KEYINPUT41), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n622), .A2(new_n623), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n625), .B1(new_n221), .B2(new_n223), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n628), .B1(new_n621), .B2(new_n220), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT102), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G190gat), .B(G218gat), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n629), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n634), .B1(new_n629), .B2(new_n632), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n605), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n629), .A2(new_n632), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n633), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n604), .A2(KEYINPUT103), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n629), .A2(new_n632), .A3(new_n634), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT94), .ZN(new_n644));
  INV_X1    g443(.A(G57gat), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(G64gat), .ZN(new_n646));
  INV_X1    g445(.A(G64gat), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(G57gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G71gat), .A2(G78gat), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT9), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n644), .B1(new_n653), .B2(KEYINPUT95), .ZN(new_n654));
  XNOR2_X1  g453(.A(G71gat), .B(G78gat), .ZN(new_n655));
  AOI22_X1  g454(.A1(new_n646), .A2(new_n648), .B1(new_n651), .B2(new_n650), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n655), .B1(new_n656), .B2(KEYINPUT94), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n644), .B(new_n655), .C1(new_n653), .C2(KEYINPUT95), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT21), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G183gat), .B(G211gat), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n235), .B1(new_n661), .B2(new_n662), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT98), .ZN(new_n671));
  XOR2_X1   g470(.A(G127gat), .B(G155gat), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT97), .ZN(new_n673));
  NAND2_X1  g472(.A1(G231gat), .A2(G233gat), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(KEYINPUT96), .Z(new_n675));
  XNOR2_X1  g474(.A(new_n673), .B(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n671), .A2(new_n676), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n669), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n679), .ZN(new_n681));
  OAI22_X1  g480(.A1(new_n681), .A2(new_n677), .B1(new_n667), .B2(new_n668), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n660), .A2(KEYINPUT10), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n625), .A2(new_n686), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n620), .A2(new_n660), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n620), .A2(new_n660), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT10), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n685), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n625), .A2(new_n686), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n688), .A2(new_n689), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n692), .B(KEYINPUT104), .C1(new_n693), .C2(KEYINPUT10), .ZN(new_n694));
  NAND2_X1  g493(.A1(G230gat), .A2(G233gat), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n691), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(G120gat), .B(G148gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(G176gat), .B(G204gat), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n697), .B(new_n698), .Z(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n695), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n700), .B1(new_n693), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n696), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n693), .A2(new_n701), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n690), .B1(new_n625), .B2(new_n686), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(new_n705), .B2(new_n701), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n700), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n643), .A2(new_n684), .A3(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n599), .A2(new_n600), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(G1gat), .ZN(G1324gat));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n563), .A2(new_n564), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n486), .B1(new_n484), .B2(KEYINPUT78), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n715), .B1(new_n716), .B2(new_n489), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n367), .B1(new_n717), .B2(new_n561), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n553), .A2(KEYINPUT37), .ZN(new_n719));
  INV_X1    g518(.A(new_n495), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n719), .A2(KEYINPUT88), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n721), .A2(new_n558), .A3(new_n530), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(KEYINPUT38), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n548), .A3(new_n549), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n581), .B1(new_n588), .B2(new_n589), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n542), .B(new_n544), .C1(new_n517), .C2(new_n524), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n590), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n455), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n718), .B1(new_n724), .B2(new_n729), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n595), .A2(new_n597), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n263), .B(new_n711), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n714), .B1(new_n732), .B2(new_n525), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n599), .A2(KEYINPUT105), .A3(new_n715), .A4(new_n711), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g534(.A(KEYINPUT16), .B(G8gat), .Z(new_n736));
  AOI21_X1  g535(.A(KEYINPUT42), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n733), .A2(new_n734), .A3(G8gat), .ZN(new_n738));
  INV_X1    g537(.A(new_n732), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n739), .A2(KEYINPUT42), .A3(new_n715), .A4(new_n736), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT106), .B1(new_n737), .B2(new_n741), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(G1325gat));
  OAI21_X1  g545(.A(G15gat), .B1(new_n732), .B2(new_n367), .ZN(new_n747));
  INV_X1    g546(.A(new_n593), .ZN(new_n748));
  OR2_X1    g547(.A1(new_n748), .A2(G15gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n732), .B2(new_n749), .ZN(G1326gat));
  NOR2_X1   g549(.A1(new_n732), .A2(new_n561), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT43), .B(G22gat), .Z(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1327gat));
  NOR3_X1   g552(.A1(new_n643), .A2(new_n684), .A3(new_n708), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n599), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(new_n203), .A3(new_n600), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT45), .ZN(new_n758));
  XOR2_X1   g557(.A(new_n708), .B(KEYINPUT107), .Z(new_n759));
  NOR3_X1   g558(.A1(new_n759), .A2(new_n264), .A3(new_n684), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(KEYINPUT108), .B1(new_n730), .B2(new_n731), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT108), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n592), .A2(new_n763), .A3(new_n598), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n643), .A2(KEYINPUT44), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n762), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n730), .A2(new_n731), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT44), .B1(new_n767), .B2(new_n643), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n761), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n769), .A2(new_n600), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n758), .B1(new_n203), .B2(new_n770), .ZN(G1328gat));
  NOR3_X1   g570(.A1(new_n755), .A2(G36gat), .A3(new_n525), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT46), .ZN(new_n773));
  INV_X1    g572(.A(G36gat), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n769), .A2(new_n715), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(G1329gat));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n593), .A2(new_n207), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n756), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT109), .B1(new_n755), .B2(new_n778), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n769), .A2(new_n368), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n783), .B(KEYINPUT47), .C1(new_n784), .C2(new_n207), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT47), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n207), .B1(new_n769), .B2(new_n368), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n787), .B2(new_n782), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(G1330gat));
  INV_X1    g588(.A(KEYINPUT48), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n766), .A2(new_n768), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n791), .A2(new_n455), .A3(new_n760), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G50gat), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n755), .A2(G50gat), .A3(new_n561), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n790), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  AOI211_X1 g595(.A(KEYINPUT48), .B(new_n794), .C1(new_n792), .C2(G50gat), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n796), .A2(new_n797), .ZN(G1331gat));
  INV_X1    g597(.A(new_n759), .ZN(new_n799));
  INV_X1    g598(.A(new_n643), .ZN(new_n800));
  NOR4_X1   g599(.A1(new_n799), .A2(new_n263), .A3(new_n683), .A4(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n762), .A2(new_n764), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT110), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n762), .A2(new_n764), .A3(KEYINPUT110), .A4(new_n801), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n804), .A2(new_n600), .A3(new_n805), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(G57gat), .ZN(G1332gat));
  NAND3_X1  g606(.A1(new_n804), .A2(new_n715), .A3(new_n805), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n809));
  XOR2_X1   g608(.A(KEYINPUT49), .B(G64gat), .Z(new_n810));
  OAI21_X1  g609(.A(new_n809), .B1(new_n808), .B2(new_n810), .ZN(G1333gat));
  NAND3_X1  g610(.A1(new_n804), .A2(new_n368), .A3(new_n805), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G71gat), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n748), .A2(G71gat), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n804), .A2(new_n805), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n813), .A2(KEYINPUT50), .A3(new_n815), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(G1334gat));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n455), .A3(new_n805), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g621(.A1(new_n264), .A2(new_n683), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n709), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(new_n766), .B2(new_n768), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n826), .A2(new_n600), .ZN(new_n827));
  INV_X1    g626(.A(G85gat), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n592), .A2(new_n598), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n823), .B1(KEYINPUT111), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n829), .A2(new_n800), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n830), .A2(KEYINPUT111), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n833), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n829), .A2(new_n800), .A3(new_n831), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n600), .A2(new_n828), .A3(new_n708), .ZN(new_n838));
  OAI22_X1  g637(.A1(new_n827), .A2(new_n828), .B1(new_n837), .B2(new_n838), .ZN(G1336gat));
  INV_X1    g638(.A(KEYINPUT52), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n799), .A2(G92gat), .A3(new_n525), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n834), .A2(new_n836), .A3(new_n841), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n826), .A2(new_n715), .ZN(new_n843));
  INV_X1    g642(.A(G92gat), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n840), .B(new_n842), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n844), .B1(new_n826), .B2(new_n715), .ZN(new_n846));
  INV_X1    g645(.A(new_n842), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT52), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n845), .A2(new_n848), .ZN(G1337gat));
  OR4_X1    g648(.A1(G99gat), .A2(new_n837), .A3(new_n748), .A4(new_n709), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n826), .A2(new_n368), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT112), .ZN(new_n852));
  OAI21_X1  g651(.A(G99gat), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n826), .A2(new_n852), .A3(new_n368), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n850), .B1(new_n853), .B2(new_n854), .ZN(G1338gat));
  NOR3_X1   g654(.A1(new_n799), .A2(G106gat), .A3(new_n561), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n834), .A2(new_n836), .A3(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT113), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n826), .A2(new_n455), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n859), .B(new_n860), .C1(new_n861), .C2(new_n370), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n370), .B1(new_n826), .B2(new_n455), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n857), .A2(new_n858), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT53), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n862), .A2(new_n865), .ZN(G1339gat));
  NOR2_X1   g665(.A1(new_n710), .A2(new_n263), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n868), .B1(new_n705), .B2(new_n701), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n696), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n868), .B(new_n695), .C1(new_n687), .C2(new_n690), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n700), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT55), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n872), .B1(new_n696), .B2(new_n869), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT55), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n263), .A2(new_n876), .A3(new_n703), .A4(new_n878), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n247), .A2(new_n243), .A3(new_n240), .A4(new_n254), .ZN(new_n880));
  OAI22_X1  g679(.A1(new_n260), .A2(new_n239), .B1(new_n241), .B2(new_n242), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n252), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AOI22_X1  g682(.A1(new_n883), .A2(new_n708), .B1(new_n637), .B2(new_n642), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n684), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  AOI22_X1  g684(.A1(new_n874), .A2(new_n875), .B1(new_n696), .B2(new_n702), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n880), .A2(new_n887), .A3(new_n882), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n880), .A2(new_n882), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT114), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n886), .A2(new_n888), .A3(new_n878), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n800), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n867), .B1(new_n885), .B2(new_n892), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n561), .A2(new_n600), .A3(new_n525), .A4(new_n593), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n263), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(G113gat), .ZN(G1340gat));
  AOI21_X1  g696(.A(G120gat), .B1(new_n895), .B2(new_n708), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n799), .A2(new_n315), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n895), .B2(new_n899), .ZN(G1341gat));
  NAND2_X1  g699(.A1(new_n895), .A2(new_n684), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g701(.A1(new_n895), .A2(new_n800), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(G134gat), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n895), .A2(new_n325), .A3(new_n800), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT115), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n905), .A2(new_n906), .A3(KEYINPUT56), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n905), .B2(KEYINPUT56), .ZN(new_n908));
  OAI221_X1 g707(.A(new_n904), .B1(KEYINPUT56), .B2(new_n905), .C1(new_n907), .C2(new_n908), .ZN(G1343gat));
  NOR3_X1   g708(.A1(new_n368), .A2(new_n715), .A3(new_n490), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n867), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n879), .A2(new_n884), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n683), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n703), .B1(new_n877), .B2(KEYINPUT55), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n870), .A2(KEYINPUT55), .A3(new_n873), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n887), .B1(new_n880), .B2(new_n882), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n643), .B1(new_n918), .B2(new_n888), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n912), .B1(new_n914), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(KEYINPUT57), .A3(new_n455), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT57), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n922), .B1(new_n893), .B2(new_n561), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n911), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n263), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n893), .A2(new_n561), .A3(new_n911), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n264), .A2(G141gat), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n925), .A2(G141gat), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT58), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n928), .B(new_n929), .ZN(G1344gat));
  NAND3_X1  g729(.A1(new_n926), .A2(new_n427), .A3(new_n708), .ZN(new_n931));
  XNOR2_X1  g730(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n932));
  AOI21_X1  g731(.A(KEYINPUT57), .B1(new_n455), .B2(KEYINPUT117), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n934), .B1(new_n920), .B2(new_n455), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n893), .A2(new_n561), .A3(new_n933), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n708), .B(new_n910), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n932), .B1(new_n937), .B2(G148gat), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n427), .A2(KEYINPUT59), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n939), .B1(new_n924), .B2(new_n708), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n931), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT118), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT118), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n943), .B(new_n931), .C1(new_n938), .C2(new_n940), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(G1345gat));
  INV_X1    g744(.A(G155gat), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n946), .B1(new_n924), .B2(new_n684), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n926), .A2(new_n946), .A3(new_n684), .ZN(new_n948));
  OR2_X1    g747(.A1(new_n947), .A2(new_n948), .ZN(G1346gat));
  AOI21_X1  g748(.A(G162gat), .B1(new_n926), .B2(new_n800), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n800), .A2(G162gat), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(new_n924), .B2(new_n951), .ZN(G1347gat));
  NOR2_X1   g751(.A1(new_n594), .A2(new_n525), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT119), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n954), .B1(new_n920), .B2(new_n490), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n893), .A2(KEYINPUT119), .A3(new_n600), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT120), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI211_X1 g758(.A(KEYINPUT120), .B(new_n953), .C1(new_n955), .C2(new_n956), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n264), .A2(G169gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT121), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n490), .A2(new_n715), .ZN(new_n964));
  OR3_X1    g763(.A1(new_n893), .A2(new_n594), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(G169gat), .B1(new_n965), .B2(new_n264), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n962), .A2(new_n963), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n963), .B1(new_n962), .B2(new_n966), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n967), .A2(new_n968), .ZN(G1348gat));
  NOR2_X1   g768(.A1(new_n709), .A2(G176gat), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n959), .A2(new_n960), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g770(.A(G176gat), .B1(new_n965), .B2(new_n799), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1349gat));
  OAI21_X1  g772(.A(G183gat), .B1(new_n965), .B2(new_n683), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n684), .A2(new_n271), .A3(new_n274), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n974), .B1(new_n957), .B2(new_n975), .ZN(new_n976));
  XOR2_X1   g775(.A(KEYINPUT122), .B(KEYINPUT60), .Z(new_n977));
  XNOR2_X1  g776(.A(new_n976), .B(new_n977), .ZN(G1350gat));
  OAI21_X1  g777(.A(G190gat), .B1(new_n965), .B2(new_n643), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(KEYINPUT123), .ZN(new_n980));
  OR2_X1    g779(.A1(new_n980), .A2(KEYINPUT61), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n959), .A2(new_n278), .A3(new_n800), .A4(new_n960), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n979), .A2(KEYINPUT123), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n980), .A2(KEYINPUT61), .ZN(new_n984));
  OAI211_X1 g783(.A(new_n981), .B(new_n982), .C1(new_n983), .C2(new_n984), .ZN(G1351gat));
  XNOR2_X1  g784(.A(KEYINPUT124), .B(G197gat), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n368), .A2(new_n964), .ZN(new_n987));
  INV_X1    g786(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n920), .A2(new_n455), .A3(new_n934), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n933), .B1(new_n893), .B2(new_n561), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n986), .B1(new_n991), .B2(new_n263), .ZN(new_n992));
  NOR3_X1   g791(.A1(new_n368), .A2(new_n561), .A3(new_n525), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n993), .B1(new_n955), .B2(new_n956), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n263), .A2(new_n986), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT125), .ZN(new_n998));
  XNOR2_X1  g797(.A(new_n997), .B(new_n998), .ZN(G1352gat));
  INV_X1    g798(.A(G204gat), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n708), .A2(new_n1000), .ZN(new_n1001));
  OR3_X1    g800(.A1(new_n994), .A2(KEYINPUT62), .A3(new_n1001), .ZN(new_n1002));
  OAI21_X1  g801(.A(KEYINPUT62), .B1(new_n994), .B2(new_n1001), .ZN(new_n1003));
  AND2_X1   g802(.A1(new_n991), .A2(new_n759), .ZN(new_n1004));
  OAI211_X1 g803(.A(new_n1002), .B(new_n1003), .C1(new_n1000), .C2(new_n1004), .ZN(G1353gat));
  INV_X1    g804(.A(G211gat), .ZN(new_n1006));
  AOI211_X1 g805(.A(new_n683), .B(new_n988), .C1(new_n989), .C2(new_n990), .ZN(new_n1007));
  AOI21_X1  g806(.A(new_n1006), .B1(new_n1007), .B2(KEYINPUT126), .ZN(new_n1008));
  AOI21_X1  g807(.A(KEYINPUT126), .B1(new_n991), .B2(new_n684), .ZN(new_n1009));
  INV_X1    g808(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g809(.A(KEYINPUT63), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g810(.A(new_n684), .B(new_n987), .C1(new_n935), .C2(new_n936), .ZN(new_n1012));
  INV_X1    g811(.A(KEYINPUT126), .ZN(new_n1013));
  OAI21_X1  g812(.A(G211gat), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g813(.A(KEYINPUT63), .ZN(new_n1015));
  NOR3_X1   g814(.A1(new_n1014), .A2(new_n1015), .A3(new_n1009), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n684), .A2(new_n1006), .ZN(new_n1017));
  OAI22_X1  g816(.A1(new_n1011), .A2(new_n1016), .B1(new_n994), .B2(new_n1017), .ZN(G1354gat));
  INV_X1    g817(.A(G218gat), .ZN(new_n1019));
  OAI21_X1  g818(.A(new_n1019), .B1(new_n994), .B2(new_n643), .ZN(new_n1020));
  OR2_X1    g819(.A1(new_n1020), .A2(KEYINPUT127), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1020), .A2(KEYINPUT127), .ZN(new_n1022));
  NOR2_X1   g821(.A1(new_n643), .A2(new_n1019), .ZN(new_n1023));
  AOI22_X1  g822(.A1(new_n1021), .A2(new_n1022), .B1(new_n991), .B2(new_n1023), .ZN(G1355gat));
endmodule


