//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 0 1 0 0 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n792, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT15), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT98), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT97), .B(G36gat), .ZN(new_n206));
  OR3_X1    g005(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n208));
  AOI22_X1  g007(.A1(G29gat), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n205), .B(new_n209), .C1(KEYINPUT15), .C2(new_n203), .ZN(new_n210));
  INV_X1    g009(.A(new_n208), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n211), .B1(new_n207), .B2(KEYINPUT96), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(KEYINPUT96), .B2(new_n207), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n206), .A2(G29gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(KEYINPUT15), .A3(new_n203), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n210), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G15gat), .B(G22gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(G1gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(G1gat), .B2(new_n218), .ZN(new_n221));
  INV_X1    g020(.A(G8gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n221), .B(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n217), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n210), .A2(new_n216), .A3(KEYINPUT17), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(new_n223), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT17), .B1(new_n210), .B2(new_n216), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n202), .B(new_n225), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(KEYINPUT99), .A2(KEYINPUT18), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n228), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(new_n223), .A3(new_n226), .ZN(new_n233));
  INV_X1    g032(.A(new_n230), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n233), .A2(new_n202), .A3(new_n225), .A4(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n217), .B(new_n224), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n202), .B(KEYINPUT13), .Z(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n231), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT95), .ZN(new_n240));
  XNOR2_X1  g039(.A(G113gat), .B(G141gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT94), .B(G197gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT11), .B(G169gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT12), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n239), .A2(new_n240), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n246), .B1(new_n239), .B2(new_n240), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G197gat), .B(G204gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT22), .ZN(new_n252));
  INV_X1    g051(.A(G211gat), .ZN(new_n253));
  INV_X1    g052(.A(G218gat), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G211gat), .B(G218gat), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n251), .A3(new_n255), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G148gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT82), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT82), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G148gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n263), .A2(new_n265), .A3(G141gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT83), .ZN(new_n267));
  INV_X1    g066(.A(G141gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT80), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT80), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(G141gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n271), .A3(G148gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT81), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT82), .B(G148gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT83), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n276), .A3(G141gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT80), .B(G141gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n278), .A2(KEYINPUT81), .A3(G148gat), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n267), .A2(new_n274), .A3(new_n277), .A4(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G155gat), .B(G162gat), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(KEYINPUT84), .A2(G155gat), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n282), .B1(KEYINPUT2), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n280), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT3), .ZN(new_n286));
  XOR2_X1   g085(.A(G141gat), .B(G148gat), .Z(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT79), .B(KEYINPUT2), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n281), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n285), .A2(new_n286), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT85), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n289), .B1(new_n280), .B2(new_n284), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(KEYINPUT85), .A3(new_n286), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT29), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n261), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G228gat), .A2(G233gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT3), .B1(new_n261), .B2(new_n297), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n294), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(KEYINPUT89), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT89), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n294), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n300), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n298), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT88), .ZN(new_n308));
  AND4_X1   g107(.A1(KEYINPUT85), .A2(new_n285), .A3(new_n286), .A4(new_n290), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT85), .B1(new_n294), .B2(new_n286), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n297), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n261), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n302), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n308), .B1(new_n313), .B2(new_n300), .ZN(new_n314));
  OAI211_X1 g113(.A(KEYINPUT88), .B(new_n299), .C1(new_n298), .C2(new_n302), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n307), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G22gat), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT90), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G78gat), .B(G106gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(KEYINPUT31), .B(G50gat), .ZN(new_n320));
  XOR2_X1   g119(.A(new_n319), .B(new_n320), .Z(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n316), .A2(new_n317), .ZN(new_n323));
  AOI211_X1 g122(.A(G22gat), .B(new_n307), .C1(new_n314), .C2(new_n315), .ZN(new_n324));
  OAI22_X1  g123(.A1(new_n318), .A2(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n314), .A2(new_n315), .ZN(new_n326));
  INV_X1    g125(.A(new_n307), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G22gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n316), .A2(new_n317), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n329), .A2(KEYINPUT90), .A3(new_n330), .A4(new_n321), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G169gat), .ZN(new_n333));
  INV_X1    g132(.A(G176gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT23), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT23), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n336), .B1(G169gat), .B2(G176gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n339), .A2(KEYINPUT25), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(KEYINPUT66), .ZN(new_n342));
  NAND3_X1  g141(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT65), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g144(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n345), .B(new_n346), .C1(G183gat), .C2(G190gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n340), .B1(new_n342), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n341), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT67), .ZN(new_n350));
  INV_X1    g149(.A(G183gat), .ZN(new_n351));
  INV_X1    g150(.A(G190gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n354));
  AND4_X1   g153(.A1(new_n349), .A2(new_n343), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT25), .B1(new_n355), .B2(new_n339), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n351), .A2(KEYINPUT27), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT27), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G183gat), .ZN(new_n359));
  AND4_X1   g158(.A1(KEYINPUT28), .A2(new_n357), .A3(new_n359), .A4(new_n352), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n357), .A2(KEYINPUT68), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT27), .B(G183gat), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n352), .B(new_n361), .C1(new_n362), .C2(KEYINPUT68), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT28), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n360), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT69), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT26), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT26), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n368), .A2(new_n333), .A3(new_n334), .A4(KEYINPUT69), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n367), .A2(new_n338), .A3(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n370), .B1(new_n351), .B2(new_n352), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n348), .B(new_n356), .C1(new_n365), .C2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G127gat), .B(G134gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT70), .ZN(new_n374));
  INV_X1    g173(.A(G113gat), .ZN(new_n375));
  INV_X1    g174(.A(G120gat), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT1), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n377), .B1(new_n375), .B2(new_n376), .ZN(new_n378));
  INV_X1    g177(.A(G134gat), .ZN(new_n379));
  OR3_X1    g178(.A1(new_n379), .A2(KEYINPUT70), .A3(G127gat), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n374), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  XOR2_X1   g180(.A(KEYINPUT71), .B(G120gat), .Z(new_n382));
  OAI211_X1 g181(.A(new_n377), .B(new_n373), .C1(new_n382), .C2(new_n375), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n372), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G227gat), .A2(G233gat), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n387), .B(KEYINPUT64), .Z(new_n388));
  AOI22_X1  g187(.A1(new_n366), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n389), .A2(new_n369), .B1(G183gat), .B2(G190gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n357), .A2(new_n359), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT68), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(G190gat), .B1(new_n357), .B2(KEYINPUT68), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT28), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n390), .B1(new_n395), .B2(new_n360), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n396), .A2(new_n384), .A3(new_n348), .A4(new_n356), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n386), .A2(new_n388), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT72), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n386), .A2(KEYINPUT72), .A3(new_n388), .A4(new_n397), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  XOR2_X1   g201(.A(G15gat), .B(G43gat), .Z(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(KEYINPUT75), .ZN(new_n404));
  XNOR2_X1  g203(.A(G71gat), .B(G99gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT33), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n402), .A2(KEYINPUT32), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n402), .A2(KEYINPUT32), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT74), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT74), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n402), .A2(new_n411), .A3(KEYINPUT32), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n406), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT33), .B1(new_n400), .B2(new_n401), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(KEYINPUT73), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n408), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n388), .ZN(new_n417));
  INV_X1    g216(.A(new_n386), .ZN(new_n418));
  INV_X1    g217(.A(new_n397), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n420), .B(KEYINPUT34), .Z(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n416), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n421), .B(new_n408), .C1(new_n413), .C2(new_n415), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n332), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT35), .ZN(new_n427));
  INV_X1    g226(.A(new_n294), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n385), .B1(new_n428), .B2(KEYINPUT3), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n296), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n294), .A2(new_n385), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(KEYINPUT4), .ZN(new_n432));
  NAND2_X1  g231(.A1(G225gat), .A2(G233gat), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n294), .B(new_n385), .ZN(new_n435));
  INV_X1    g234(.A(new_n433), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT5), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n430), .A2(new_n432), .A3(KEYINPUT5), .A4(new_n433), .ZN(new_n440));
  XNOR2_X1  g239(.A(G57gat), .B(G85gat), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT87), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  XOR2_X1   g242(.A(G1gat), .B(G29gat), .Z(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT92), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n439), .A2(new_n440), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n447), .B1(new_n439), .B2(new_n440), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n450), .A2(new_n451), .A3(KEYINPUT6), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n439), .A2(new_n447), .A3(new_n440), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n453), .A2(KEYINPUT6), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n427), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G8gat), .B(G36gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(G64gat), .B(G92gat), .ZN(new_n457));
  XOR2_X1   g256(.A(new_n456), .B(new_n457), .Z(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n372), .A2(G226gat), .A3(G233gat), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n372), .A2(KEYINPUT76), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT76), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n396), .A2(new_n462), .A3(new_n348), .A4(new_n356), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n461), .A2(new_n297), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(G226gat), .A2(G233gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n460), .B1(new_n466), .B2(KEYINPUT77), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT77), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n464), .A2(new_n468), .A3(new_n465), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n261), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n461), .A2(new_n463), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(G226gat), .A3(G233gat), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n372), .A2(new_n297), .A3(new_n465), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n312), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n459), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n474), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n464), .A2(new_n468), .A3(new_n465), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n468), .B1(new_n464), .B2(new_n465), .ZN(new_n478));
  NOR3_X1   g277(.A1(new_n477), .A2(new_n478), .A3(new_n460), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n476), .B(new_n458), .C1(new_n479), .C2(new_n261), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT30), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n481), .A2(KEYINPUT78), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n475), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n470), .A2(new_n474), .ZN(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT78), .B(KEYINPUT30), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n458), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT91), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n483), .A2(KEYINPUT91), .A3(new_n486), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n455), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n426), .A2(new_n491), .A3(KEYINPUT93), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT93), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n439), .A2(new_n440), .ZN(new_n494));
  INV_X1    g293(.A(new_n447), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT6), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n439), .A2(new_n440), .A3(new_n449), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n453), .A2(KEYINPUT6), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT35), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n483), .A2(KEYINPUT91), .A3(new_n486), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT91), .B1(new_n483), .B2(new_n486), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n325), .A2(new_n331), .A3(new_n423), .A4(new_n424), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n493), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n496), .B1(new_n495), .B2(new_n494), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n499), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n487), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT35), .B1(new_n504), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n332), .A2(new_n508), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT36), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n425), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n423), .A2(KEYINPUT36), .A3(new_n424), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n430), .A2(new_n432), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n436), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n517), .A2(KEYINPUT39), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT39), .B1(new_n435), .B2(new_n436), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n519), .B1(new_n516), .B2(new_n436), .ZN(new_n520));
  NOR3_X1   g319(.A1(new_n518), .A2(new_n520), .A3(new_n449), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n521), .A2(KEYINPUT40), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n450), .B1(new_n521), .B2(KEYINPUT40), .ZN(new_n523));
  AND4_X1   g322(.A1(new_n489), .A2(new_n490), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT37), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n458), .B1(new_n484), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n467), .A2(new_n469), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n261), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n472), .A2(new_n473), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n525), .B1(new_n529), .B2(new_n312), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT38), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n496), .A2(new_n497), .B1(KEYINPUT6), .B2(new_n453), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(new_n533), .A3(new_n480), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT38), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT37), .B1(new_n470), .B2(new_n474), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(new_n526), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n331), .B(new_n325), .C1(new_n534), .C2(new_n537), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n511), .B(new_n515), .C1(new_n524), .C2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n250), .B1(new_n510), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G71gat), .B(G78gat), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n541), .A2(KEYINPUT100), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(KEYINPUT100), .ZN(new_n543));
  XNOR2_X1  g342(.A(G57gat), .B(G64gat), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n542), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  OAI211_X1 g346(.A(KEYINPUT100), .B(new_n541), .C1(new_n544), .C2(new_n545), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n549), .A2(KEYINPUT21), .ZN(new_n550));
  NAND2_X1  g349(.A1(G231gat), .A2(G233gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G127gat), .B(G155gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT20), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n552), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G183gat), .B(G211gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT102), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n555), .B(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n224), .B1(KEYINPUT21), .B2(new_n549), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT101), .B(KEYINPUT19), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n559), .B(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G85gat), .A2(G92gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT7), .ZN(new_n565));
  NAND2_X1  g364(.A1(G99gat), .A2(G106gat), .ZN(new_n566));
  INV_X1    g365(.A(G85gat), .ZN(new_n567));
  INV_X1    g366(.A(G92gat), .ZN(new_n568));
  AOI22_X1  g367(.A1(KEYINPUT8), .A2(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G99gat), .B(G106gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n572), .A2(KEYINPUT10), .A3(new_n549), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT104), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n570), .B(new_n571), .Z(new_n575));
  NAND3_X1  g374(.A1(new_n565), .A2(new_n571), .A3(new_n569), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT103), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(new_n577), .A3(new_n549), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n549), .A2(new_n577), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n572), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT10), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n574), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AOI211_X1 g382(.A(KEYINPUT104), .B(KEYINPUT10), .C1(new_n578), .C2(new_n580), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n573), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G230gat), .A2(G233gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n586), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n578), .A2(new_n588), .A3(new_n580), .ZN(new_n589));
  XNOR2_X1  g388(.A(G120gat), .B(G148gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(G176gat), .B(G204gat), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n590), .B(new_n591), .Z(new_n592));
  NAND3_X1  g391(.A1(new_n587), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n592), .B1(new_n587), .B2(new_n589), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  AND2_X1   g396(.A1(G232gat), .A2(G233gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n217), .A2(new_n572), .B1(KEYINPUT41), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n226), .A2(new_n575), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n599), .B1(new_n600), .B2(new_n228), .ZN(new_n601));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n598), .A2(KEYINPUT41), .ZN(new_n604));
  XNOR2_X1  g403(.A(G134gat), .B(G162gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  OR2_X1    g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n563), .A2(new_n597), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n540), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n507), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g415(.A1(new_n501), .A2(new_n502), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT105), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT42), .ZN(new_n620));
  XOR2_X1   g419(.A(KEYINPUT16), .B(G8gat), .Z(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NOR4_X1   g421(.A1(new_n618), .A2(new_n619), .A3(new_n620), .A4(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n618), .A2(new_n622), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT105), .B1(new_n624), .B2(KEYINPUT42), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n222), .B1(new_n613), .B2(new_n617), .ZN(new_n626));
  OAI22_X1  g425(.A1(new_n626), .A2(new_n620), .B1(new_n618), .B2(new_n622), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n623), .B1(new_n625), .B2(new_n627), .ZN(G1325gat));
  OAI21_X1  g427(.A(G15gat), .B1(new_n612), .B2(new_n515), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n425), .A2(G15gat), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n629), .B1(new_n612), .B2(new_n630), .ZN(G1326gat));
  INV_X1    g430(.A(new_n332), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n612), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(KEYINPUT43), .B(G22gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(G1327gat));
  INV_X1    g434(.A(G29gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n563), .A2(new_n596), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n637), .A2(new_n609), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n540), .A2(new_n636), .A3(new_n614), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT45), .ZN(new_n640));
  AND2_X1   g439(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n641));
  NOR2_X1   g440(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n510), .A2(new_n539), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n643), .B1(new_n644), .B2(new_n610), .ZN(new_n645));
  AOI211_X1 g444(.A(new_n609), .B(new_n641), .C1(new_n510), .C2(new_n539), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n637), .A2(new_n250), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n614), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n640), .B1(new_n650), .B2(new_n636), .ZN(G1328gat));
  NOR3_X1   g450(.A1(new_n637), .A2(new_n206), .A3(new_n609), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n540), .A2(new_n617), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT46), .Z(new_n654));
  OAI211_X1 g453(.A(new_n617), .B(new_n648), .C1(new_n645), .C2(new_n646), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n655), .A2(KEYINPUT107), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n206), .B1(new_n655), .B2(KEYINPUT107), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(G1329gat));
  INV_X1    g457(.A(new_n515), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n659), .B(new_n648), .C1(new_n645), .C2(new_n646), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(G43gat), .ZN(new_n661));
  INV_X1    g460(.A(G43gat), .ZN(new_n662));
  INV_X1    g461(.A(new_n425), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n540), .A2(new_n662), .A3(new_n663), .A4(new_n638), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT47), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n661), .A2(KEYINPUT47), .A3(new_n664), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(G1330gat));
  INV_X1    g468(.A(G50gat), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n632), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n647), .A2(new_n648), .A3(new_n671), .ZN(new_n672));
  OR2_X1    g471(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n540), .A2(new_n332), .A3(new_n638), .ZN(new_n674));
  AOI22_X1  g473(.A1(new_n674), .A2(new_n670), .B1(KEYINPUT108), .B2(KEYINPUT48), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n672), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n673), .B1(new_n672), .B2(new_n675), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(G1331gat));
  NOR3_X1   g477(.A1(new_n563), .A2(new_n610), .A3(new_n249), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n597), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT109), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n644), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n614), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g483(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n617), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT110), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n688), .A2(KEYINPUT111), .ZN(new_n689));
  NOR2_X1   g488(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(KEYINPUT111), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n690), .B1(new_n689), .B2(new_n691), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(G1333gat));
  NAND3_X1  g493(.A1(new_n682), .A2(G71gat), .A3(new_n659), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n425), .B(KEYINPUT112), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n682), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n695), .B1(new_n698), .B2(G71gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g499(.A1(new_n682), .A2(new_n332), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G78gat), .ZN(G1335gat));
  INV_X1    g501(.A(new_n563), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT113), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n703), .A2(new_n704), .A3(new_n249), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT113), .B1(new_n563), .B2(new_n250), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n596), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n647), .A2(new_n614), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G85gat), .ZN(new_n710));
  INV_X1    g509(.A(new_n707), .ZN(new_n711));
  AND2_X1   g510(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n712));
  NOR2_X1   g511(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n644), .A2(new_n610), .A3(new_n711), .A4(new_n715), .ZN(new_n716));
  AOI211_X1 g515(.A(new_n609), .B(new_n707), .C1(new_n510), .C2(new_n539), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n717), .B2(new_n712), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n614), .A2(new_n567), .A3(new_n597), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n710), .B1(new_n719), .B2(new_n720), .ZN(G1336gat));
  OAI211_X1 g520(.A(new_n617), .B(new_n708), .C1(new_n645), .C2(new_n646), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(G92gat), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n718), .A2(new_n568), .A3(new_n617), .A4(new_n597), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT52), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT52), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n723), .A2(new_n724), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(G1337gat));
  INV_X1    g528(.A(G99gat), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n659), .B(new_n708), .C1(new_n645), .C2(new_n646), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n730), .B1(new_n731), .B2(KEYINPUT115), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(KEYINPUT115), .B2(new_n731), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n663), .A2(new_n730), .A3(new_n597), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT116), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n719), .B2(new_n735), .ZN(G1338gat));
  INV_X1    g535(.A(G106gat), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n632), .A2(new_n737), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n708), .B(new_n738), .C1(new_n645), .C2(new_n646), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT53), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT117), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n632), .A2(new_n596), .ZN(new_n743));
  INV_X1    g542(.A(new_n716), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n609), .B1(new_n510), .B2(new_n539), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n712), .B1(new_n745), .B2(new_n711), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n743), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n737), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n740), .A2(KEYINPUT117), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n742), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n739), .A2(new_n741), .ZN(new_n752));
  AOI21_X1  g551(.A(G106gat), .B1(new_n718), .B2(new_n743), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n749), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n751), .A2(new_n754), .ZN(G1339gat));
  NAND2_X1  g554(.A1(new_n679), .A2(new_n596), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n588), .B(new_n573), .C1(new_n583), .C2(new_n584), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n587), .A2(KEYINPUT54), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT54), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n585), .A2(new_n761), .A3(new_n586), .ZN(new_n762));
  INV_X1    g561(.A(new_n592), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n757), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n764), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n766), .A2(new_n759), .A3(KEYINPUT55), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n765), .A2(new_n593), .A3(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n231), .A2(new_n235), .A3(new_n238), .A4(new_n246), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n202), .B1(new_n233), .B2(new_n225), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n236), .A2(new_n237), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n245), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n607), .A2(new_n773), .A3(new_n608), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n768), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n765), .A2(new_n249), .A3(new_n767), .A4(new_n593), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n773), .B1(new_n594), .B2(new_n595), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT118), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n773), .B(new_n779), .C1(new_n594), .C2(new_n595), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n776), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n775), .B1(new_n781), .B2(new_n609), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n756), .B1(new_n782), .B2(new_n703), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(new_n504), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n617), .A2(new_n507), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n250), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(new_n375), .ZN(G1340gat));
  NOR2_X1   g588(.A1(new_n787), .A2(new_n596), .ZN(new_n790));
  MUX2_X1   g589(.A(G120gat), .B(new_n382), .S(new_n790), .Z(G1341gat));
  NOR2_X1   g590(.A1(new_n787), .A2(new_n563), .ZN(new_n792));
  XOR2_X1   g591(.A(KEYINPUT119), .B(G127gat), .Z(new_n793));
  XNOR2_X1  g592(.A(new_n792), .B(new_n793), .ZN(G1342gat));
  OAI21_X1  g593(.A(G134gat), .B1(new_n787), .B2(new_n609), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n617), .A2(new_n609), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n796), .A2(new_n379), .A3(new_n614), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT56), .B1(new_n785), .B2(new_n798), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n785), .A2(KEYINPUT56), .A3(new_n798), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n795), .B1(new_n799), .B2(new_n800), .ZN(G1343gat));
  NAND2_X1  g600(.A1(new_n783), .A2(new_n332), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n515), .ZN(new_n803));
  NOR4_X1   g602(.A1(new_n802), .A2(G141gat), .A3(new_n250), .A4(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n803), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n332), .A2(KEYINPUT57), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n610), .B1(new_n776), .B2(new_n777), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n563), .B1(new_n807), .B2(new_n775), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT120), .ZN(new_n809));
  AOI22_X1  g608(.A1(new_n808), .A2(new_n809), .B1(new_n596), .B2(new_n679), .ZN(new_n810));
  OAI211_X1 g609(.A(KEYINPUT120), .B(new_n563), .C1(new_n807), .C2(new_n775), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n806), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT57), .B1(new_n783), .B2(new_n332), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n249), .B(new_n805), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n278), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n804), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT121), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n816), .A2(new_n817), .A3(KEYINPUT58), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(KEYINPUT58), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n817), .A2(KEYINPUT58), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n816), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n818), .A2(new_n821), .ZN(G1344gat));
  INV_X1    g621(.A(new_n802), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n823), .A2(new_n275), .A3(new_n597), .A4(new_n805), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n810), .A2(new_n811), .ZN(new_n825));
  INV_X1    g624(.A(new_n806), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n813), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n803), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI211_X1 g628(.A(KEYINPUT59), .B(new_n275), .C1(new_n829), .C2(new_n597), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n632), .B1(new_n808), .B2(new_n756), .ZN(new_n832));
  OAI22_X1  g631(.A1(new_n784), .A2(new_n806), .B1(new_n832), .B2(KEYINPUT57), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n833), .A2(new_n597), .A3(new_n805), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n831), .B1(new_n834), .B2(G148gat), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n824), .B1(new_n830), .B2(new_n835), .ZN(G1345gat));
  XNOR2_X1  g635(.A(KEYINPUT84), .B(G155gat), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n823), .A2(new_n703), .A3(new_n805), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n838), .A2(KEYINPUT122), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(KEYINPUT122), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n703), .A2(new_n837), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(new_n829), .B2(new_n842), .ZN(G1346gat));
  NAND2_X1  g642(.A1(new_n829), .A2(new_n610), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT123), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n829), .A2(KEYINPUT123), .A3(new_n610), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(G162gat), .A3(new_n847), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n659), .A2(G162gat), .A3(new_n507), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n823), .A2(new_n796), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(G1347gat));
  NAND2_X1  g650(.A1(new_n783), .A2(new_n507), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n617), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n696), .A2(new_n854), .A3(new_n332), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n856), .A2(new_n333), .A3(new_n250), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n854), .A2(new_n504), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT124), .ZN(new_n859));
  OR3_X1    g658(.A1(new_n852), .A2(new_n859), .A3(KEYINPUT125), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT125), .B1(new_n852), .B2(new_n859), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n249), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n857), .B1(new_n862), .B2(new_n333), .ZN(G1348gat));
  NAND4_X1  g662(.A1(new_n860), .A2(new_n334), .A3(new_n597), .A4(new_n861), .ZN(new_n864));
  OAI21_X1  g663(.A(G176gat), .B1(new_n856), .B2(new_n596), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(G1349gat));
  OR4_X1    g665(.A1(new_n391), .A2(new_n852), .A3(new_n859), .A4(new_n563), .ZN(new_n867));
  OAI21_X1  g666(.A(G183gat), .B1(new_n856), .B2(new_n563), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g669(.A1(new_n860), .A2(new_n352), .A3(new_n610), .A4(new_n861), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n853), .A2(new_n610), .A3(new_n855), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT61), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n872), .A2(new_n873), .A3(G190gat), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n872), .B2(G190gat), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(G1351gat));
  NAND3_X1  g675(.A1(new_n515), .A2(new_n507), .A3(new_n617), .ZN(new_n877));
  XOR2_X1   g676(.A(new_n877), .B(KEYINPUT126), .Z(new_n878));
  AND2_X1   g677(.A1(new_n833), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(G197gat), .A3(new_n249), .ZN(new_n880));
  INV_X1    g679(.A(G197gat), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n802), .A2(new_n877), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(new_n250), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n880), .A2(new_n883), .ZN(G1352gat));
  OR3_X1    g683(.A1(new_n882), .A2(G204gat), .A3(new_n596), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n885), .A2(KEYINPUT62), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n879), .A2(new_n597), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(G204gat), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n885), .A2(KEYINPUT62), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(G1353gat));
  NOR2_X1   g689(.A1(new_n877), .A2(new_n563), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n253), .B1(new_n833), .B2(new_n891), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n892), .A2(KEYINPUT63), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(KEYINPUT63), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n703), .A2(new_n253), .ZN(new_n895));
  OAI22_X1  g694(.A1(new_n893), .A2(new_n894), .B1(new_n882), .B2(new_n895), .ZN(G1354gat));
  OAI21_X1  g695(.A(new_n254), .B1(new_n882), .B2(new_n609), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n897), .A2(KEYINPUT127), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(KEYINPUT127), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n609), .A2(new_n254), .ZN(new_n900));
  AOI22_X1  g699(.A1(new_n898), .A2(new_n899), .B1(new_n879), .B2(new_n900), .ZN(G1355gat));
endmodule


