

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U325 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n387) );
  XNOR2_X1 U326 ( .A(n388), .B(n387), .ZN(n427) );
  INV_X1 U327 ( .A(KEYINPUT55), .ZN(n450) );
  XNOR2_X1 U328 ( .A(n450), .B(KEYINPUT119), .ZN(n451) );
  XNOR2_X1 U329 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U330 ( .A(n366), .B(n365), .Z(n572) );
  XNOR2_X1 U331 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U332 ( .A(n457), .B(n456), .ZN(G1349GAT) );
  XNOR2_X1 U333 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n293) );
  XNOR2_X1 U334 ( .A(n293), .B(KEYINPUT86), .ZN(n294) );
  XOR2_X1 U335 ( .A(n294), .B(KEYINPUT19), .Z(n296) );
  XNOR2_X1 U336 ( .A(G169GAT), .B(G183GAT), .ZN(n295) );
  XNOR2_X1 U337 ( .A(n296), .B(n295), .ZN(n446) );
  XOR2_X1 U338 ( .A(G120GAT), .B(G71GAT), .Z(n358) );
  XOR2_X1 U339 ( .A(G15GAT), .B(G127GAT), .Z(n389) );
  XOR2_X1 U340 ( .A(n358), .B(n389), .Z(n298) );
  NAND2_X1 U341 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U343 ( .A(G134GAT), .B(KEYINPUT0), .Z(n341) );
  XOR2_X1 U344 ( .A(n299), .B(n341), .Z(n307) );
  XOR2_X1 U345 ( .A(KEYINPUT20), .B(G99GAT), .Z(n301) );
  XNOR2_X1 U346 ( .A(G43GAT), .B(G190GAT), .ZN(n300) );
  XNOR2_X1 U347 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U348 ( .A(G176GAT), .B(KEYINPUT85), .Z(n303) );
  XNOR2_X1 U349 ( .A(G113GAT), .B(KEYINPUT87), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U351 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U352 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U353 ( .A(n446), .B(n308), .ZN(n532) );
  XNOR2_X1 U354 ( .A(G211GAT), .B(G218GAT), .ZN(n309) );
  XNOR2_X1 U355 ( .A(n309), .B(KEYINPUT88), .ZN(n310) );
  XOR2_X1 U356 ( .A(n310), .B(KEYINPUT21), .Z(n312) );
  XNOR2_X1 U357 ( .A(G197GAT), .B(G204GAT), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n442) );
  XOR2_X1 U359 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n314) );
  XNOR2_X1 U360 ( .A(G141GAT), .B(KEYINPUT89), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n314), .B(n313), .ZN(n339) );
  XOR2_X1 U362 ( .A(G22GAT), .B(G155GAT), .Z(n392) );
  XOR2_X1 U363 ( .A(n339), .B(n392), .Z(n316) );
  NAND2_X1 U364 ( .A1(G228GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U366 ( .A(KEYINPUT90), .B(KEYINPUT23), .Z(n318) );
  XNOR2_X1 U367 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U369 ( .A(n320), .B(n319), .Z(n324) );
  XNOR2_X1 U370 ( .A(G50GAT), .B(KEYINPUT77), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n321), .B(G162GAT), .ZN(n413) );
  XNOR2_X1 U372 ( .A(G106GAT), .B(G78GAT), .ZN(n322) );
  XNOR2_X1 U373 ( .A(n322), .B(G148GAT), .ZN(n349) );
  XNOR2_X1 U374 ( .A(n413), .B(n349), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U376 ( .A(n442), .B(n325), .ZN(n473) );
  XOR2_X1 U377 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n327) );
  XNOR2_X1 U378 ( .A(KEYINPUT93), .B(KEYINPUT1), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n327), .B(n326), .ZN(n345) );
  XOR2_X1 U380 ( .A(G85GAT), .B(G155GAT), .Z(n329) );
  XNOR2_X1 U381 ( .A(G29GAT), .B(G162GAT), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U383 ( .A(KEYINPUT6), .B(G148GAT), .Z(n331) );
  XNOR2_X1 U384 ( .A(G120GAT), .B(G127GAT), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U386 ( .A(n333), .B(n332), .Z(n338) );
  XOR2_X1 U387 ( .A(KEYINPUT5), .B(G57GAT), .Z(n335) );
  NAND2_X1 U388 ( .A1(G225GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U389 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U390 ( .A(KEYINPUT4), .B(n336), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n338), .B(n337), .ZN(n340) );
  XOR2_X1 U392 ( .A(n340), .B(n339), .Z(n343) );
  XOR2_X1 U393 ( .A(G113GAT), .B(G1GAT), .Z(n381) );
  XNOR2_X1 U394 ( .A(n381), .B(n341), .ZN(n342) );
  XNOR2_X1 U395 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U396 ( .A(n345), .B(n344), .Z(n517) );
  XOR2_X1 U397 ( .A(KEYINPUT76), .B(KEYINPUT31), .Z(n347) );
  XNOR2_X1 U398 ( .A(G204GAT), .B(KEYINPUT75), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n347), .B(n346), .ZN(n366) );
  XNOR2_X1 U400 ( .A(G176GAT), .B(G92GAT), .ZN(n348) );
  XNOR2_X1 U401 ( .A(n348), .B(G64GAT), .ZN(n441) );
  XNOR2_X1 U402 ( .A(n349), .B(n441), .ZN(n352) );
  XOR2_X1 U403 ( .A(KEYINPUT13), .B(KEYINPUT72), .Z(n351) );
  XNOR2_X1 U404 ( .A(G57GAT), .B(KEYINPUT73), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n351), .B(n350), .ZN(n393) );
  XNOR2_X1 U406 ( .A(n352), .B(n393), .ZN(n357) );
  XNOR2_X1 U407 ( .A(KEYINPUT33), .B(KEYINPUT74), .ZN(n354) );
  AND2_X1 U408 ( .A1(G230GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U410 ( .A(n355), .B(KEYINPUT32), .Z(n356) );
  XNOR2_X1 U411 ( .A(n357), .B(n356), .ZN(n359) );
  XOR2_X1 U412 ( .A(G99GAT), .B(G85GAT), .Z(n409) );
  XOR2_X1 U413 ( .A(n358), .B(n409), .Z(n360) );
  NAND2_X1 U414 ( .A1(n359), .A2(n360), .ZN(n364) );
  INV_X1 U415 ( .A(n359), .ZN(n362) );
  INV_X1 U416 ( .A(n360), .ZN(n361) );
  NAND2_X1 U417 ( .A1(n362), .A2(n361), .ZN(n363) );
  NAND2_X1 U418 ( .A1(n364), .A2(n363), .ZN(n365) );
  XOR2_X1 U419 ( .A(KEYINPUT41), .B(n572), .Z(n550) );
  XOR2_X1 U420 ( .A(KEYINPUT69), .B(KEYINPUT8), .Z(n368) );
  XNOR2_X1 U421 ( .A(G43GAT), .B(G29GAT), .ZN(n367) );
  XNOR2_X1 U422 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U423 ( .A(KEYINPUT7), .B(n369), .Z(n423) );
  XOR2_X1 U424 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n371) );
  XNOR2_X1 U425 ( .A(KEYINPUT68), .B(KEYINPUT30), .ZN(n370) );
  XNOR2_X1 U426 ( .A(n371), .B(n370), .ZN(n385) );
  XOR2_X1 U427 ( .A(G141GAT), .B(G22GAT), .Z(n373) );
  XNOR2_X1 U428 ( .A(G50GAT), .B(G36GAT), .ZN(n372) );
  XNOR2_X1 U429 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U430 ( .A(G8GAT), .B(G15GAT), .Z(n375) );
  XNOR2_X1 U431 ( .A(G169GAT), .B(G197GAT), .ZN(n374) );
  XNOR2_X1 U432 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U433 ( .A(n377), .B(n376), .Z(n383) );
  XOR2_X1 U434 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n379) );
  NAND2_X1 U435 ( .A1(G229GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U438 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U439 ( .A(n385), .B(n384), .Z(n386) );
  XNOR2_X1 U440 ( .A(n423), .B(n386), .ZN(n502) );
  INV_X1 U441 ( .A(n502), .ZN(n567) );
  NAND2_X1 U442 ( .A1(n550), .A2(n567), .ZN(n388) );
  XOR2_X1 U443 ( .A(G8GAT), .B(KEYINPUT80), .Z(n436) );
  XOR2_X1 U444 ( .A(n436), .B(G78GAT), .Z(n391) );
  XNOR2_X1 U445 ( .A(n389), .B(G211GAT), .ZN(n390) );
  XNOR2_X1 U446 ( .A(n391), .B(n390), .ZN(n397) );
  XOR2_X1 U447 ( .A(n393), .B(n392), .Z(n395) );
  NAND2_X1 U448 ( .A1(G231GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U449 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U450 ( .A(n397), .B(n396), .Z(n399) );
  XNOR2_X1 U451 ( .A(G183GAT), .B(G71GAT), .ZN(n398) );
  XNOR2_X1 U452 ( .A(n399), .B(n398), .ZN(n407) );
  XOR2_X1 U453 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n401) );
  XNOR2_X1 U454 ( .A(G1GAT), .B(G64GAT), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U456 ( .A(KEYINPUT15), .B(KEYINPUT83), .Z(n403) );
  XNOR2_X1 U457 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n402) );
  XNOR2_X1 U458 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U459 ( .A(n405), .B(n404), .Z(n406) );
  XNOR2_X1 U460 ( .A(n407), .B(n406), .ZN(n577) );
  XNOR2_X1 U461 ( .A(G36GAT), .B(G190GAT), .ZN(n408) );
  XNOR2_X1 U462 ( .A(n408), .B(KEYINPUT79), .ZN(n439) );
  XOR2_X1 U463 ( .A(n439), .B(n409), .Z(n411) );
  NAND2_X1 U464 ( .A1(G232GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U465 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U466 ( .A(n412), .B(KEYINPUT9), .Z(n415) );
  XNOR2_X1 U467 ( .A(n413), .B(KEYINPUT11), .ZN(n414) );
  XNOR2_X1 U468 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U469 ( .A(KEYINPUT78), .B(G106GAT), .Z(n417) );
  XNOR2_X1 U470 ( .A(G134GAT), .B(G218GAT), .ZN(n416) );
  XNOR2_X1 U471 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U472 ( .A(n419), .B(n418), .Z(n425) );
  XOR2_X1 U473 ( .A(KEYINPUT64), .B(KEYINPUT10), .Z(n421) );
  XNOR2_X1 U474 ( .A(G92GAT), .B(KEYINPUT66), .ZN(n420) );
  XNOR2_X1 U475 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U476 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U477 ( .A(n425), .B(n424), .ZN(n460) );
  INV_X1 U478 ( .A(n460), .ZN(n561) );
  NOR2_X1 U479 ( .A1(n577), .A2(n561), .ZN(n426) );
  AND2_X1 U480 ( .A1(n427), .A2(n426), .ZN(n428) );
  XNOR2_X1 U481 ( .A(n428), .B(KEYINPUT47), .ZN(n434) );
  XOR2_X1 U482 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n430) );
  XOR2_X1 U483 ( .A(KEYINPUT36), .B(n460), .Z(n579) );
  NAND2_X1 U484 ( .A1(n579), .A2(n577), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n431) );
  NOR2_X1 U486 ( .A1(n572), .A2(n431), .ZN(n432) );
  NAND2_X1 U487 ( .A1(n432), .A2(n502), .ZN(n433) );
  NAND2_X1 U488 ( .A1(n434), .A2(n433), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n435), .B(KEYINPUT48), .ZN(n531) );
  XOR2_X1 U490 ( .A(KEYINPUT94), .B(n436), .Z(n438) );
  NAND2_X1 U491 ( .A1(G226GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n440) );
  XOR2_X1 U493 ( .A(n440), .B(n439), .Z(n444) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U495 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U496 ( .A(n446), .B(n445), .ZN(n466) );
  NAND2_X1 U497 ( .A1(n531), .A2(n466), .ZN(n448) );
  XOR2_X1 U498 ( .A(KEYINPUT54), .B(KEYINPUT118), .Z(n447) );
  XNOR2_X1 U499 ( .A(n448), .B(n447), .ZN(n449) );
  NAND2_X1 U500 ( .A1(n517), .A2(n449), .ZN(n565) );
  NOR2_X1 U501 ( .A1(n473), .A2(n565), .ZN(n452) );
  NOR2_X1 U502 ( .A1(n532), .A2(n453), .ZN(n562) );
  NAND2_X1 U503 ( .A1(n562), .A2(n550), .ZN(n457) );
  XOR2_X1 U504 ( .A(KEYINPUT120), .B(KEYINPUT57), .Z(n455) );
  XNOR2_X1 U505 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n454) );
  XOR2_X1 U506 ( .A(KEYINPUT34), .B(KEYINPUT97), .Z(n459) );
  XNOR2_X1 U507 ( .A(G1GAT), .B(KEYINPUT98), .ZN(n458) );
  XNOR2_X1 U508 ( .A(n459), .B(n458), .ZN(n479) );
  OR2_X1 U509 ( .A1(n502), .A2(n572), .ZN(n492) );
  XOR2_X1 U510 ( .A(KEYINPUT16), .B(KEYINPUT84), .Z(n462) );
  NAND2_X1 U511 ( .A1(n460), .A2(n577), .ZN(n461) );
  XNOR2_X1 U512 ( .A(n462), .B(n461), .ZN(n477) );
  XOR2_X1 U513 ( .A(KEYINPUT95), .B(KEYINPUT26), .Z(n464) );
  NAND2_X1 U514 ( .A1(n473), .A2(n532), .ZN(n463) );
  XNOR2_X1 U515 ( .A(n464), .B(n463), .ZN(n566) );
  XOR2_X1 U516 ( .A(KEYINPUT27), .B(n466), .Z(n472) );
  NOR2_X1 U517 ( .A1(n566), .A2(n472), .ZN(n465) );
  XOR2_X1 U518 ( .A(KEYINPUT96), .B(n465), .Z(n470) );
  INV_X1 U519 ( .A(n466), .ZN(n521) );
  NOR2_X1 U520 ( .A1(n521), .A2(n532), .ZN(n467) );
  NOR2_X1 U521 ( .A1(n473), .A2(n467), .ZN(n468) );
  XNOR2_X1 U522 ( .A(KEYINPUT25), .B(n468), .ZN(n469) );
  NAND2_X1 U523 ( .A1(n470), .A2(n469), .ZN(n471) );
  NAND2_X1 U524 ( .A1(n517), .A2(n471), .ZN(n476) );
  NOR2_X1 U525 ( .A1(n517), .A2(n472), .ZN(n530) );
  XNOR2_X1 U526 ( .A(KEYINPUT28), .B(n473), .ZN(n535) );
  INV_X1 U527 ( .A(n535), .ZN(n526) );
  AND2_X1 U528 ( .A1(n526), .A2(n532), .ZN(n474) );
  NAND2_X1 U529 ( .A1(n530), .A2(n474), .ZN(n475) );
  NAND2_X1 U530 ( .A1(n476), .A2(n475), .ZN(n488) );
  NAND2_X1 U531 ( .A1(n477), .A2(n488), .ZN(n503) );
  OR2_X1 U532 ( .A1(n492), .A2(n503), .ZN(n485) );
  NOR2_X1 U533 ( .A1(n517), .A2(n485), .ZN(n478) );
  XOR2_X1 U534 ( .A(n479), .B(n478), .Z(G1324GAT) );
  NOR2_X1 U535 ( .A1(n521), .A2(n485), .ZN(n480) );
  XOR2_X1 U536 ( .A(G8GAT), .B(n480), .Z(G1325GAT) );
  NOR2_X1 U537 ( .A1(n485), .A2(n532), .ZN(n484) );
  XOR2_X1 U538 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n482) );
  XNOR2_X1 U539 ( .A(G15GAT), .B(KEYINPUT100), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(G1326GAT) );
  NOR2_X1 U542 ( .A1(n526), .A2(n485), .ZN(n486) );
  XOR2_X1 U543 ( .A(G22GAT), .B(n486), .Z(G1327GAT) );
  XNOR2_X1 U544 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n487), .B(KEYINPUT39), .ZN(n495) );
  NAND2_X1 U546 ( .A1(n579), .A2(n488), .ZN(n489) );
  NOR2_X1 U547 ( .A1(n577), .A2(n489), .ZN(n491) );
  XNOR2_X1 U548 ( .A(KEYINPUT37), .B(KEYINPUT102), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n491), .B(n490), .ZN(n516) );
  NOR2_X1 U550 ( .A1(n516), .A2(n492), .ZN(n493) );
  XOR2_X1 U551 ( .A(KEYINPUT38), .B(n493), .Z(n500) );
  NOR2_X1 U552 ( .A1(n517), .A2(n500), .ZN(n494) );
  XOR2_X1 U553 ( .A(n495), .B(n494), .Z(G1328GAT) );
  NOR2_X1 U554 ( .A1(n521), .A2(n500), .ZN(n496) );
  XOR2_X1 U555 ( .A(G36GAT), .B(n496), .Z(G1329GAT) );
  NOR2_X1 U556 ( .A1(n500), .A2(n532), .ZN(n498) );
  XNOR2_X1 U557 ( .A(KEYINPUT40), .B(KEYINPUT103), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n499), .ZN(G1330GAT) );
  NOR2_X1 U560 ( .A1(n500), .A2(n526), .ZN(n501) );
  XOR2_X1 U561 ( .A(G50GAT), .B(n501), .Z(G1331GAT) );
  XNOR2_X1 U562 ( .A(KEYINPUT42), .B(KEYINPUT105), .ZN(n506) );
  NAND2_X1 U563 ( .A1(n550), .A2(n502), .ZN(n515) );
  NOR2_X1 U564 ( .A1(n515), .A2(n503), .ZN(n504) );
  XOR2_X1 U565 ( .A(KEYINPUT104), .B(n504), .Z(n510) );
  NOR2_X1 U566 ( .A1(n517), .A2(n510), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(n507), .ZN(G1332GAT) );
  NOR2_X1 U569 ( .A1(n521), .A2(n510), .ZN(n508) );
  XOR2_X1 U570 ( .A(G64GAT), .B(n508), .Z(G1333GAT) );
  NOR2_X1 U571 ( .A1(n510), .A2(n532), .ZN(n509) );
  XOR2_X1 U572 ( .A(G71GAT), .B(n509), .Z(G1334GAT) );
  NOR2_X1 U573 ( .A1(n526), .A2(n510), .ZN(n514) );
  XOR2_X1 U574 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n512) );
  XNOR2_X1 U575 ( .A(G78GAT), .B(KEYINPUT106), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  OR2_X1 U578 ( .A1(n516), .A2(n515), .ZN(n525) );
  NOR2_X1 U579 ( .A1(n517), .A2(n525), .ZN(n519) );
  XNOR2_X1 U580 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(n520), .ZN(G1336GAT) );
  NOR2_X1 U583 ( .A1(n521), .A2(n525), .ZN(n522) );
  XOR2_X1 U584 ( .A(KEYINPUT110), .B(n522), .Z(n523) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(n523), .ZN(G1337GAT) );
  NOR2_X1 U586 ( .A1(n532), .A2(n525), .ZN(n524) );
  XOR2_X1 U587 ( .A(G99GAT), .B(n524), .Z(G1338GAT) );
  NOR2_X1 U588 ( .A1(n526), .A2(n525), .ZN(n528) );
  XNOR2_X1 U589 ( .A(KEYINPUT111), .B(KEYINPUT44), .ZN(n527) );
  XNOR2_X1 U590 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n537) );
  NAND2_X1 U593 ( .A1(n531), .A2(n530), .ZN(n547) );
  NOR2_X1 U594 ( .A1(n532), .A2(n547), .ZN(n533) );
  XNOR2_X1 U595 ( .A(n533), .B(KEYINPUT113), .ZN(n534) );
  NOR2_X1 U596 ( .A1(n535), .A2(n534), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n543), .A2(n567), .ZN(n536) );
  XNOR2_X1 U598 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U601 ( .A1(n543), .A2(n550), .ZN(n539) );
  XNOR2_X1 U602 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  NAND2_X1 U603 ( .A1(n577), .A2(n543), .ZN(n541) );
  XNOR2_X1 U604 ( .A(n541), .B(KEYINPUT50), .ZN(n542) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U607 ( .A1(n543), .A2(n561), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U609 ( .A(G134GAT), .B(n546), .ZN(G1343GAT) );
  NOR2_X1 U610 ( .A1(n566), .A2(n547), .ZN(n548) );
  XOR2_X1 U611 ( .A(KEYINPUT117), .B(n548), .Z(n555) );
  NAND2_X1 U612 ( .A1(n567), .A2(n555), .ZN(n549) );
  XNOR2_X1 U613 ( .A(G141GAT), .B(n549), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n552) );
  NAND2_X1 U615 ( .A1(n555), .A2(n550), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U618 ( .A1(n577), .A2(n555), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n554), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U620 ( .A1(n561), .A2(n555), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n556), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U622 ( .A1(n562), .A2(n567), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U624 ( .A1(n577), .A2(n562), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U626 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n559), .B(KEYINPUT121), .ZN(n560) );
  XOR2_X1 U628 ( .A(KEYINPUT122), .B(n560), .Z(n564) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1351GAT) );
  XOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT123), .Z(n569) );
  NOR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n580) );
  NAND2_X1 U633 ( .A1(n580), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n571) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n574) );
  NAND2_X1 U638 ( .A1(n580), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n576) );
  XOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT124), .Z(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n580), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n584) );
  XOR2_X1 U645 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n582) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(G1355GAT) );
endmodule

