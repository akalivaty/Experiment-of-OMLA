//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n551,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n608, new_n610, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G221), .A2(G220), .A3(G219), .A4(G218), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n453), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n467), .A2(new_n469), .A3(G137), .A4(new_n465), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n466), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n472), .A2(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n467), .A2(new_n469), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n465), .A2(G112), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(KEYINPUT3), .B(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT69), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n483), .B1(G124), .B2(new_n486), .ZN(new_n487));
  XOR2_X1   g062(.A(new_n487), .B(KEYINPUT70), .Z(G162));
  NAND4_X1  g063(.A1(new_n467), .A2(new_n469), .A3(G138), .A4(new_n465), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT71), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n484), .A2(new_n491), .A3(G138), .A4(new_n465), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n490), .A2(new_n492), .A3(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n489), .A2(KEYINPUT71), .A3(new_n494), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n467), .A2(new_n469), .A3(G126), .A4(G2105), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n493), .A2(new_n495), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  NAND2_X1  g077(.A1(G75), .A2(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G62), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n503), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(KEYINPUT72), .A2(KEYINPUT6), .A3(G651), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n510), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  OR2_X1    g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n514), .A2(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G88), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n509), .A2(new_n517), .A3(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NAND2_X1  g098(.A1(new_n516), .A2(G51), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n518), .A2(new_n519), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n527), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n524), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n520), .A2(G89), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(G168));
  NAND2_X1  g106(.A1(G77), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G64), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n506), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n520), .A2(G90), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n516), .A2(G52), .ZN(new_n537));
  AND3_X1   g112(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(G171));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G56), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n506), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n513), .B1(new_n541), .B2(KEYINPUT73), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n542), .B1(KEYINPUT73), .B2(new_n541), .ZN(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT74), .B(G43), .ZN(new_n544));
  AOI22_X1  g119(.A1(G81), .A2(new_n520), .B1(new_n516), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT75), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n549), .A2(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(new_n516), .A2(G53), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT76), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  XOR2_X1   g133(.A(KEYINPUT76), .B(KEYINPUT9), .Z(new_n559));
  NAND3_X1  g134(.A1(new_n516), .A2(G53), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n506), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G651), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n520), .A2(G91), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n561), .A2(new_n567), .ZN(G299));
  NAND3_X1  g143(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(G301));
  INV_X1    g144(.A(G168), .ZN(G286));
  INV_X1    g145(.A(G74), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n513), .B1(new_n506), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n572), .B1(G49), .B2(new_n516), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n520), .A2(G87), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(G288));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n518), .B2(new_n519), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT77), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n580), .A2(G73), .A3(G543), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n577), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n514), .A2(new_n515), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n584), .A2(G48), .A3(G543), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n584), .A2(G86), .A3(new_n527), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(new_n520), .A2(G85), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n516), .A2(G47), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n527), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n588), .B(new_n589), .C1(new_n513), .C2(new_n590), .ZN(G290));
  INV_X1    g166(.A(G868), .ZN(new_n592));
  NOR2_X1   g167(.A1(G301), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n520), .A2(G92), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n506), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(new_n516), .B2(G54), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT78), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n593), .B1(new_n602), .B2(new_n592), .ZN(G284));
  AOI21_X1  g178(.A(new_n593), .B1(new_n602), .B2(new_n592), .ZN(G321));
  NAND2_X1  g179(.A1(G299), .A2(new_n592), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n592), .B2(G168), .ZN(G297));
  XOR2_X1   g181(.A(G297), .B(KEYINPUT79), .Z(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n602), .B1(new_n608), .B2(G860), .ZN(G148));
  NOR2_X1   g184(.A1(new_n546), .A2(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n602), .A2(new_n608), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT80), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n610), .B1(new_n612), .B2(G868), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n484), .A2(new_n465), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n615), .A2(new_n466), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XOR2_X1   g192(.A(KEYINPUT81), .B(KEYINPUT13), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT82), .B(G2100), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT83), .ZN(new_n621));
  AND2_X1   g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n479), .A2(G135), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT84), .Z(new_n625));
  NAND2_X1  g200(.A1(new_n486), .A2(G123), .ZN(new_n626));
  OR2_X1    g201(.A1(G99), .A2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n627), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G2096), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(G2096), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n620), .A2(new_n621), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n619), .B1(new_n622), .B2(new_n632), .ZN(new_n633));
  NAND4_X1  g208(.A1(new_n623), .A2(new_n630), .A3(new_n631), .A4(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2427), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT86), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(KEYINPUT14), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT87), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n636), .B2(new_n638), .ZN(new_n642));
  XOR2_X1   g217(.A(G2443), .B(G2446), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT88), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(G14), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n648), .A2(new_n650), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g232(.A1(new_n657), .A2(KEYINPUT17), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n655), .A2(new_n656), .ZN(new_n659));
  AOI21_X1  g234(.A(KEYINPUT18), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n657), .B2(KEYINPUT18), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n660), .B(new_n662), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2100), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT89), .B(G2096), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(G227));
  XOR2_X1   g241(.A(G1971), .B(G1976), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  AND2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT20), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n668), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n668), .B2(new_n674), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G229));
  NOR2_X1   g259(.A1(G29), .A2(G35), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(G162), .B2(G29), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT29), .ZN(new_n687));
  INV_X1    g262(.A(G2090), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT31), .B(G11), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT30), .B(G28), .Z(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(G29), .ZN(new_n692));
  INV_X1    g267(.A(G29), .ZN(new_n693));
  INV_X1    g268(.A(G34), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n694), .A2(KEYINPUT24), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(KEYINPUT24), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n693), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G160), .B2(new_n693), .ZN(new_n698));
  OAI22_X1  g273(.A1(new_n629), .A2(new_n693), .B1(G2084), .B2(new_n698), .ZN(new_n699));
  AOI211_X1 g274(.A(new_n692), .B(new_n699), .C1(G2084), .C2(new_n698), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G5), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G171), .B2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(G1961), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n701), .A2(G21), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G168), .B2(new_n701), .ZN(new_n707));
  INV_X1    g282(.A(G1966), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n693), .A2(G26), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT28), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n486), .A2(G128), .ZN(new_n712));
  NOR2_X1   g287(.A1(G104), .A2(G2105), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT94), .ZN(new_n714));
  INV_X1    g289(.A(G116), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n466), .B1(new_n715), .B2(G2105), .ZN(new_n716));
  AOI22_X1  g291(.A1(G140), .A2(new_n479), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n711), .B1(new_n718), .B2(G29), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT95), .B(G2067), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n700), .A2(new_n705), .A3(new_n709), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n693), .A2(G33), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT25), .Z(new_n725));
  INV_X1    g300(.A(G139), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(new_n615), .ZN(new_n727));
  NAND2_X1  g302(.A1(G115), .A2(G2104), .ZN(new_n728));
  INV_X1    g303(.A(G127), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n478), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n727), .B1(G2105), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT96), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n723), .B1(new_n732), .B2(new_n693), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G2072), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n701), .A2(G20), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT23), .Z(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G299), .B2(G16), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1956), .ZN(new_n738));
  NAND2_X1  g313(.A1(G164), .A2(G29), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G27), .B2(G29), .ZN(new_n740));
  INV_X1    g315(.A(G2078), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n738), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G19), .ZN(new_n745));
  OR3_X1    g320(.A1(new_n745), .A2(KEYINPUT92), .A3(G16), .ZN(new_n746));
  OAI21_X1  g321(.A(KEYINPUT92), .B1(new_n745), .B2(G16), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n746), .B(new_n747), .C1(new_n547), .C2(new_n701), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT93), .B(G1341), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NOR4_X1   g325(.A1(new_n722), .A2(new_n734), .A3(new_n744), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n693), .A2(G32), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n479), .A2(G141), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT97), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n486), .A2(G129), .ZN(new_n755));
  NAND3_X1  g330(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT26), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n758), .A2(new_n759), .B1(G105), .B2(new_n474), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n754), .A2(new_n755), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT98), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n752), .B1(new_n765), .B2(new_n693), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT27), .B(G1996), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT99), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n766), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n701), .A2(G4), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n602), .B2(new_n701), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1348), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n689), .A2(new_n751), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n693), .A2(G25), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n486), .A2(G119), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n465), .A2(G107), .ZN(new_n777));
  OAI21_X1  g352(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n479), .A2(G131), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n775), .B1(new_n782), .B2(new_n693), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT35), .B(G1991), .Z(new_n784));
  XOR2_X1   g359(.A(new_n783), .B(new_n784), .Z(new_n785));
  MUX2_X1   g360(.A(G24), .B(G290), .S(G16), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1986), .ZN(new_n787));
  MUX2_X1   g362(.A(G23), .B(G288), .S(G16), .Z(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT33), .B(G1976), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(G16), .A2(G22), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G166), .B2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT90), .B(G1971), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  MUX2_X1   g369(.A(G6), .B(G305), .S(G16), .Z(new_n795));
  XOR2_X1   g370(.A(KEYINPUT32), .B(G1981), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n790), .A2(new_n794), .A3(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT91), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT34), .ZN(new_n800));
  AOI211_X1 g375(.A(new_n785), .B(new_n787), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(KEYINPUT36), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(KEYINPUT36), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n774), .B1(new_n804), .B2(new_n805), .ZN(G311));
  INV_X1    g381(.A(G311), .ZN(G150));
  NAND2_X1  g382(.A1(new_n602), .A2(G559), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT38), .ZN(new_n809));
  NAND2_X1  g384(.A1(G80), .A2(G543), .ZN(new_n810));
  INV_X1    g385(.A(G67), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n506), .B2(new_n811), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n812), .A2(G651), .B1(new_n516), .B2(G55), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n520), .A2(G93), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n546), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n815), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n817), .A2(new_n543), .A3(new_n545), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n809), .B(new_n819), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n820), .A2(KEYINPUT39), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n820), .A2(KEYINPUT39), .ZN(new_n822));
  NOR3_X1   g397(.A1(new_n821), .A2(new_n822), .A3(G860), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n815), .A2(G860), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT37), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n823), .A2(new_n825), .ZN(G145));
  NAND2_X1  g401(.A1(new_n486), .A2(G130), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n465), .A2(G118), .ZN(new_n828));
  OAI21_X1  g403(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n479), .A2(G142), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n617), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n781), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n732), .B(G164), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n834), .B(new_n835), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n763), .A2(new_n764), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(new_n718), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n718), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n841), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n838), .A2(new_n839), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n836), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(G162), .B(G160), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(new_n629), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n834), .B(new_n835), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n849), .A2(new_n844), .A3(new_n842), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n846), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(G37), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n846), .A2(new_n850), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n853), .B(KEYINPUT40), .C1(new_n848), .C2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT40), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n854), .A2(new_n848), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n851), .A2(new_n852), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n855), .A2(new_n859), .ZN(G395));
  XNOR2_X1  g435(.A(new_n819), .B(KEYINPUT102), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n612), .B(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n565), .A2(new_n566), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(new_n560), .B2(new_n558), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n601), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(G299), .A2(new_n596), .A3(new_n600), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(G288), .A2(G290), .ZN(new_n869));
  NAND2_X1  g444(.A1(G288), .A2(G290), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT103), .ZN(new_n872));
  XNOR2_X1  g447(.A(G303), .B(G305), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n869), .A2(new_n875), .A3(new_n870), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n872), .A2(new_n876), .A3(new_n873), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(KEYINPUT42), .Z(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n865), .A2(new_n866), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT41), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n862), .A2(new_n883), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n868), .A2(new_n880), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n880), .B1(new_n868), .B2(new_n884), .ZN(new_n886));
  OAI21_X1  g461(.A(G868), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n887), .B1(G868), .B2(new_n817), .ZN(G295));
  OAI21_X1  g463(.A(new_n887), .B1(G868), .B2(new_n817), .ZN(G331));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT43), .ZN(new_n891));
  NAND2_X1  g466(.A1(G301), .A2(KEYINPUT104), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(G301), .A2(KEYINPUT104), .ZN(new_n894));
  OAI21_X1  g469(.A(G286), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n894), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(G168), .A3(new_n892), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n867), .B1(new_n898), .B2(new_n819), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n895), .A2(new_n897), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n816), .A2(new_n818), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n900), .A2(KEYINPUT105), .A3(new_n901), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n899), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n819), .A2(new_n897), .A3(new_n895), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n902), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n883), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n878), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT106), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n913), .A3(new_n852), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n906), .A2(new_n909), .A3(new_n878), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n878), .B1(new_n906), .B2(new_n909), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT106), .B1(new_n917), .B2(G37), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n891), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n915), .A2(new_n852), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n904), .A2(new_n907), .A3(new_n905), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n883), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(KEYINPUT107), .A3(new_n883), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n899), .A2(new_n902), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n920), .B1(new_n927), .B2(new_n911), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n928), .A2(new_n891), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n890), .B1(new_n919), .B2(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n914), .A2(new_n918), .A3(new_n891), .A4(new_n915), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n931), .B(KEYINPUT44), .C1(new_n928), .C2(new_n891), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n932), .A2(KEYINPUT108), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(KEYINPUT108), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(G397));
  INV_X1    g510(.A(G1384), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n490), .A2(new_n492), .A3(KEYINPUT4), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n495), .A2(new_n498), .A3(new_n497), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT45), .B1(new_n939), .B2(KEYINPUT109), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n489), .A2(KEYINPUT71), .A3(new_n494), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n941), .A2(new_n499), .ZN(new_n942));
  AOI21_X1  g517(.A(G1384), .B1(new_n942), .B2(new_n493), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n940), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G40), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n472), .A2(new_n476), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g525(.A(new_n718), .B(G2067), .Z(new_n951));
  XNOR2_X1  g526(.A(new_n781), .B(new_n784), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n765), .A2(G1996), .ZN(new_n953));
  INV_X1    g528(.A(G1996), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n837), .A2(new_n954), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n951), .B(new_n952), .C1(new_n953), .C2(new_n955), .ZN(new_n956));
  XOR2_X1   g531(.A(G290), .B(G1986), .Z(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n950), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n961), .B(new_n936), .C1(new_n937), .C2(new_n938), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n501), .A2(KEYINPUT111), .A3(new_n961), .A4(new_n936), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G2084), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n949), .B1(new_n939), .B2(KEYINPUT50), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n939), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n936), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n948), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n708), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n969), .A2(G168), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(G8), .ZN(new_n976));
  AOI21_X1  g551(.A(G168), .B1(new_n969), .B2(new_n974), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT51), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n975), .A2(new_n979), .A3(G8), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT62), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT62), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n978), .A2(new_n983), .A3(new_n980), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n501), .A2(new_n936), .A3(new_n948), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n573), .A2(G1976), .A3(new_n574), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n985), .A2(G8), .A3(new_n986), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n987), .A2(KEYINPUT112), .A3(KEYINPUT52), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT112), .B1(new_n987), .B2(KEYINPUT52), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G8), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(new_n943), .B2(new_n948), .ZN(new_n992));
  INV_X1    g567(.A(G1976), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT52), .B1(G288), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n992), .A2(new_n986), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(G305), .A2(G1981), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n997));
  INV_X1    g572(.A(G1981), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n583), .A2(new_n585), .A3(new_n586), .A4(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n996), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT49), .ZN(new_n1001));
  NAND3_X1  g576(.A1(G305), .A2(KEYINPUT113), .A3(G1981), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n992), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1001), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n995), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n990), .A2(new_n1006), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n968), .A2(new_n688), .A3(new_n962), .ZN(new_n1008));
  XNOR2_X1  g583(.A(KEYINPUT110), .B(G1971), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n949), .B1(new_n939), .B2(new_n970), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1009), .B1(new_n1010), .B2(new_n972), .ZN(new_n1011));
  OAI21_X1  g586(.A(G8), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n1013));
  NOR3_X1   g588(.A1(G166), .A2(new_n1013), .A3(new_n991), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n966), .A2(new_n688), .A3(new_n968), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1009), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n973), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1016), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(G8), .A3(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1007), .A2(new_n1017), .A3(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n971), .A2(new_n741), .A3(new_n948), .A4(new_n972), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1010), .A2(KEYINPUT53), .A3(new_n741), .A4(new_n972), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n948), .B1(new_n943), .B2(new_n961), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1029), .B1(new_n964), .B2(new_n965), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1027), .B(new_n1028), .C1(new_n1030), .C2(G1961), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G171), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1024), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n982), .A2(new_n984), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT49), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1036), .A2(new_n992), .A3(new_n1003), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1037), .B(new_n995), .C1(new_n989), .C2(new_n988), .ZN(new_n1038));
  XOR2_X1   g613(.A(new_n999), .B(KEYINPUT114), .Z(new_n1039));
  NOR2_X1   g614(.A1(G288), .A2(G1976), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n1040), .B(KEYINPUT115), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1039), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n992), .ZN(new_n1043));
  OAI22_X1  g618(.A1(new_n1023), .A2(new_n1038), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT63), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G168), .A2(G8), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1046), .B1(new_n969), .B2(new_n974), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1047), .A2(KEYINPUT116), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n1049));
  AOI211_X1 g624(.A(new_n1049), .B(new_n1046), .C1(new_n969), .C2(new_n974), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1045), .B1(new_n1051), .B2(new_n1024), .ZN(new_n1052));
  AOI211_X1 g627(.A(new_n991), .B(new_n1016), .C1(new_n1018), .C2(new_n1020), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(new_n1038), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1021), .A2(G8), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1045), .B1(new_n1055), .B2(new_n1016), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1054), .B(new_n1056), .C1(new_n1050), .C2(new_n1048), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1044), .B1(new_n1052), .B2(new_n1057), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1034), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT123), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT111), .B1(new_n943), .B2(new_n961), .ZN(new_n1061));
  INV_X1    g636(.A(new_n965), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n968), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n704), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n948), .A2(KEYINPUT53), .A3(new_n741), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(new_n943), .B2(KEYINPUT45), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n946), .A2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1064), .A2(G301), .A3(new_n1027), .A4(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1032), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1060), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT54), .B1(new_n1031), .B2(G171), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1027), .B(new_n1067), .C1(new_n1030), .C2(G1961), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G171), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT124), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT124), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(new_n1076), .A3(G171), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1072), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g653(.A(KEYINPUT123), .B(KEYINPUT54), .C1(new_n1032), .C2(new_n1068), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n1071), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT118), .B1(new_n558), .B2(new_n560), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n558), .A2(KEYINPUT118), .A3(new_n560), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(new_n567), .A3(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1084), .A2(new_n1085), .B1(KEYINPUT57), .B2(new_n864), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT56), .B(G2072), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1010), .A2(new_n972), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(G1956), .B1(new_n968), .B2(new_n962), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1086), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n985), .A2(G2067), .ZN(new_n1091));
  INV_X1    g666(.A(G1348), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n1063), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1090), .B1(new_n1093), .B2(new_n601), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n864), .A2(KEYINPUT57), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1083), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1097), .A2(new_n1081), .A3(new_n863), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1085), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1096), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1956), .ZN(new_n1101));
  INV_X1    g676(.A(new_n962), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1101), .B1(new_n1029), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1010), .A2(new_n972), .A3(new_n1087), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1100), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1094), .A2(new_n1095), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1095), .B1(new_n1094), .B2(new_n1105), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n601), .B1(new_n1093), .B2(KEYINPUT60), .ZN(new_n1109));
  AOI21_X1  g684(.A(G1348), .B1(new_n966), .B2(new_n968), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT60), .ZN(new_n1111));
  INV_X1    g686(.A(new_n601), .ZN(new_n1112));
  NOR4_X1   g687(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .A4(new_n1091), .ZN(new_n1113));
  OAI22_X1  g688(.A1(new_n1109), .A2(new_n1113), .B1(KEYINPUT60), .B2(new_n1093), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n547), .A2(KEYINPUT121), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1010), .A2(new_n954), .A3(new_n972), .ZN(new_n1116));
  XOR2_X1   g691(.A(KEYINPUT58), .B(G1341), .Z(new_n1117));
  NAND2_X1  g692(.A1(new_n985), .A2(new_n1117), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1116), .A2(KEYINPUT120), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT120), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1115), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g698(.A(KEYINPUT59), .B(new_n1115), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1114), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1090), .A2(new_n1105), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT61), .B1(new_n1126), .B2(KEYINPUT122), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n1129));
  AOI211_X1 g704(.A(new_n1128), .B(new_n1129), .C1(new_n1090), .C2(new_n1105), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1108), .B1(new_n1125), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1024), .B1(new_n978), .B2(new_n980), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1080), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n960), .B1(new_n1059), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n765), .A2(new_n951), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT46), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n950), .A2(new_n954), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1136), .A2(new_n950), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1139), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1140));
  XNOR2_X1  g715(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1140), .B(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n951), .B1(new_n953), .B2(new_n955), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n782), .A2(new_n784), .ZN(new_n1144));
  OAI22_X1  g719(.A1(new_n1143), .A2(new_n1144), .B1(G2067), .B2(new_n718), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n950), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n956), .A2(new_n950), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT126), .ZN(new_n1148));
  NOR2_X1   g723(.A1(G290), .A2(G1986), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n950), .A2(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT48), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n956), .A2(new_n1152), .A3(new_n950), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1148), .A2(new_n1151), .A3(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1142), .A2(new_n1146), .A3(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT127), .B1(new_n1135), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1094), .A2(new_n1105), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(KEYINPUT119), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1094), .A2(new_n1095), .A3(new_n1105), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1093), .A2(KEYINPUT60), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1093), .A2(KEYINPUT60), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n1112), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1113), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1161), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1160), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(KEYINPUT123), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1072), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1077), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1076), .B1(new_n1073), .B2(G171), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1172), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1069), .A2(new_n1060), .A3(new_n1070), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1171), .A2(new_n1133), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1169), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1034), .A2(new_n1058), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n959), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1155), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1156), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g759(.A1(G227), .A2(new_n463), .ZN(new_n1186));
  NAND2_X1  g760(.A1(new_n683), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g761(.A1(G401), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g762(.A(new_n1188), .B1(new_n857), .B2(new_n858), .ZN(new_n1189));
  NOR2_X1   g763(.A1(new_n919), .A2(new_n929), .ZN(new_n1190));
  NOR2_X1   g764(.A1(new_n1189), .A2(new_n1190), .ZN(G308));
  OAI221_X1 g765(.A(new_n1188), .B1(new_n857), .B2(new_n858), .C1(new_n919), .C2(new_n929), .ZN(G225));
endmodule


