

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769;

  NAND2_X2 U376 ( .A1(n636), .A2(G953), .ZN(n667) );
  XNOR2_X1 U377 ( .A(n424), .B(n590), .ZN(n768) );
  AND2_X1 U378 ( .A1(n594), .A2(n593), .ZN(n394) );
  XNOR2_X1 U379 ( .A(n589), .B(KEYINPUT41), .ZN(n710) );
  NAND2_X1 U380 ( .A1(n701), .A2(n698), .ZN(n589) );
  NOR2_X1 U381 ( .A1(n696), .A2(n697), .ZN(n701) );
  BUF_X1 U382 ( .A(n611), .Z(n354) );
  XNOR2_X1 U383 ( .A(n597), .B(n358), .ZN(n697) );
  INV_X1 U384 ( .A(KEYINPUT38), .ZN(n358) );
  XNOR2_X1 U385 ( .A(n586), .B(KEYINPUT1), .ZN(n611) );
  OR2_X1 U386 ( .A1(n672), .A2(G902), .ZN(n525) );
  XOR2_X1 U387 ( .A(KEYINPUT10), .B(n462), .Z(n753) );
  XNOR2_X1 U388 ( .A(KEYINPUT66), .B(KEYINPUT67), .ZN(n450) );
  NOR2_X1 U389 ( .A1(G953), .A2(G237), .ZN(n490) );
  XNOR2_X1 U390 ( .A(n357), .B(n470), .ZN(n654) );
  XNOR2_X1 U391 ( .A(n471), .B(n469), .ZN(n357) );
  XNOR2_X1 U392 ( .A(n471), .B(n452), .ZN(n642) );
  XNOR2_X2 U393 ( .A(n499), .B(n498), .ZN(n556) );
  XNOR2_X1 U394 ( .A(n368), .B(n404), .ZN(n627) );
  XNOR2_X2 U395 ( .A(n642), .B(n643), .ZN(n644) );
  XNOR2_X2 U396 ( .A(n633), .B(n632), .ZN(n634) );
  XOR2_X2 U397 ( .A(n480), .B(KEYINPUT94), .Z(n481) );
  XNOR2_X2 U398 ( .A(n405), .B(n505), .ZN(n650) );
  AND2_X4 U399 ( .A1(n411), .A2(n415), .ZN(n663) );
  XNOR2_X2 U400 ( .A(n625), .B(KEYINPUT76), .ZN(n411) );
  XNOR2_X2 U401 ( .A(n355), .B(n550), .ZN(n711) );
  NAND2_X2 U402 ( .A1(n549), .A2(n605), .ZN(n355) );
  NAND2_X2 U403 ( .A1(n356), .A2(n567), .ZN(n568) );
  XNOR2_X2 U404 ( .A(n561), .B(KEYINPUT87), .ZN(n356) );
  XNOR2_X2 U405 ( .A(n574), .B(n527), .ZN(n605) );
  NOR2_X1 U406 ( .A1(n768), .A2(n765), .ZN(n370) );
  INV_X1 U407 ( .A(G953), .ZN(n514) );
  BUF_X1 U408 ( .A(G128), .Z(n360) );
  AND2_X2 U409 ( .A1(n401), .A2(n361), .ZN(n400) );
  NAND2_X1 U410 ( .A1(n437), .A2(n434), .ZN(n574) );
  INV_X1 U411 ( .A(KEYINPUT48), .ZN(n404) );
  NOR2_X2 U412 ( .A1(n391), .A2(n683), .ZN(n735) );
  XNOR2_X1 U413 ( .A(n609), .B(n608), .ZN(n391) );
  NOR2_X1 U414 ( .A1(n684), .A2(n382), .ZN(n598) );
  NAND2_X1 U415 ( .A1(n410), .A2(n535), .ZN(n409) );
  AND2_X1 U416 ( .A1(n556), .A2(n536), .ZN(n606) );
  AND2_X1 U417 ( .A1(n439), .A2(n438), .ZN(n437) );
  XNOR2_X1 U418 ( .A(n508), .B(G478), .ZN(n535) );
  NOR2_X1 U419 ( .A1(n664), .A2(G902), .ZN(n461) );
  XNOR2_X1 U420 ( .A(n443), .B(n413), .ZN(n738) );
  XNOR2_X1 U421 ( .A(n450), .B(G131), .ZN(n486) );
  XNOR2_X1 U422 ( .A(KEYINPUT88), .B(KEYINPUT36), .ZN(n608) );
  XNOR2_X1 U423 ( .A(G140), .B(G137), .ZN(n519) );
  INV_X1 U424 ( .A(n744), .ZN(n359) );
  NAND2_X1 U425 ( .A1(n371), .A2(n369), .ZN(n368) );
  XNOR2_X1 U426 ( .A(n370), .B(KEYINPUT46), .ZN(n369) );
  XNOR2_X2 U427 ( .A(n512), .B(KEYINPUT22), .ZN(n547) );
  INV_X1 U428 ( .A(n738), .ZN(n423) );
  AND2_X1 U429 ( .A1(n432), .A2(n440), .ZN(n431) );
  NOR2_X1 U430 ( .A1(n437), .A2(KEYINPUT30), .ZN(n430) );
  XNOR2_X1 U431 ( .A(n394), .B(KEYINPUT73), .ZN(n393) );
  XNOR2_X1 U432 ( .A(n735), .B(n390), .ZN(n389) );
  INV_X1 U433 ( .A(KEYINPUT86), .ZN(n390) );
  XNOR2_X1 U434 ( .A(n584), .B(KEYINPUT69), .ZN(n604) );
  NAND2_X1 U435 ( .A1(n576), .A2(n611), .ZN(n396) );
  NAND2_X1 U436 ( .A1(n441), .A2(G902), .ZN(n438) );
  XNOR2_X1 U437 ( .A(n455), .B(n380), .ZN(n379) );
  XNOR2_X1 U438 ( .A(G110), .B(KEYINPUT24), .ZN(n455) );
  XNOR2_X1 U439 ( .A(KEYINPUT95), .B(KEYINPUT23), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n507), .B(n503), .ZN(n407) );
  XNOR2_X1 U441 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n501) );
  XNOR2_X1 U442 ( .A(n377), .B(n376), .ZN(n504) );
  INV_X1 U443 ( .A(KEYINPUT8), .ZN(n376) );
  XNOR2_X1 U444 ( .A(n421), .B(G107), .ZN(n500) );
  INV_X1 U445 ( .A(G116), .ZN(n421) );
  XNOR2_X1 U446 ( .A(G107), .B(G104), .ZN(n515) );
  XNOR2_X1 U447 ( .A(n386), .B(G146), .ZN(n385) );
  XNOR2_X1 U448 ( .A(n419), .B(KEYINPUT75), .ZN(n516) );
  INV_X1 U449 ( .A(G110), .ZN(n419) );
  XNOR2_X1 U450 ( .A(n381), .B(KEYINPUT39), .ZN(n619) );
  NAND2_X1 U451 ( .A1(n580), .A2(n598), .ZN(n381) );
  INV_X1 U452 ( .A(KEYINPUT68), .ZN(n610) );
  AND2_X1 U453 ( .A1(n603), .A2(n393), .ZN(n392) );
  XOR2_X1 U454 ( .A(KEYINPUT12), .B(KEYINPUT97), .Z(n489) );
  XNOR2_X1 U455 ( .A(KEYINPUT100), .B(KEYINPUT98), .ZN(n488) );
  OR2_X1 U456 ( .A1(G902), .A2(G237), .ZN(n474) );
  XNOR2_X1 U457 ( .A(G116), .B(G146), .ZN(n447) );
  XNOR2_X1 U458 ( .A(G143), .B(G113), .ZN(n484) );
  XOR2_X1 U459 ( .A(KEYINPUT99), .B(G140), .Z(n485) );
  NAND2_X1 U460 ( .A1(G237), .A2(G234), .ZN(n477) );
  XNOR2_X1 U461 ( .A(n537), .B(KEYINPUT105), .ZN(n700) );
  NOR2_X1 U462 ( .A1(n606), .A2(n618), .ZN(n537) );
  NAND2_X1 U463 ( .A1(n399), .A2(n398), .ZN(n397) );
  NOR2_X1 U464 ( .A1(n696), .A2(KEYINPUT19), .ZN(n398) );
  OR2_X1 U465 ( .A1(n642), .A2(n435), .ZN(n434) );
  NAND2_X1 U466 ( .A1(n453), .A2(n436), .ZN(n435) );
  INV_X1 U467 ( .A(G902), .ZN(n436) );
  INV_X1 U468 ( .A(G122), .ZN(n422) );
  XNOR2_X1 U469 ( .A(G113), .B(KEYINPUT91), .ZN(n443) );
  XNOR2_X1 U470 ( .A(n414), .B(KEYINPUT3), .ZN(n413) );
  INV_X1 U471 ( .A(G119), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n396), .B(KEYINPUT107), .ZN(n549) );
  AND2_X1 U473 ( .A1(n604), .A2(n388), .ZN(n613) );
  AND2_X1 U474 ( .A1(n606), .A2(n605), .ZN(n388) );
  NOR2_X1 U475 ( .A1(n588), .A2(n587), .ZN(n591) );
  XNOR2_X1 U476 ( .A(n409), .B(n408), .ZN(n618) );
  INV_X1 U477 ( .A(KEYINPUT104), .ZN(n408) );
  XNOR2_X1 U478 ( .A(n613), .B(KEYINPUT112), .ZN(n607) );
  XNOR2_X1 U479 ( .A(n384), .B(n559), .ZN(n662) );
  NAND2_X1 U480 ( .A1(n558), .A2(n557), .ZN(n384) );
  NAND2_X1 U481 ( .A1(n395), .A2(n690), .ZN(n691) );
  OR2_X1 U482 ( .A1(n577), .A2(n578), .ZN(n382) );
  XNOR2_X1 U483 ( .A(n538), .B(KEYINPUT65), .ZN(n576) );
  XNOR2_X1 U484 ( .A(n420), .B(n417), .ZN(n739) );
  XNOR2_X1 U485 ( .A(n516), .B(n418), .ZN(n417) );
  XNOR2_X1 U486 ( .A(n483), .B(n500), .ZN(n420) );
  INV_X1 U487 ( .A(KEYINPUT16), .ZN(n418) );
  AND2_X1 U488 ( .A1(n504), .A2(G221), .ZN(n375) );
  XNOR2_X1 U489 ( .A(n456), .B(n379), .ZN(n378) );
  XNOR2_X1 U490 ( .A(n407), .B(n406), .ZN(n405) );
  XNOR2_X1 U491 ( .A(n500), .B(n366), .ZN(n406) );
  XNOR2_X1 U492 ( .A(n387), .B(n385), .ZN(n517) );
  XNOR2_X1 U493 ( .A(n516), .B(n515), .ZN(n387) );
  XNOR2_X1 U494 ( .A(n654), .B(n655), .ZN(n656) );
  XNOR2_X1 U495 ( .A(n426), .B(n425), .ZN(n765) );
  XNOR2_X1 U496 ( .A(KEYINPUT110), .B(KEYINPUT40), .ZN(n425) );
  OR2_X1 U497 ( .A1(n433), .A2(n476), .ZN(n361) );
  XNOR2_X1 U498 ( .A(n460), .B(n459), .ZN(n362) );
  XNOR2_X1 U499 ( .A(n422), .B(G104), .ZN(n483) );
  AND2_X1 U500 ( .A1(n399), .A2(n433), .ZN(n363) );
  AND2_X1 U501 ( .A1(n434), .A2(n428), .ZN(n364) );
  AND2_X1 U502 ( .A1(n383), .A2(n442), .ZN(n365) );
  XOR2_X1 U503 ( .A(G134), .B(G122), .Z(n366) );
  INV_X1 U504 ( .A(KEYINPUT30), .ZN(n440) );
  INV_X1 U505 ( .A(KEYINPUT19), .ZN(n476) );
  XNOR2_X1 U506 ( .A(n372), .B(n610), .ZN(n371) );
  NAND2_X1 U507 ( .A1(n400), .A2(n397), .ZN(n367) );
  NAND2_X1 U508 ( .A1(n400), .A2(n397), .ZN(n592) );
  XNOR2_X2 U509 ( .A(n530), .B(KEYINPUT32), .ZN(n562) );
  XNOR2_X1 U510 ( .A(n378), .B(n375), .ZN(n457) );
  BUF_X1 U511 ( .A(n662), .Z(n403) );
  BUF_X1 U512 ( .A(n540), .Z(n552) );
  BUF_X1 U513 ( .A(n579), .Z(n597) );
  NAND2_X1 U514 ( .A1(n392), .A2(n389), .ZN(n372) );
  INV_X1 U515 ( .A(n374), .ZN(n583) );
  NAND2_X1 U516 ( .A1(n374), .A2(n681), .ZN(n538) );
  XNOR2_X2 U517 ( .A(n461), .B(n362), .ZN(n374) );
  AND2_X1 U518 ( .A1(n583), .A2(n373), .ZN(n682) );
  INV_X1 U519 ( .A(n681), .ZN(n373) );
  NOR2_X1 U520 ( .A1(n605), .A2(n374), .ZN(n528) );
  NAND2_X1 U521 ( .A1(n544), .A2(n374), .ZN(n545) );
  NAND2_X1 U522 ( .A1(n514), .A2(G234), .ZN(n377) );
  NAND2_X1 U523 ( .A1(n662), .A2(KEYINPUT44), .ZN(n383) );
  NAND2_X1 U524 ( .A1(n514), .A2(G227), .ZN(n386) );
  INV_X1 U525 ( .A(n396), .ZN(n395) );
  INV_X1 U526 ( .A(n579), .ZN(n399) );
  NAND2_X1 U527 ( .A1(n579), .A2(KEYINPUT19), .ZN(n401) );
  NAND2_X1 U528 ( .A1(n592), .A2(n481), .ZN(n482) );
  AND2_X1 U529 ( .A1(n631), .A2(n630), .ZN(n415) );
  NAND2_X1 U530 ( .A1(n663), .A2(G478), .ZN(n651) );
  NAND2_X1 U531 ( .A1(n560), .A2(n365), .ZN(n561) );
  INV_X1 U532 ( .A(n535), .ZN(n536) );
  INV_X1 U533 ( .A(n409), .ZN(n731) );
  INV_X1 U534 ( .A(n556), .ZN(n410) );
  NAND2_X1 U535 ( .A1(n680), .A2(n411), .ZN(n716) );
  XNOR2_X2 U536 ( .A(n412), .B(n473), .ZN(n579) );
  NAND2_X1 U537 ( .A1(n654), .A2(n472), .ZN(n412) );
  XNOR2_X1 U538 ( .A(n497), .B(n496), .ZN(n633) );
  XOR2_X2 U539 ( .A(G146), .B(G125), .Z(n462) );
  XNOR2_X2 U540 ( .A(n518), .B(n423), .ZN(n471) );
  XNOR2_X2 U541 ( .A(n752), .B(G101), .ZN(n518) );
  XNOR2_X2 U542 ( .A(n506), .B(KEYINPUT4), .ZN(n752) );
  XNOR2_X2 U543 ( .A(G143), .B(G128), .ZN(n506) );
  NAND2_X1 U544 ( .A1(n710), .A2(n591), .ZN(n424) );
  AND2_X1 U545 ( .A1(n619), .A2(n606), .ZN(n426) );
  NAND2_X1 U546 ( .A1(n429), .A2(n427), .ZN(n575) );
  NAND2_X1 U547 ( .A1(n437), .A2(n364), .ZN(n427) );
  NOR2_X1 U548 ( .A1(n696), .A2(n440), .ZN(n428) );
  NOR2_X1 U549 ( .A1(n431), .A2(n430), .ZN(n429) );
  NAND2_X1 U550 ( .A1(n434), .A2(n433), .ZN(n432) );
  INV_X1 U551 ( .A(n696), .ZN(n433) );
  NAND2_X1 U552 ( .A1(n642), .A2(n441), .ZN(n439) );
  INV_X1 U553 ( .A(n453), .ZN(n441) );
  BUF_X1 U554 ( .A(n663), .Z(n669) );
  AND2_X1 U555 ( .A1(n548), .A2(n641), .ZN(n442) );
  XNOR2_X1 U556 ( .A(n700), .B(KEYINPUT82), .ZN(n593) );
  INV_X1 U557 ( .A(n727), .ZN(n601) );
  AND2_X1 U558 ( .A1(n602), .A2(n601), .ZN(n603) );
  INV_X1 U559 ( .A(G137), .ZN(n446) );
  XNOR2_X1 U560 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U561 ( .A(n449), .B(n448), .ZN(n451) );
  INV_X1 U562 ( .A(KEYINPUT84), .ZN(n622) );
  XNOR2_X1 U563 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U564 ( .A(KEYINPUT74), .B(KEYINPUT5), .Z(n445) );
  NAND2_X1 U565 ( .A1(G210), .A2(n490), .ZN(n444) );
  XNOR2_X1 U566 ( .A(n445), .B(n444), .ZN(n449) );
  XNOR2_X1 U567 ( .A(n486), .B(G134), .ZN(n520) );
  XNOR2_X1 U568 ( .A(n451), .B(n520), .ZN(n452) );
  XNOR2_X1 U569 ( .A(KEYINPUT96), .B(G472), .ZN(n453) );
  XNOR2_X1 U570 ( .A(n360), .B(G119), .ZN(n454) );
  XNOR2_X1 U571 ( .A(n454), .B(n519), .ZN(n456) );
  XNOR2_X1 U572 ( .A(n457), .B(n753), .ZN(n664) );
  XOR2_X1 U573 ( .A(KEYINPUT25), .B(KEYINPUT77), .Z(n460) );
  XNOR2_X1 U574 ( .A(n436), .B(KEYINPUT15), .ZN(n630) );
  INV_X1 U575 ( .A(n630), .ZN(n472) );
  NAND2_X1 U576 ( .A1(G234), .A2(n472), .ZN(n458) );
  XNOR2_X1 U577 ( .A(KEYINPUT20), .B(n458), .ZN(n509) );
  NAND2_X1 U578 ( .A1(n509), .A2(G217), .ZN(n459) );
  XNOR2_X1 U579 ( .A(n739), .B(n462), .ZN(n470) );
  XOR2_X1 U580 ( .A(KEYINPUT90), .B(KEYINPUT17), .Z(n464) );
  NAND2_X1 U581 ( .A1(G224), .A2(n514), .ZN(n463) );
  XNOR2_X1 U582 ( .A(n464), .B(n463), .ZN(n468) );
  XOR2_X1 U583 ( .A(KEYINPUT18), .B(KEYINPUT78), .Z(n466) );
  XNOR2_X1 U584 ( .A(KEYINPUT92), .B(KEYINPUT79), .ZN(n465) );
  XNOR2_X1 U585 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U586 ( .A(n468), .B(n467), .Z(n469) );
  NAND2_X1 U587 ( .A1(n474), .A2(G210), .ZN(n473) );
  NAND2_X1 U588 ( .A1(G214), .A2(n474), .ZN(n475) );
  XNOR2_X1 U589 ( .A(KEYINPUT93), .B(n475), .ZN(n696) );
  XNOR2_X1 U590 ( .A(n477), .B(KEYINPUT14), .ZN(n478) );
  NAND2_X1 U591 ( .A1(G952), .A2(n478), .ZN(n708) );
  NOR2_X1 U592 ( .A1(G953), .A2(n708), .ZN(n572) );
  NAND2_X1 U593 ( .A1(G902), .A2(n478), .ZN(n569) );
  OR2_X1 U594 ( .A1(n514), .A2(G898), .ZN(n742) );
  NOR2_X1 U595 ( .A1(n569), .A2(n742), .ZN(n479) );
  NOR2_X1 U596 ( .A1(n572), .A2(n479), .ZN(n480) );
  XNOR2_X2 U597 ( .A(n482), .B(KEYINPUT0), .ZN(n540) );
  XNOR2_X1 U598 ( .A(n753), .B(n483), .ZN(n497) );
  XNOR2_X1 U599 ( .A(n485), .B(n484), .ZN(n487) );
  XNOR2_X1 U600 ( .A(n486), .B(n487), .ZN(n495) );
  XNOR2_X1 U601 ( .A(n489), .B(n488), .ZN(n493) );
  NAND2_X1 U602 ( .A1(n490), .A2(G214), .ZN(n491) );
  XNOR2_X1 U603 ( .A(n491), .B(KEYINPUT11), .ZN(n492) );
  XNOR2_X1 U604 ( .A(n492), .B(n493), .ZN(n494) );
  NAND2_X1 U605 ( .A1(n633), .A2(n436), .ZN(n499) );
  XOR2_X1 U606 ( .A(KEYINPUT13), .B(G475), .Z(n498) );
  XOR2_X1 U607 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n502) );
  XNOR2_X1 U608 ( .A(n502), .B(n501), .ZN(n503) );
  NAND2_X1 U609 ( .A1(G217), .A2(n504), .ZN(n505) );
  XNOR2_X1 U610 ( .A(n506), .B(KEYINPUT101), .ZN(n507) );
  NAND2_X1 U611 ( .A1(n650), .A2(n436), .ZN(n508) );
  NOR2_X1 U612 ( .A1(n556), .A2(n535), .ZN(n698) );
  NAND2_X1 U613 ( .A1(n509), .A2(G221), .ZN(n510) );
  XOR2_X1 U614 ( .A(KEYINPUT21), .B(n510), .Z(n681) );
  NAND2_X1 U615 ( .A1(n698), .A2(n681), .ZN(n511) );
  NOR2_X2 U616 ( .A1(n540), .A2(n511), .ZN(n512) );
  AND2_X1 U617 ( .A1(n547), .A2(n583), .ZN(n513) );
  NAND2_X1 U618 ( .A1(n574), .A2(n513), .ZN(n563) );
  XNOR2_X1 U619 ( .A(n518), .B(n517), .ZN(n521) );
  XNOR2_X1 U620 ( .A(n520), .B(n519), .ZN(n754) );
  XNOR2_X1 U621 ( .A(n521), .B(n754), .ZN(n672) );
  XNOR2_X1 U622 ( .A(KEYINPUT71), .B(G469), .ZN(n523) );
  INV_X1 U623 ( .A(KEYINPUT70), .ZN(n522) );
  XNOR2_X1 U624 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X2 U625 ( .A(n525), .B(n524), .ZN(n586) );
  INV_X1 U626 ( .A(KEYINPUT44), .ZN(n531) );
  OR2_X1 U627 ( .A1(n354), .A2(n531), .ZN(n526) );
  NOR2_X1 U628 ( .A1(n563), .A2(n526), .ZN(n533) );
  XNOR2_X1 U629 ( .A(KEYINPUT106), .B(KEYINPUT6), .ZN(n527) );
  AND2_X1 U630 ( .A1(n528), .A2(n354), .ZN(n529) );
  NAND2_X1 U631 ( .A1(n547), .A2(n529), .ZN(n530) );
  NOR2_X1 U632 ( .A1(n562), .A2(n531), .ZN(n532) );
  NOR2_X1 U633 ( .A1(n532), .A2(n533), .ZN(n534) );
  XNOR2_X1 U634 ( .A(n534), .B(KEYINPUT64), .ZN(n560) );
  INV_X1 U635 ( .A(n574), .ZN(n690) );
  NOR2_X1 U636 ( .A1(n540), .A2(n691), .ZN(n539) );
  XOR2_X1 U637 ( .A(KEYINPUT31), .B(n539), .Z(n732) );
  NAND2_X1 U638 ( .A1(n574), .A2(n576), .ZN(n541) );
  INV_X1 U639 ( .A(n586), .ZN(n578) );
  OR2_X1 U640 ( .A1(n541), .A2(n578), .ZN(n542) );
  NOR2_X1 U641 ( .A1(n552), .A2(n542), .ZN(n720) );
  OR2_X1 U642 ( .A1(n732), .A2(n720), .ZN(n543) );
  NAND2_X1 U643 ( .A1(n593), .A2(n543), .ZN(n548) );
  INV_X1 U644 ( .A(n605), .ZN(n544) );
  NOR2_X1 U645 ( .A1(n545), .A2(n354), .ZN(n546) );
  NAND2_X1 U646 ( .A1(n547), .A2(n546), .ZN(n641) );
  XNOR2_X1 U647 ( .A(KEYINPUT72), .B(KEYINPUT33), .ZN(n550) );
  INV_X1 U648 ( .A(n552), .ZN(n553) );
  NAND2_X1 U649 ( .A1(n711), .A2(n553), .ZN(n555) );
  INV_X1 U650 ( .A(KEYINPUT34), .ZN(n554) );
  XNOR2_X1 U651 ( .A(n555), .B(n554), .ZN(n558) );
  NAND2_X1 U652 ( .A1(n535), .A2(n556), .ZN(n600) );
  INV_X1 U653 ( .A(n600), .ZN(n557) );
  XNOR2_X1 U654 ( .A(KEYINPUT80), .B(KEYINPUT35), .ZN(n559) );
  BUF_X1 U655 ( .A(n562), .Z(n767) );
  OR2_X1 U656 ( .A1(n563), .A2(n354), .ZN(n724) );
  NAND2_X1 U657 ( .A1(n767), .A2(n724), .ZN(n564) );
  NOR2_X1 U658 ( .A1(n564), .A2(KEYINPUT44), .ZN(n566) );
  INV_X1 U659 ( .A(n403), .ZN(n565) );
  NAND2_X1 U660 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X2 U661 ( .A(n568), .B(KEYINPUT45), .ZN(n743) );
  OR2_X1 U662 ( .A1(n514), .A2(n569), .ZN(n570) );
  NOR2_X1 U663 ( .A1(G900), .A2(n570), .ZN(n571) );
  NOR2_X1 U664 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U665 ( .A(KEYINPUT81), .B(n573), .ZN(n581) );
  NAND2_X1 U666 ( .A1(n581), .A2(n575), .ZN(n577) );
  INV_X1 U667 ( .A(n576), .ZN(n684) );
  INV_X1 U668 ( .A(n697), .ZN(n580) );
  XNOR2_X1 U669 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n590) );
  AND2_X1 U670 ( .A1(n681), .A2(n581), .ZN(n582) );
  NAND2_X1 U671 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U672 ( .A1(n604), .A2(n690), .ZN(n585) );
  XNOR2_X1 U673 ( .A(n585), .B(KEYINPUT28), .ZN(n588) );
  XNOR2_X1 U674 ( .A(n586), .B(KEYINPUT109), .ZN(n587) );
  NAND2_X1 U675 ( .A1(n367), .A2(n591), .ZN(n595) );
  NOR2_X1 U676 ( .A1(KEYINPUT47), .A2(n595), .ZN(n594) );
  INV_X1 U677 ( .A(n595), .ZN(n728) );
  NAND2_X1 U678 ( .A1(n700), .A2(n728), .ZN(n596) );
  NAND2_X1 U679 ( .A1(n596), .A2(KEYINPUT47), .ZN(n602) );
  INV_X1 U680 ( .A(n597), .ZN(n616) );
  NAND2_X1 U681 ( .A1(n616), .A2(n598), .ZN(n599) );
  NOR2_X1 U682 ( .A1(n600), .A2(n599), .ZN(n727) );
  NAND2_X1 U683 ( .A1(n607), .A2(n363), .ZN(n609) );
  INV_X1 U684 ( .A(n354), .ZN(n683) );
  NOR2_X1 U685 ( .A1(n354), .A2(n696), .ZN(n612) );
  AND2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U687 ( .A(n614), .B(KEYINPUT43), .ZN(n615) );
  NOR2_X1 U688 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U689 ( .A(n617), .B(KEYINPUT108), .ZN(n766) );
  NAND2_X1 U690 ( .A1(n619), .A2(n618), .ZN(n737) );
  INV_X1 U691 ( .A(n737), .ZN(n620) );
  NOR2_X1 U692 ( .A1(n766), .A2(n620), .ZN(n626) );
  AND2_X1 U693 ( .A1(n626), .A2(KEYINPUT2), .ZN(n621) );
  NAND2_X1 U694 ( .A1(n627), .A2(n621), .ZN(n623) );
  XNOR2_X1 U695 ( .A(n623), .B(n622), .ZN(n624) );
  NAND2_X1 U696 ( .A1(n743), .A2(n624), .ZN(n625) );
  AND2_X1 U697 ( .A1(n627), .A2(n626), .ZN(n756) );
  NAND2_X1 U698 ( .A1(n743), .A2(n756), .ZN(n629) );
  INV_X1 U699 ( .A(KEYINPUT2), .ZN(n628) );
  NAND2_X1 U700 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U701 ( .A1(n663), .A2(G475), .ZN(n635) );
  XOR2_X1 U702 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n632) );
  XNOR2_X1 U703 ( .A(n635), .B(n634), .ZN(n637) );
  INV_X1 U704 ( .A(G952), .ZN(n636) );
  NAND2_X1 U705 ( .A1(n637), .A2(n667), .ZN(n639) );
  INV_X1 U706 ( .A(KEYINPUT60), .ZN(n638) );
  XNOR2_X1 U707 ( .A(n639), .B(n638), .ZN(G60) );
  XOR2_X1 U708 ( .A(G101), .B(KEYINPUT115), .Z(n640) );
  XNOR2_X1 U709 ( .A(n641), .B(n640), .ZN(G3) );
  NAND2_X1 U710 ( .A1(n663), .A2(G472), .ZN(n645) );
  XNOR2_X1 U711 ( .A(KEYINPUT113), .B(KEYINPUT62), .ZN(n643) );
  XNOR2_X1 U712 ( .A(n645), .B(n644), .ZN(n646) );
  NAND2_X1 U713 ( .A1(n646), .A2(n667), .ZN(n649) );
  XOR2_X1 U714 ( .A(KEYINPUT114), .B(KEYINPUT63), .Z(n647) );
  XNOR2_X1 U715 ( .A(n647), .B(KEYINPUT89), .ZN(n648) );
  XNOR2_X1 U716 ( .A(n649), .B(n648), .ZN(G57) );
  XNOR2_X1 U717 ( .A(n651), .B(n650), .ZN(n652) );
  NAND2_X1 U718 ( .A1(n652), .A2(n667), .ZN(n653) );
  XNOR2_X1 U719 ( .A(n653), .B(KEYINPUT121), .ZN(G63) );
  NAND2_X1 U720 ( .A1(n663), .A2(G210), .ZN(n657) );
  XOR2_X1 U721 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n655) );
  XNOR2_X1 U722 ( .A(n657), .B(n656), .ZN(n658) );
  NAND2_X1 U723 ( .A1(n658), .A2(n667), .ZN(n660) );
  XNOR2_X1 U724 ( .A(KEYINPUT85), .B(KEYINPUT56), .ZN(n659) );
  XNOR2_X1 U725 ( .A(n660), .B(n659), .ZN(G51) );
  XOR2_X1 U726 ( .A(G122), .B(KEYINPUT126), .Z(n661) );
  XNOR2_X1 U727 ( .A(n403), .B(n661), .ZN(G24) );
  NAND2_X1 U728 ( .A1(n669), .A2(G217), .ZN(n666) );
  XNOR2_X1 U729 ( .A(n664), .B(KEYINPUT122), .ZN(n665) );
  XNOR2_X1 U730 ( .A(n666), .B(n665), .ZN(n668) );
  INV_X1 U731 ( .A(n667), .ZN(n675) );
  NOR2_X1 U732 ( .A1(n668), .A2(n675), .ZN(G66) );
  NAND2_X1 U733 ( .A1(n669), .A2(G469), .ZN(n674) );
  XNOR2_X1 U734 ( .A(KEYINPUT119), .B(KEYINPUT57), .ZN(n670) );
  XNOR2_X1 U735 ( .A(n670), .B(KEYINPUT58), .ZN(n671) );
  XNOR2_X1 U736 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U737 ( .A(n674), .B(n673), .ZN(n676) );
  NOR2_X1 U738 ( .A1(n676), .A2(n675), .ZN(G54) );
  NOR2_X1 U739 ( .A1(n359), .A2(KEYINPUT2), .ZN(n679) );
  NOR2_X1 U740 ( .A1(n756), .A2(KEYINPUT2), .ZN(n677) );
  XOR2_X1 U741 ( .A(KEYINPUT83), .B(n677), .Z(n678) );
  NOR2_X1 U742 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U743 ( .A(KEYINPUT49), .B(n682), .ZN(n688) );
  NAND2_X1 U744 ( .A1(n684), .A2(n683), .ZN(n686) );
  XOR2_X1 U745 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n685) );
  XNOR2_X1 U746 ( .A(n686), .B(n685), .ZN(n687) );
  NAND2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U748 ( .A1(n690), .A2(n689), .ZN(n693) );
  INV_X1 U749 ( .A(n691), .ZN(n692) );
  NOR2_X1 U750 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U751 ( .A(KEYINPUT51), .B(n694), .ZN(n695) );
  NAND2_X1 U752 ( .A1(n695), .A2(n710), .ZN(n706) );
  NAND2_X1 U753 ( .A1(n697), .A2(n696), .ZN(n699) );
  NAND2_X1 U754 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U755 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U756 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U757 ( .A1(n704), .A2(n711), .ZN(n705) );
  NAND2_X1 U758 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U759 ( .A(KEYINPUT52), .B(n707), .Z(n709) );
  NOR2_X1 U760 ( .A1(n709), .A2(n708), .ZN(n714) );
  NAND2_X1 U761 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U762 ( .A1(n712), .A2(n514), .ZN(n713) );
  NOR2_X1 U763 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U764 ( .A1(n716), .A2(n715), .ZN(n718) );
  XOR2_X1 U765 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n717) );
  XNOR2_X1 U766 ( .A(n718), .B(n717), .ZN(G75) );
  NAND2_X1 U767 ( .A1(n720), .A2(n606), .ZN(n719) );
  XNOR2_X1 U768 ( .A(n719), .B(G104), .ZN(G6) );
  XOR2_X1 U769 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n722) );
  NAND2_X1 U770 ( .A1(n720), .A2(n731), .ZN(n721) );
  XNOR2_X1 U771 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U772 ( .A(G107), .B(n723), .ZN(G9) );
  XNOR2_X1 U773 ( .A(G110), .B(n724), .ZN(G12) );
  XOR2_X1 U774 ( .A(n360), .B(KEYINPUT29), .Z(n726) );
  NAND2_X1 U775 ( .A1(n728), .A2(n731), .ZN(n725) );
  XNOR2_X1 U776 ( .A(n726), .B(n725), .ZN(G30) );
  XOR2_X1 U777 ( .A(G143), .B(n727), .Z(G45) );
  NAND2_X1 U778 ( .A1(n728), .A2(n606), .ZN(n729) );
  XNOR2_X1 U779 ( .A(n729), .B(G146), .ZN(G48) );
  NAND2_X1 U780 ( .A1(n606), .A2(n732), .ZN(n730) );
  XNOR2_X1 U781 ( .A(G113), .B(n730), .ZN(G15) );
  NAND2_X1 U782 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U783 ( .A(n733), .B(KEYINPUT116), .ZN(n734) );
  XNOR2_X1 U784 ( .A(G116), .B(n734), .ZN(G18) );
  XNOR2_X1 U785 ( .A(n735), .B(G125), .ZN(n736) );
  XNOR2_X1 U786 ( .A(n736), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U787 ( .A(G134), .B(n737), .ZN(G36) );
  XNOR2_X1 U788 ( .A(G101), .B(n738), .ZN(n740) );
  XNOR2_X1 U789 ( .A(n740), .B(n739), .ZN(n741) );
  NAND2_X1 U790 ( .A1(n742), .A2(n741), .ZN(n751) );
  INV_X1 U791 ( .A(n743), .ZN(n744) );
  NOR2_X1 U792 ( .A1(n744), .A2(G953), .ZN(n749) );
  NAND2_X1 U793 ( .A1(G953), .A2(G224), .ZN(n745) );
  XNOR2_X1 U794 ( .A(KEYINPUT61), .B(n745), .ZN(n746) );
  NAND2_X1 U795 ( .A1(n746), .A2(G898), .ZN(n747) );
  XNOR2_X1 U796 ( .A(n747), .B(KEYINPUT123), .ZN(n748) );
  NOR2_X1 U797 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U798 ( .A(n751), .B(n750), .ZN(G69) );
  XNOR2_X1 U799 ( .A(n752), .B(n753), .ZN(n755) );
  XNOR2_X1 U800 ( .A(n755), .B(n754), .ZN(n759) );
  XOR2_X1 U801 ( .A(KEYINPUT124), .B(n756), .Z(n757) );
  XNOR2_X1 U802 ( .A(n759), .B(n757), .ZN(n758) );
  NAND2_X1 U803 ( .A1(n758), .A2(n514), .ZN(n764) );
  XNOR2_X1 U804 ( .A(G227), .B(n759), .ZN(n760) );
  NAND2_X1 U805 ( .A1(n760), .A2(G900), .ZN(n761) );
  XOR2_X1 U806 ( .A(KEYINPUT125), .B(n761), .Z(n762) );
  NAND2_X1 U807 ( .A1(G953), .A2(n762), .ZN(n763) );
  NAND2_X1 U808 ( .A1(n764), .A2(n763), .ZN(G72) );
  XOR2_X1 U809 ( .A(G131), .B(n765), .Z(G33) );
  XOR2_X1 U810 ( .A(G140), .B(n766), .Z(G42) );
  XNOR2_X1 U811 ( .A(G119), .B(n767), .ZN(G21) );
  XNOR2_X1 U812 ( .A(G137), .B(KEYINPUT127), .ZN(n769) );
  XNOR2_X1 U813 ( .A(n769), .B(n768), .ZN(G39) );
endmodule

