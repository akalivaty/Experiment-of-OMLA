//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n531, new_n532, new_n533, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n545, new_n547, new_n548, new_n549, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1128, new_n1129, new_n1130,
    new_n1131;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT68), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n465), .A2(new_n471), .A3(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n462), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n468), .B2(new_n470), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n467), .A2(G2105), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n475), .A2(G137), .B1(G101), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n474), .A2(new_n478), .ZN(G160));
  AOI21_X1  g054(.A(new_n462), .B1(new_n468), .B2(new_n470), .ZN(new_n480));
  MUX2_X1   g055(.A(G100), .B(G112), .S(G2105), .Z(new_n481));
  AOI22_X1  g056(.A1(G124), .A2(new_n480), .B1(new_n481), .B2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n475), .A2(G136), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT69), .Z(G162));
  OAI21_X1  g060(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n488), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n489));
  AOI21_X1  g064(.A(KEYINPUT70), .B1(new_n488), .B2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(G138), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n496), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n465), .A2(new_n471), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n493), .B1(new_n495), .B2(new_n498), .ZN(G164));
  AND2_X1   g074(.A1(KEYINPUT6), .A2(G651), .ZN(new_n500));
  NOR2_X1   g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G50), .ZN(new_n505));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  INV_X1    g081(.A(new_n502), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n505), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n510), .A2(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  NAND2_X1  g090(.A1(new_n507), .A2(G89), .ZN(new_n516));
  NAND2_X1  g091(.A1(G63), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(new_n508), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n504), .A2(G51), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT71), .B(KEYINPUT7), .ZN(new_n522));
  AND3_X1   g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n522), .B(new_n523), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n519), .A2(new_n520), .A3(new_n521), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n521), .ZN(new_n526));
  XOR2_X1   g101(.A(KEYINPUT5), .B(G543), .Z(new_n527));
  AOI21_X1  g102(.A(new_n527), .B1(new_n516), .B2(new_n517), .ZN(new_n528));
  OAI21_X1  g103(.A(KEYINPUT72), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n525), .A2(new_n529), .ZN(G168));
  NOR2_X1   g105(.A1(new_n527), .A2(new_n502), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n531), .A2(G90), .B1(new_n504), .B2(G52), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n512), .B2(new_n533), .ZN(G301));
  INV_X1    g109(.A(G301), .ZN(G171));
  INV_X1    g110(.A(G81), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n507), .A2(G543), .ZN(new_n537));
  XOR2_X1   g112(.A(KEYINPUT73), .B(G43), .Z(new_n538));
  OAI22_X1  g113(.A1(new_n509), .A2(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n512), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  XOR2_X1   g117(.A(new_n542), .B(KEYINPUT74), .Z(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  AND3_X1   g119(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G36), .ZN(G176));
  XOR2_X1   g121(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n547));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n545), .A2(new_n549), .ZN(G188));
  INV_X1    g125(.A(G53), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT77), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n551), .B1(new_n552), .B2(KEYINPUT9), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n504), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT76), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n552), .B1(new_n555), .B2(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n556), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n504), .A2(new_n553), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g135(.A(KEYINPUT78), .B(G65), .Z(new_n561));
  AOI22_X1  g136(.A1(new_n561), .A2(new_n508), .B1(G78), .B2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G91), .ZN(new_n563));
  OAI22_X1  g138(.A1(new_n562), .A2(new_n512), .B1(new_n509), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(G299));
  INV_X1    g141(.A(G168), .ZN(G286));
  NAND2_X1  g142(.A1(new_n531), .A2(G87), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n504), .A2(G49), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  AOI22_X1  g146(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n512), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT79), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n573), .B(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n531), .A2(G86), .B1(new_n504), .B2(G48), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(G305));
  NAND2_X1  g152(.A1(G72), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G60), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n527), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT80), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n512), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n582), .B1(new_n581), .B2(new_n580), .ZN(new_n583));
  XNOR2_X1  g158(.A(KEYINPUT81), .B(G85), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n531), .A2(new_n584), .B1(new_n504), .B2(G47), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(G290));
  INV_X1    g161(.A(KEYINPUT10), .ZN(new_n587));
  INV_X1    g162(.A(G92), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n509), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n531), .A2(KEYINPUT10), .A3(G92), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n589), .A2(new_n590), .B1(G54), .B2(new_n504), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n508), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n512), .B1(new_n592), .B2(KEYINPUT82), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(KEYINPUT82), .B2(new_n592), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(new_n596), .B2(G301), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G284));
  XNOR2_X1  g174(.A(new_n598), .B(KEYINPUT83), .ZN(G321));
  OAI21_X1  g175(.A(KEYINPUT84), .B1(new_n565), .B2(G868), .ZN(new_n601));
  NOR2_X1   g176(.A1(G168), .A2(new_n596), .ZN(new_n602));
  MUX2_X1   g177(.A(new_n601), .B(KEYINPUT84), .S(new_n602), .Z(G297));
  XOR2_X1   g178(.A(G297), .B(KEYINPUT85), .Z(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n595), .B1(new_n605), .B2(G860), .ZN(G148));
  INV_X1    g181(.A(new_n595), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(G559), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(new_n596), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(new_n596), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g187(.A1(new_n465), .A2(new_n471), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(new_n476), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  INV_X1    g191(.A(G2100), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  AOI22_X1  g194(.A1(G123), .A2(new_n480), .B1(new_n475), .B2(G135), .ZN(new_n620));
  NOR3_X1   g195(.A1(new_n462), .A2(KEYINPUT86), .A3(G111), .ZN(new_n621));
  OAI21_X1  g196(.A(KEYINPUT86), .B1(new_n462), .B2(G111), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n622), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n620), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(G2096), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n618), .A2(new_n619), .A3(new_n626), .ZN(G156));
  XOR2_X1   g202(.A(G2451), .B(G2454), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT87), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT15), .B(G2435), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2438), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2427), .Z(new_n637));
  OAI21_X1  g212(.A(KEYINPUT14), .B1(new_n637), .B2(G2430), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n638), .B1(G2430), .B2(new_n637), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n634), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n634), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(new_n642), .A3(G14), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(G401));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  NOR3_X1   g224(.A1(new_n646), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT18), .ZN(new_n651));
  INV_X1    g226(.A(new_n647), .ZN(new_n652));
  AND2_X1   g227(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n648), .B1(new_n653), .B2(new_n645), .ZN(new_n654));
  INV_X1    g229(.A(new_n653), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n654), .B1(new_n646), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n646), .A2(new_n649), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n652), .B1(new_n657), .B2(KEYINPUT17), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n651), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(new_n625), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2100), .ZN(G227));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1956), .B(G2474), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1961), .B(G1966), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n663), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n663), .A2(new_n666), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT20), .Z(new_n670));
  AOI211_X1 g245(.A(new_n668), .B(new_n670), .C1(new_n663), .C2(new_n667), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT88), .Z(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1981), .B(G1986), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n674), .B(new_n677), .ZN(G229));
  NOR2_X1   g253(.A1(G6), .A2(G16), .ZN(new_n679));
  INV_X1    g254(.A(G305), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(G16), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT32), .B(G1981), .Z(new_n682));
  XOR2_X1   g257(.A(new_n681), .B(new_n682), .Z(new_n683));
  NOR2_X1   g258(.A1(G16), .A2(G23), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT92), .ZN(new_n685));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n685), .B1(G288), .B2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT33), .B(G1976), .Z(new_n688));
  XOR2_X1   g263(.A(new_n687), .B(new_n688), .Z(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(G22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT93), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(G303), .B2(G16), .ZN(new_n692));
  INV_X1    g267(.A(G1971), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n683), .A2(new_n689), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT91), .B(KEYINPUT34), .Z(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n699), .A2(KEYINPUT89), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(KEYINPUT89), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n702), .A2(G25), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n475), .A2(G131), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n480), .A2(G119), .ZN(new_n705));
  MUX2_X1   g280(.A(G95), .B(G107), .S(G2105), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G2104), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n703), .B1(new_n709), .B2(new_n702), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT90), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT35), .B(G1991), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  MUX2_X1   g288(.A(G24), .B(G290), .S(G16), .Z(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(G1986), .Z(new_n715));
  NAND4_X1  g290(.A1(new_n697), .A2(new_n698), .A3(new_n713), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT36), .ZN(new_n717));
  NOR2_X1   g292(.A1(G29), .A2(G33), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n476), .A2(G103), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT25), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n476), .A2(KEYINPUT25), .A3(G103), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n721), .A2(new_n722), .B1(G139), .B2(new_n475), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n613), .A2(G127), .ZN(new_n724));
  NAND2_X1  g299(.A1(G115), .A2(G2104), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n462), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT98), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n723), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n727), .B2(new_n726), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n718), .B1(new_n729), .B2(G29), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT99), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G2072), .ZN(new_n732));
  NOR2_X1   g307(.A1(G171), .A2(new_n686), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G5), .B2(new_n686), .ZN(new_n734));
  INV_X1    g309(.A(G1961), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n702), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT24), .B(G34), .ZN(new_n738));
  AOI22_X1  g313(.A1(G160), .A2(G29), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n699), .A2(G32), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT26), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n475), .A2(G141), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n480), .A2(G129), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI211_X1 g320(.A(new_n742), .B(new_n745), .C1(G105), .C2(new_n476), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n740), .B1(new_n746), .B2(new_n699), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT27), .B(G1996), .ZN(new_n749));
  OAI221_X1 g324(.A(new_n736), .B1(G2084), .B2(new_n739), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT100), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n702), .A2(G35), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G162), .B2(new_n702), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT29), .Z(new_n756));
  INV_X1    g331(.A(G2090), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n752), .A2(new_n753), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n686), .A2(G19), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n543), .B2(new_n686), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(G1341), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n737), .A2(G27), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT101), .Z(new_n764));
  INV_X1    g339(.A(G164), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(new_n702), .ZN(new_n766));
  INV_X1    g341(.A(G2078), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n734), .A2(new_n735), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n748), .A2(new_n749), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT31), .B(G11), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT30), .B(G28), .Z(new_n772));
  OAI221_X1 g347(.A(new_n771), .B1(G29), .B2(new_n772), .C1(new_n624), .C2(new_n737), .ZN(new_n773));
  NOR4_X1   g348(.A1(new_n768), .A2(new_n769), .A3(new_n770), .A4(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G4), .A2(G16), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT94), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n607), .B2(new_n686), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT95), .B(G1348), .Z(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G2084), .B2(new_n739), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n737), .A2(G26), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT28), .ZN(new_n782));
  AOI22_X1  g357(.A1(G128), .A2(new_n480), .B1(new_n475), .B2(G140), .ZN(new_n783));
  NOR2_X1   g358(.A1(G104), .A2(G2105), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT96), .ZN(new_n785));
  OAI21_X1  g360(.A(G2104), .B1(new_n462), .B2(G116), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n783), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AND3_X1   g362(.A1(new_n787), .A2(KEYINPUT97), .A3(G29), .ZN(new_n788));
  AOI21_X1  g363(.A(KEYINPUT97), .B1(new_n787), .B2(G29), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n782), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G2067), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n762), .A2(new_n774), .A3(new_n780), .A4(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n756), .A2(new_n757), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n686), .A2(G20), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT23), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n565), .B2(new_n686), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(G1956), .Z(new_n798));
  NOR2_X1   g373(.A1(G16), .A2(G21), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G168), .B2(G16), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(G1966), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(G1966), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n777), .A2(new_n778), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n798), .A2(new_n801), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  NOR4_X1   g379(.A1(new_n759), .A2(new_n793), .A3(new_n794), .A4(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n717), .A2(new_n732), .A3(new_n805), .ZN(G150));
  INV_X1    g381(.A(G150), .ZN(G311));
  NAND2_X1  g382(.A1(new_n504), .A2(G55), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT102), .B(G93), .Z(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n509), .B2(new_n809), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(new_n512), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(G860), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT37), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n595), .A2(G559), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT38), .Z(new_n818));
  INV_X1    g393(.A(new_n813), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n543), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(new_n542), .B2(new_n819), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n818), .B(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT39), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT103), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n826), .B(new_n814), .C1(new_n823), .C2(new_n822), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n824), .A2(new_n825), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n816), .B1(new_n827), .B2(new_n828), .ZN(G145));
  XNOR2_X1  g404(.A(new_n615), .B(new_n708), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n462), .A2(G106), .ZN(new_n831));
  NAND2_X1  g406(.A1(G118), .A2(G2105), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n467), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n480), .A2(G130), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT106), .Z(new_n835));
  AOI211_X1 g410(.A(new_n833), .B(new_n835), .C1(G142), .C2(new_n475), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n830), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n492), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT70), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n462), .B2(G114), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n488), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n486), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(KEYINPUT105), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n498), .A2(new_n495), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT105), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n491), .A2(new_n845), .A3(new_n492), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n787), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n837), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n729), .B(new_n746), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(G162), .B(new_n624), .ZN(new_n852));
  XNOR2_X1  g427(.A(G160), .B(KEYINPUT104), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(G37), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n854), .B2(new_n851), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g432(.A1(new_n595), .A2(G299), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n858), .A2(KEYINPUT107), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n595), .A2(G299), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n858), .B2(KEYINPUT107), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT41), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n821), .B(new_n609), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(new_n862), .B2(new_n864), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n866), .A2(KEYINPUT42), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(KEYINPUT42), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(G305), .B(G303), .ZN(new_n870));
  XOR2_X1   g445(.A(G290), .B(G288), .Z(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n867), .A2(new_n872), .A3(new_n868), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n596), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n819), .A2(G868), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(G295));
  NAND2_X1  g453(.A1(new_n874), .A2(new_n875), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(G868), .ZN(new_n880));
  INV_X1    g455(.A(new_n877), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n880), .A2(KEYINPUT108), .A3(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT108), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(new_n876), .B2(new_n877), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(G331));
  XNOR2_X1  g460(.A(G168), .B(G301), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n821), .B(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n863), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n862), .B2(new_n887), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n889), .A2(new_n872), .ZN(new_n890));
  INV_X1    g465(.A(G37), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n872), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n893), .A2(KEYINPUT43), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(KEYINPUT43), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n895), .B1(new_n894), .B2(new_n896), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(G397));
  INV_X1    g474(.A(KEYINPUT126), .ZN(new_n900));
  INV_X1    g475(.A(G1384), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n847), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT45), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n472), .A2(new_n473), .ZN(new_n905));
  OAI211_X1 g480(.A(G40), .B(new_n477), .C1(new_n905), .C2(new_n462), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n746), .B(G1996), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n787), .B(new_n791), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XOR2_X1   g485(.A(new_n708), .B(new_n712), .Z(new_n911));
  OAI21_X1  g486(.A(new_n907), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g487(.A1(G290), .A2(G1986), .ZN(new_n913));
  NOR2_X1   g488(.A1(G290), .A2(G1986), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n907), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  XOR2_X1   g491(.A(new_n916), .B(KEYINPUT109), .Z(new_n917));
  NAND2_X1  g492(.A1(new_n575), .A2(KEYINPUT111), .ZN(new_n918));
  NAND3_X1  g493(.A1(G305), .A2(new_n918), .A3(G1981), .ZN(new_n919));
  INV_X1    g494(.A(G1981), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n575), .B(new_n576), .C1(KEYINPUT111), .C2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT49), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n919), .A2(KEYINPUT49), .A3(new_n921), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n902), .A2(new_n906), .ZN(new_n926));
  INV_X1    g501(.A(G8), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n924), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n928), .ZN(new_n930));
  INV_X1    g505(.A(G1976), .ZN(new_n931));
  NOR2_X1   g506(.A1(G288), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT52), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT52), .B1(G288), .B2(new_n931), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n928), .B(new_n934), .C1(new_n931), .C2(G288), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n929), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  OAI211_X1 g511(.A(G303), .B(G8), .C1(KEYINPUT110), .C2(KEYINPUT55), .ZN(new_n937));
  NAND2_X1  g512(.A1(KEYINPUT110), .A2(KEYINPUT55), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n937), .B(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT50), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(G164), .B2(G1384), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n847), .A2(KEYINPUT50), .A3(new_n901), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n906), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n903), .B1(G164), .B2(G1384), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n847), .A2(KEYINPUT45), .A3(new_n901), .ZN(new_n946));
  INV_X1    g521(.A(G40), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n474), .A2(new_n478), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n757), .A2(new_n944), .B1(new_n949), .B2(new_n693), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n940), .B1(new_n950), .B2(new_n927), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n840), .A2(new_n841), .ZN(new_n952));
  AOI22_X1  g527(.A1(G126), .A2(new_n480), .B1(new_n952), .B2(new_n487), .ZN(new_n953));
  AOI21_X1  g528(.A(G1384), .B1(new_n844), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n954), .A2(new_n941), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n955), .A2(new_n906), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n847), .A2(new_n941), .A3(new_n901), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(new_n757), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n949), .A2(new_n693), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n927), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n940), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n936), .A2(new_n951), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n966), .A2(new_n957), .A3(new_n948), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n967), .A2(new_n778), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n902), .A2(new_n906), .A3(G2067), .ZN(new_n969));
  OAI211_X1 g544(.A(KEYINPUT60), .B(new_n595), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n969), .B1(new_n778), .B2(new_n967), .ZN(new_n971));
  OR2_X1    g546(.A1(new_n595), .A2(KEYINPUT60), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n595), .A2(KEYINPUT60), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n970), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G1996), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n945), .A2(new_n946), .A3(new_n976), .A4(new_n948), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT115), .ZN(new_n978));
  XOR2_X1   g553(.A(KEYINPUT58), .B(G1341), .Z(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n902), .B2(new_n906), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n978), .B1(new_n977), .B2(new_n980), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n543), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT59), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT59), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n985), .B(new_n543), .C1(new_n981), .C2(new_n982), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n975), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT57), .ZN(new_n988));
  INV_X1    g563(.A(new_n560), .ZN(new_n989));
  INV_X1    g564(.A(new_n564), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n560), .A2(KEYINPUT57), .A3(new_n564), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(KEYINPUT56), .B(G2072), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n945), .A2(new_n946), .A3(new_n948), .A4(new_n994), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n993), .B(new_n995), .C1(G1956), .C2(new_n944), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n995), .B1(new_n944), .B2(G1956), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n991), .A2(new_n992), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n997), .B2(new_n999), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n996), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT61), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n997), .A2(new_n999), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(new_n996), .A3(KEYINPUT61), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT117), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT117), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1005), .A2(new_n996), .A3(new_n1008), .A4(KEYINPUT61), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n987), .A2(new_n1004), .A3(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n971), .A2(new_n607), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1012), .B(KEYINPUT114), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1005), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n996), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1011), .A2(new_n1015), .A3(KEYINPUT118), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT120), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n525), .A2(G8), .A3(new_n529), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT119), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1018), .B(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n954), .A2(KEYINPUT45), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n953), .A2(new_n845), .B1(new_n495), .B2(new_n498), .ZN(new_n1022));
  AOI21_X1  g597(.A(G1384), .B1(new_n1022), .B2(new_n843), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n948), .B(new_n1021), .C1(new_n1023), .C2(KEYINPUT45), .ZN(new_n1024));
  INV_X1    g599(.A(G1966), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n1027));
  INV_X1    g602(.A(G2084), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n956), .A2(new_n1027), .A3(new_n1028), .A4(new_n957), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n966), .A2(new_n957), .A3(new_n1028), .A4(new_n948), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT112), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1026), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1020), .B1(new_n1032), .B2(G8), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1017), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n1024), .A2(new_n1025), .B1(new_n1030), .B2(KEYINPUT112), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n927), .B1(new_n1036), .B2(new_n1029), .ZN(new_n1037));
  OAI211_X1 g612(.A(KEYINPUT120), .B(KEYINPUT51), .C1(new_n1037), .C2(new_n1020), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1032), .A2(G8), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1039), .A2(new_n1034), .A3(new_n1018), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1035), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1032), .A2(G8), .A3(G286), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n945), .A2(new_n946), .A3(new_n767), .A4(new_n948), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g621(.A(KEYINPUT121), .B(G1961), .Z(new_n1047));
  NAND2_X1  g622(.A1(new_n967), .A2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1045), .A2(G2078), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n904), .A2(new_n948), .A3(new_n1021), .A4(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1046), .A2(new_n1048), .A3(G301), .A4(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT123), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1044), .A2(new_n1045), .B1(new_n967), .B2(new_n1047), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT123), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(G301), .A4(new_n1050), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n1057));
  INV_X1    g632(.A(new_n946), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n904), .A2(new_n948), .A3(new_n1049), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1046), .B(new_n1048), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1057), .B1(new_n1060), .B2(G171), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1056), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT124), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1056), .A2(KEYINPUT124), .A3(new_n1061), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(G301), .B1(new_n1053), .B2(new_n1050), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1067), .A2(KEYINPUT122), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1053), .A2(new_n1050), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1069), .A2(KEYINPUT122), .A3(G171), .ZN(new_n1070));
  OR2_X1    g645(.A1(new_n1060), .A2(G171), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n1057), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1043), .A2(new_n1066), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT118), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1016), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1043), .A2(KEYINPUT62), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n1043), .B2(KEYINPUT62), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n965), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(G288), .A2(G1976), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n929), .A2(new_n1082), .B1(new_n920), .B2(new_n680), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n929), .A2(new_n933), .A3(new_n935), .ZN(new_n1084));
  OAI22_X1  g659(.A1(new_n1083), .A2(new_n930), .B1(new_n963), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT113), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1039), .A2(G286), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1086), .B1(new_n964), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1084), .A2(new_n962), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1090), .A2(KEYINPUT113), .A3(new_n951), .A4(new_n1087), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT63), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1089), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1092), .B1(new_n940), .B2(new_n961), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1090), .A2(new_n1087), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1085), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n917), .B1(new_n1081), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n907), .A2(new_n976), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1098), .B(KEYINPUT46), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n909), .A2(new_n746), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n907), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT47), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n709), .A2(new_n712), .ZN(new_n1104));
  OAI22_X1  g679(.A1(new_n910), .A2(new_n1104), .B1(G2067), .B2(new_n787), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n907), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n907), .A2(new_n914), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT125), .B(KEYINPUT48), .ZN(new_n1108));
  OR2_X1    g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n912), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1103), .A2(new_n1106), .A3(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n900), .B1(new_n1097), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1112), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1085), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1066), .A2(new_n1073), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(new_n1121), .A3(new_n1043), .ZN(new_n1122));
  OAI22_X1  g697(.A1(new_n1122), .A2(new_n1016), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1117), .B1(new_n1123), .B2(new_n965), .ZN(new_n1124));
  OAI211_X1 g699(.A(KEYINPUT126), .B(new_n1114), .C1(new_n1124), .C2(new_n917), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1113), .A2(new_n1125), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g701(.A1(new_n894), .A2(new_n896), .ZN(new_n1128));
  NOR3_X1   g702(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1129));
  XOR2_X1   g703(.A(new_n1129), .B(KEYINPUT127), .Z(new_n1130));
  NOR2_X1   g704(.A1(new_n1130), .A2(G229), .ZN(new_n1131));
  NAND3_X1  g705(.A1(new_n1128), .A2(new_n1131), .A3(new_n856), .ZN(G225));
  INV_X1    g706(.A(G225), .ZN(G308));
endmodule


