

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740;

  XNOR2_X1 U371 ( .A(n410), .B(n443), .ZN(n364) );
  XNOR2_X1 U372 ( .A(n409), .B(G110), .ZN(n480) );
  XNOR2_X1 U373 ( .A(n411), .B(G113), .ZN(n410) );
  XNOR2_X1 U374 ( .A(n457), .B(n456), .ZN(n556) );
  AND2_X4 U375 ( .A1(n647), .A2(n646), .ZN(n704) );
  NAND2_X2 U376 ( .A1(n526), .A2(n618), .ZN(n528) );
  XNOR2_X2 U377 ( .A(n365), .B(n350), .ZN(n526) );
  XNOR2_X2 U378 ( .A(n719), .B(n491), .ZN(n673) );
  AND2_X2 U379 ( .A1(n582), .A2(n430), .ZN(n538) );
  XNOR2_X2 U380 ( .A(n486), .B(n431), .ZN(n726) );
  XNOR2_X2 U381 ( .A(n472), .B(KEYINPUT4), .ZN(n486) );
  AND2_X1 U382 ( .A1(n368), .A2(n366), .ZN(n398) );
  NOR2_X1 U383 ( .A1(n563), .A2(n348), .ZN(n367) );
  XNOR2_X1 U384 ( .A(n537), .B(KEYINPUT31), .ZN(n698) );
  XNOR2_X1 U385 ( .A(n442), .B(n441), .ZN(n508) );
  XNOR2_X1 U386 ( .A(n608), .B(n392), .ZN(n695) );
  XNOR2_X1 U387 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U388 ( .A(n726), .B(G146), .ZN(n450) );
  XNOR2_X1 U389 ( .A(n587), .B(KEYINPUT28), .ZN(n588) );
  XNOR2_X1 U390 ( .A(G134), .B(G131), .ZN(n431) );
  INV_X1 U391 ( .A(G119), .ZN(n409) );
  XNOR2_X1 U392 ( .A(KEYINPUT80), .B(KEYINPUT3), .ZN(n443) );
  INV_X1 U393 ( .A(G101), .ZN(n411) );
  XNOR2_X1 U394 ( .A(n397), .B(KEYINPUT96), .ZN(n396) );
  XNOR2_X2 U395 ( .A(n407), .B(n405), .ZN(n719) );
  XNOR2_X2 U396 ( .A(n545), .B(KEYINPUT22), .ZN(n551) );
  INV_X1 U397 ( .A(n594), .ZN(n402) );
  XNOR2_X1 U398 ( .A(n432), .B(G125), .ZN(n485) );
  XNOR2_X1 U399 ( .A(n599), .B(n598), .ZN(n617) );
  INV_X1 U400 ( .A(KEYINPUT102), .ZN(n598) );
  NAND2_X1 U401 ( .A1(n695), .A2(n390), .ZN(n599) );
  AND2_X1 U402 ( .A1(n597), .A2(n391), .ZN(n390) );
  XNOR2_X1 U403 ( .A(n495), .B(KEYINPUT92), .ZN(n608) );
  XNOR2_X1 U404 ( .A(n496), .B(KEYINPUT93), .ZN(n594) );
  AND2_X1 U405 ( .A1(n361), .A2(n387), .ZN(n615) );
  NOR2_X1 U406 ( .A1(n351), .A2(n700), .ZN(n361) );
  NOR2_X1 U407 ( .A1(n738), .A2(n737), .ZN(n388) );
  NAND2_X1 U408 ( .A1(n564), .A2(KEYINPUT64), .ZN(n395) );
  INV_X1 U409 ( .A(n583), .ZN(n577) );
  OR2_X1 U410 ( .A1(n668), .A2(G902), .ZN(n399) );
  OR2_X1 U411 ( .A1(n648), .A2(G902), .ZN(n452) );
  INV_X1 U412 ( .A(G140), .ZN(n421) );
  XNOR2_X1 U413 ( .A(G110), .B(G107), .ZN(n436) );
  XNOR2_X1 U414 ( .A(G104), .B(G101), .ZN(n437) );
  XNOR2_X1 U415 ( .A(n483), .B(KEYINPUT17), .ZN(n484) );
  INV_X1 U416 ( .A(KEYINPUT81), .ZN(n483) );
  AND2_X1 U417 ( .A1(G224), .A2(n733), .ZN(n488) );
  XNOR2_X1 U418 ( .A(n408), .B(n364), .ZN(n407) );
  XNOR2_X1 U419 ( .A(n480), .B(n481), .ZN(n408) );
  NOR2_X1 U420 ( .A1(n606), .A2(n605), .ZN(n607) );
  INV_X1 U421 ( .A(KEYINPUT78), .ZN(n527) );
  XNOR2_X1 U422 ( .A(n394), .B(n393), .ZN(n357) );
  INV_X1 U423 ( .A(KEYINPUT34), .ZN(n393) );
  XNOR2_X1 U424 ( .A(n385), .B(n383), .ZN(n558) );
  XNOR2_X1 U425 ( .A(n468), .B(n384), .ZN(n383) );
  INV_X1 U426 ( .A(G475), .ZN(n384) );
  BUF_X1 U427 ( .A(n602), .Z(n362) );
  INV_X2 U428 ( .A(G953), .ZN(n733) );
  INV_X1 U429 ( .A(KEYINPUT100), .ZN(n392) );
  OR2_X1 U430 ( .A1(n740), .A2(n657), .ZN(n563) );
  XNOR2_X1 U431 ( .A(G119), .B(G116), .ZN(n444) );
  XOR2_X1 U432 ( .A(G137), .B(KEYINPUT5), .Z(n445) );
  NOR2_X1 U433 ( .A1(n547), .A2(n658), .ZN(n397) );
  XNOR2_X1 U434 ( .A(n401), .B(n400), .ZN(n547) );
  INV_X1 U435 ( .A(KEYINPUT94), .ZN(n400) );
  XNOR2_X1 U436 ( .A(G902), .B(KEYINPUT15), .ZN(n641) );
  XNOR2_X1 U437 ( .A(G113), .B(G143), .ZN(n458) );
  XNOR2_X1 U438 ( .A(G131), .B(G140), .ZN(n459) );
  XOR2_X1 U439 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n460) );
  XNOR2_X1 U440 ( .A(n485), .B(n389), .ZN(n465) );
  INV_X1 U441 ( .A(KEYINPUT10), .ZN(n389) );
  INV_X1 U442 ( .A(G116), .ZN(n406) );
  INV_X1 U443 ( .A(n596), .ZN(n391) );
  XNOR2_X1 U444 ( .A(n550), .B(KEYINPUT98), .ZN(n586) );
  XNOR2_X1 U445 ( .A(n590), .B(KEYINPUT1), .ZN(n602) );
  XNOR2_X1 U446 ( .A(G134), .B(G122), .ZN(n469) );
  XNOR2_X1 U447 ( .A(KEYINPUT73), .B(KEYINPUT8), .ZN(n413) );
  NOR2_X1 U448 ( .A1(n732), .A2(n641), .ZN(n640) );
  NAND2_X1 U449 ( .A1(n380), .A2(n379), .ZN(n378) );
  INV_X1 U450 ( .A(KEYINPUT32), .ZN(n382) );
  NOR2_X1 U451 ( .A1(n349), .A2(n374), .ZN(n373) );
  OR2_X1 U452 ( .A1(n597), .A2(n382), .ZN(n374) );
  XNOR2_X1 U453 ( .A(n386), .B(n479), .ZN(n494) );
  XNOR2_X1 U454 ( .A(KEYINPUT91), .B(G478), .ZN(n479) );
  OR2_X1 U455 ( .A1(n705), .A2(G902), .ZN(n386) );
  NAND2_X1 U456 ( .A1(n356), .A2(n578), .ZN(n606) );
  AND2_X1 U457 ( .A1(n579), .A2(n577), .ZN(n356) );
  XNOR2_X1 U458 ( .A(n358), .B(KEYINPUT87), .ZN(n360) );
  INV_X1 U459 ( .A(n597), .ZN(n379) );
  INV_X1 U460 ( .A(n551), .ZN(n375) );
  XOR2_X1 U461 ( .A(n661), .B(KEYINPUT59), .Z(n662) );
  XNOR2_X1 U462 ( .A(n450), .B(n440), .ZN(n668) );
  XNOR2_X1 U463 ( .A(n488), .B(KEYINPUT18), .ZN(n489) );
  XNOR2_X1 U464 ( .A(n653), .B(KEYINPUT79), .ZN(n711) );
  NOR2_X1 U465 ( .A1(n603), .A2(n620), .ZN(n700) );
  AND2_X1 U466 ( .A1(n617), .A2(n600), .ZN(n601) );
  NAND2_X1 U467 ( .A1(n357), .A2(n559), .ZN(n561) );
  NAND2_X1 U468 ( .A1(n376), .A2(n372), .ZN(n740) );
  AND2_X1 U469 ( .A1(n381), .A2(n377), .ZN(n376) );
  NAND2_X1 U470 ( .A1(n375), .A2(n373), .ZN(n372) );
  NAND2_X1 U471 ( .A1(n378), .A2(n382), .ZN(n377) );
  INV_X1 U472 ( .A(n695), .ZN(n693) );
  AND2_X1 U473 ( .A1(KEYINPUT44), .A2(KEYINPUT64), .ZN(n348) );
  XOR2_X1 U474 ( .A(n549), .B(KEYINPUT97), .Z(n349) );
  AND2_X1 U475 ( .A1(G210), .A2(n492), .ZN(n350) );
  OR2_X1 U476 ( .A1(n604), .A2(n691), .ZN(n351) );
  INV_X1 U477 ( .A(G146), .ZN(n432) );
  XOR2_X1 U478 ( .A(n406), .B(G107), .Z(n352) );
  AND2_X1 U479 ( .A1(n370), .A2(n562), .ZN(n353) );
  AND2_X1 U480 ( .A1(n375), .A2(n379), .ZN(n354) );
  NOR2_X1 U481 ( .A1(n554), .A2(KEYINPUT64), .ZN(n355) );
  XNOR2_X1 U482 ( .A(n487), .B(n486), .ZN(n490) );
  INV_X1 U483 ( .A(n586), .ZN(n570) );
  XNOR2_X1 U484 ( .A(n388), .B(KEYINPUT46), .ZN(n387) );
  XNOR2_X2 U485 ( .A(n600), .B(KEYINPUT19), .ZN(n592) );
  NAND2_X1 U486 ( .A1(n555), .A2(n539), .ZN(n358) );
  NAND2_X1 U487 ( .A1(n359), .A2(n402), .ZN(n401) );
  NAND2_X1 U488 ( .A1(n404), .A2(n403), .ZN(n359) );
  NAND2_X1 U489 ( .A1(n360), .A2(n550), .ZN(n404) );
  XNOR2_X1 U490 ( .A(n589), .B(n588), .ZN(n591) );
  NAND2_X1 U491 ( .A1(n353), .A2(n369), .ZN(n368) );
  NAND2_X1 U492 ( .A1(n398), .A2(n396), .ZN(n565) );
  XNOR2_X2 U493 ( .A(n363), .B(n535), .ZN(n541) );
  NOR2_X2 U494 ( .A1(n592), .A2(n534), .ZN(n363) );
  XNOR2_X1 U495 ( .A(n364), .B(n448), .ZN(n449) );
  NAND2_X1 U496 ( .A1(n673), .A2(n641), .ZN(n365) );
  NAND2_X1 U497 ( .A1(n367), .A2(n395), .ZN(n366) );
  NAND2_X1 U498 ( .A1(n371), .A2(n660), .ZN(n369) );
  NAND2_X1 U499 ( .A1(n660), .A2(n355), .ZN(n370) );
  INV_X1 U500 ( .A(n563), .ZN(n371) );
  INV_X1 U501 ( .A(n349), .ZN(n380) );
  NAND2_X1 U502 ( .A1(n551), .A2(n382), .ZN(n381) );
  INV_X1 U503 ( .A(n494), .ZN(n557) );
  NAND2_X1 U504 ( .A1(n494), .A2(n558), .ZN(n495) );
  OR2_X1 U505 ( .A1(n661), .A2(G902), .ZN(n385) );
  XNOR2_X2 U506 ( .A(n528), .B(n527), .ZN(n600) );
  NAND2_X1 U507 ( .A1(n556), .A2(n555), .ZN(n394) );
  XNOR2_X2 U508 ( .A(G143), .B(G128), .ZN(n472) );
  XNOR2_X2 U509 ( .A(n399), .B(G469), .ZN(n590) );
  INV_X1 U510 ( .A(n404), .ZN(n680) );
  INV_X1 U511 ( .A(n698), .ZN(n403) );
  XNOR2_X1 U512 ( .A(n482), .B(n352), .ZN(n405) );
  XNOR2_X1 U513 ( .A(n485), .B(n484), .ZN(n487) );
  XNOR2_X1 U514 ( .A(n490), .B(n489), .ZN(n491) );
  INV_X1 U515 ( .A(KEYINPUT107), .ZN(n587) );
  XNOR2_X1 U516 ( .A(n541), .B(KEYINPUT83), .ZN(n555) );
  XNOR2_X1 U517 ( .A(n424), .B(KEYINPUT25), .ZN(n425) );
  NOR2_X1 U518 ( .A1(n611), .A2(n592), .ZN(n593) );
  INV_X1 U519 ( .A(n711), .ZN(n654) );
  XNOR2_X1 U520 ( .A(n607), .B(KEYINPUT39), .ZN(n616) );
  XNOR2_X1 U521 ( .A(n639), .B(n638), .ZN(G75) );
  NAND2_X1 U522 ( .A1(G234), .A2(G237), .ZN(n412) );
  XNOR2_X1 U523 ( .A(KEYINPUT14), .B(n412), .ZN(n532) );
  NAND2_X1 U524 ( .A1(G952), .A2(n532), .ZN(n529) );
  XOR2_X1 U525 ( .A(n480), .B(KEYINPUT24), .Z(n416) );
  NAND2_X1 U526 ( .A1(n733), .A2(G234), .ZN(n414) );
  XNOR2_X1 U527 ( .A(n414), .B(n413), .ZN(n476) );
  NAND2_X1 U528 ( .A1(G221), .A2(n476), .ZN(n415) );
  XNOR2_X1 U529 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U530 ( .A(KEYINPUT23), .B(KEYINPUT84), .Z(n418) );
  XNOR2_X1 U531 ( .A(G128), .B(KEYINPUT85), .ZN(n417) );
  XNOR2_X1 U532 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U533 ( .A(n420), .B(n419), .ZN(n422) );
  XNOR2_X1 U534 ( .A(n421), .B(G137), .ZN(n435) );
  XOR2_X1 U535 ( .A(n435), .B(n465), .Z(n725) );
  XNOR2_X1 U536 ( .A(n422), .B(n725), .ZN(n708) );
  NOR2_X1 U537 ( .A1(G902), .A2(n708), .ZN(n426) );
  NAND2_X1 U538 ( .A1(G234), .A2(n641), .ZN(n423) );
  XNOR2_X1 U539 ( .A(KEYINPUT20), .B(n423), .ZN(n427) );
  NAND2_X1 U540 ( .A1(n427), .A2(G217), .ZN(n424) );
  XNOR2_X2 U541 ( .A(n426), .B(n425), .ZN(n582) );
  NAND2_X1 U542 ( .A1(n427), .A2(G221), .ZN(n428) );
  XOR2_X1 U543 ( .A(n428), .B(KEYINPUT21), .Z(n584) );
  INV_X1 U544 ( .A(KEYINPUT86), .ZN(n429) );
  XNOR2_X1 U545 ( .A(n584), .B(n429), .ZN(n542) );
  INV_X1 U546 ( .A(n542), .ZN(n430) );
  NAND2_X1 U547 ( .A1(n733), .A2(G227), .ZN(n433) );
  XNOR2_X1 U548 ( .A(n433), .B(KEYINPUT70), .ZN(n434) );
  XNOR2_X1 U549 ( .A(n435), .B(n434), .ZN(n439) );
  XNOR2_X1 U550 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U551 ( .A(n439), .B(n438), .ZN(n440) );
  NAND2_X1 U552 ( .A1(n538), .A2(n602), .ZN(n442) );
  INV_X1 U553 ( .A(KEYINPUT69), .ZN(n441) );
  XNOR2_X1 U554 ( .A(n508), .B(KEYINPUT99), .ZN(n455) );
  XNOR2_X1 U555 ( .A(n445), .B(n444), .ZN(n447) );
  NOR2_X1 U556 ( .A1(G953), .A2(G237), .ZN(n463) );
  NAND2_X1 U557 ( .A1(n463), .A2(G210), .ZN(n446) );
  XNOR2_X1 U558 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U559 ( .A(n450), .B(n449), .ZN(n648) );
  XNOR2_X1 U560 ( .A(G472), .B(KEYINPUT67), .ZN(n451) );
  XNOR2_X2 U561 ( .A(n452), .B(n451), .ZN(n550) );
  INV_X1 U562 ( .A(KEYINPUT95), .ZN(n453) );
  XNOR2_X1 U563 ( .A(n453), .B(KEYINPUT6), .ZN(n454) );
  XNOR2_X1 U564 ( .A(n550), .B(n454), .ZN(n597) );
  NAND2_X1 U565 ( .A1(n455), .A2(n597), .ZN(n457) );
  XNOR2_X1 U566 ( .A(KEYINPUT66), .B(KEYINPUT33), .ZN(n456) );
  INV_X1 U567 ( .A(n556), .ZN(n523) );
  XOR2_X1 U568 ( .A(G122), .B(G104), .Z(n482) );
  XNOR2_X1 U569 ( .A(n458), .B(n482), .ZN(n462) );
  XNOR2_X1 U570 ( .A(n460), .B(n459), .ZN(n461) );
  XOR2_X1 U571 ( .A(n462), .B(n461), .Z(n467) );
  NAND2_X1 U572 ( .A1(G214), .A2(n463), .ZN(n464) );
  XNOR2_X1 U573 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U574 ( .A(n467), .B(n466), .ZN(n661) );
  XNOR2_X1 U575 ( .A(KEYINPUT88), .B(KEYINPUT13), .ZN(n468) );
  XOR2_X1 U576 ( .A(KEYINPUT90), .B(KEYINPUT9), .Z(n470) );
  XNOR2_X1 U577 ( .A(n470), .B(n469), .ZN(n475) );
  XOR2_X1 U578 ( .A(KEYINPUT89), .B(KEYINPUT7), .Z(n471) );
  XNOR2_X1 U579 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U580 ( .A(n473), .B(n352), .ZN(n474) );
  XOR2_X1 U581 ( .A(n475), .B(n474), .Z(n478) );
  NAND2_X1 U582 ( .A1(G217), .A2(n476), .ZN(n477) );
  XNOR2_X1 U583 ( .A(n478), .B(n477), .ZN(n705) );
  NOR2_X1 U584 ( .A1(n558), .A2(n557), .ZN(n544) );
  INV_X1 U585 ( .A(n544), .ZN(n513) );
  XNOR2_X1 U586 ( .A(KEYINPUT16), .B(KEYINPUT68), .ZN(n481) );
  OR2_X1 U587 ( .A1(G237), .A2(G902), .ZN(n492) );
  INV_X1 U588 ( .A(n526), .ZN(n624) );
  XOR2_X1 U589 ( .A(n624), .B(KEYINPUT38), .Z(n605) );
  INV_X1 U590 ( .A(n605), .ZN(n497) );
  NAND2_X1 U591 ( .A1(G214), .A2(n492), .ZN(n618) );
  NOR2_X1 U592 ( .A1(n497), .A2(n618), .ZN(n493) );
  NOR2_X1 U593 ( .A1(n513), .A2(n493), .ZN(n499) );
  NOR2_X1 U594 ( .A1(n494), .A2(n558), .ZN(n697) );
  INV_X1 U595 ( .A(n697), .ZN(n687) );
  NAND2_X1 U596 ( .A1(n687), .A2(n608), .ZN(n496) );
  NAND2_X1 U597 ( .A1(n497), .A2(n618), .ZN(n512) );
  NOR2_X1 U598 ( .A1(n594), .A2(n512), .ZN(n498) );
  NOR2_X1 U599 ( .A1(n499), .A2(n498), .ZN(n500) );
  NOR2_X1 U600 ( .A1(n523), .A2(n500), .ZN(n501) );
  XNOR2_X1 U601 ( .A(n501), .B(KEYINPUT115), .ZN(n519) );
  INV_X1 U602 ( .A(n550), .ZN(n540) );
  NOR2_X1 U603 ( .A1(n584), .A2(n582), .ZN(n502) );
  XOR2_X1 U604 ( .A(KEYINPUT49), .B(n502), .Z(n503) );
  NOR2_X1 U605 ( .A1(n540), .A2(n503), .ZN(n504) );
  XOR2_X1 U606 ( .A(KEYINPUT114), .B(n504), .Z(n507) );
  NOR2_X1 U607 ( .A1(n538), .A2(n362), .ZN(n505) );
  XNOR2_X1 U608 ( .A(n505), .B(KEYINPUT50), .ZN(n506) );
  NOR2_X1 U609 ( .A1(n507), .A2(n506), .ZN(n510) );
  OR2_X1 U610 ( .A1(n508), .A2(n550), .ZN(n536) );
  INV_X1 U611 ( .A(n536), .ZN(n509) );
  NOR2_X1 U612 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U613 ( .A(KEYINPUT51), .B(n511), .ZN(n517) );
  NOR2_X1 U614 ( .A1(n513), .A2(n512), .ZN(n515) );
  XNOR2_X1 U615 ( .A(KEYINPUT41), .B(KEYINPUT109), .ZN(n514) );
  XOR2_X1 U616 ( .A(n515), .B(n514), .Z(n612) );
  INV_X1 U617 ( .A(n612), .ZN(n516) );
  NAND2_X1 U618 ( .A1(n517), .A2(n516), .ZN(n518) );
  NAND2_X1 U619 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U620 ( .A(n520), .B(KEYINPUT116), .ZN(n521) );
  XOR2_X1 U621 ( .A(KEYINPUT52), .B(n521), .Z(n522) );
  NOR2_X1 U622 ( .A1(n529), .A2(n522), .ZN(n525) );
  NOR2_X1 U623 ( .A1(n523), .A2(n612), .ZN(n524) );
  NOR2_X1 U624 ( .A1(n525), .A2(n524), .ZN(n637) );
  NOR2_X1 U625 ( .A1(n529), .A2(G953), .ZN(n530) );
  XNOR2_X1 U626 ( .A(n530), .B(KEYINPUT82), .ZN(n575) );
  AND2_X1 U627 ( .A1(G953), .A2(G902), .ZN(n531) );
  NAND2_X1 U628 ( .A1(n532), .A2(n531), .ZN(n573) );
  NOR2_X1 U629 ( .A1(n573), .A2(G898), .ZN(n533) );
  NOR2_X1 U630 ( .A1(n575), .A2(n533), .ZN(n534) );
  INV_X1 U631 ( .A(KEYINPUT0), .ZN(n535) );
  OR2_X1 U632 ( .A1(n541), .A2(n536), .ZN(n537) );
  NAND2_X1 U633 ( .A1(n538), .A2(n590), .ZN(n569) );
  INV_X1 U634 ( .A(n569), .ZN(n539) );
  NOR2_X1 U635 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U636 ( .A1(n544), .A2(n543), .ZN(n545) );
  INV_X1 U637 ( .A(n582), .ZN(n548) );
  NOR2_X1 U638 ( .A1(n548), .A2(n362), .ZN(n546) );
  AND2_X1 U639 ( .A1(n354), .A2(n546), .ZN(n658) );
  NAND2_X1 U640 ( .A1(n548), .A2(n362), .ZN(n549) );
  NOR2_X1 U641 ( .A1(n551), .A2(n570), .ZN(n553) );
  NOR2_X1 U642 ( .A1(n362), .A2(n582), .ZN(n552) );
  AND2_X1 U643 ( .A1(n553), .A2(n552), .ZN(n657) );
  INV_X1 U644 ( .A(KEYINPUT44), .ZN(n554) );
  NAND2_X1 U645 ( .A1(n558), .A2(n557), .ZN(n580) );
  INV_X1 U646 ( .A(n580), .ZN(n559) );
  XNOR2_X1 U647 ( .A(KEYINPUT77), .B(KEYINPUT35), .ZN(n560) );
  XNOR2_X2 U648 ( .A(n561), .B(n560), .ZN(n660) );
  NAND2_X1 U649 ( .A1(n554), .A2(KEYINPUT64), .ZN(n562) );
  INV_X1 U650 ( .A(n660), .ZN(n564) );
  XNOR2_X2 U651 ( .A(n565), .B(KEYINPUT45), .ZN(n712) );
  INV_X1 U652 ( .A(n712), .ZN(n566) );
  INV_X1 U653 ( .A(KEYINPUT2), .ZN(n630) );
  NAND2_X1 U654 ( .A1(n566), .A2(n630), .ZN(n568) );
  INV_X1 U655 ( .A(KEYINPUT74), .ZN(n567) );
  XNOR2_X1 U656 ( .A(n568), .B(n567), .ZN(n634) );
  XNOR2_X1 U657 ( .A(n569), .B(KEYINPUT105), .ZN(n579) );
  NAND2_X1 U658 ( .A1(n570), .A2(n618), .ZN(n572) );
  XOR2_X1 U659 ( .A(KEYINPUT30), .B(KEYINPUT106), .Z(n571) );
  XNOR2_X1 U660 ( .A(n572), .B(n571), .ZN(n578) );
  XOR2_X1 U661 ( .A(KEYINPUT101), .B(n573), .Z(n574) );
  NOR2_X1 U662 ( .A1(G900), .A2(n574), .ZN(n576) );
  NOR2_X1 U663 ( .A1(n576), .A2(n575), .ZN(n583) );
  OR2_X1 U664 ( .A1(n624), .A2(n580), .ZN(n581) );
  NOR2_X1 U665 ( .A1(n606), .A2(n581), .ZN(n691) );
  NOR2_X1 U666 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U667 ( .A1(n585), .A2(n584), .ZN(n596) );
  NOR2_X1 U668 ( .A1(n586), .A2(n596), .ZN(n589) );
  NAND2_X1 U669 ( .A1(n591), .A2(n590), .ZN(n611) );
  XNOR2_X1 U670 ( .A(n593), .B(KEYINPUT71), .ZN(n692) );
  NOR2_X1 U671 ( .A1(n692), .A2(n594), .ZN(n595) );
  XOR2_X1 U672 ( .A(KEYINPUT47), .B(n595), .Z(n604) );
  XOR2_X1 U673 ( .A(KEYINPUT36), .B(n601), .Z(n603) );
  INV_X1 U674 ( .A(n362), .ZN(n620) );
  NOR2_X1 U675 ( .A1(n608), .A2(n616), .ZN(n610) );
  XNOR2_X1 U676 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n609) );
  XNOR2_X1 U677 ( .A(n610), .B(n609), .ZN(n738) );
  OR2_X1 U678 ( .A1(n612), .A2(n611), .ZN(n614) );
  XOR2_X1 U679 ( .A(KEYINPUT42), .B(KEYINPUT110), .Z(n613) );
  XNOR2_X1 U680 ( .A(n614), .B(n613), .ZN(n737) );
  XNOR2_X1 U681 ( .A(KEYINPUT48), .B(n615), .ZN(n628) );
  NOR2_X1 U682 ( .A1(n616), .A2(n687), .ZN(n702) );
  INV_X1 U683 ( .A(n702), .ZN(n626) );
  NAND2_X1 U684 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U685 ( .A(KEYINPUT103), .B(n619), .ZN(n621) );
  NAND2_X1 U686 ( .A1(n621), .A2(n620), .ZN(n623) );
  XNOR2_X1 U687 ( .A(KEYINPUT104), .B(KEYINPUT43), .ZN(n622) );
  XNOR2_X1 U688 ( .A(n623), .B(n622), .ZN(n625) );
  NAND2_X1 U689 ( .A1(n625), .A2(n624), .ZN(n703) );
  AND2_X1 U690 ( .A1(n626), .A2(n703), .ZN(n627) );
  NAND2_X1 U691 ( .A1(n628), .A2(n627), .ZN(n732) );
  NOR2_X1 U692 ( .A1(n732), .A2(n630), .ZN(n629) );
  NAND2_X1 U693 ( .A1(n712), .A2(n629), .ZN(n646) );
  AND2_X1 U694 ( .A1(n630), .A2(n732), .ZN(n631) );
  XNOR2_X1 U695 ( .A(n631), .B(KEYINPUT75), .ZN(n632) );
  NAND2_X1 U696 ( .A1(n646), .A2(n632), .ZN(n633) );
  NOR2_X1 U697 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U698 ( .A1(G953), .A2(n635), .ZN(n636) );
  NAND2_X1 U699 ( .A1(n637), .A2(n636), .ZN(n639) );
  XNOR2_X1 U700 ( .A(KEYINPUT53), .B(KEYINPUT117), .ZN(n638) );
  NAND2_X1 U701 ( .A1(n712), .A2(n640), .ZN(n645) );
  XOR2_X1 U702 ( .A(KEYINPUT76), .B(n641), .Z(n642) );
  NAND2_X1 U703 ( .A1(n642), .A2(KEYINPUT2), .ZN(n643) );
  XOR2_X1 U704 ( .A(KEYINPUT65), .B(n643), .Z(n644) );
  NAND2_X1 U705 ( .A1(n645), .A2(n644), .ZN(n647) );
  NAND2_X1 U706 ( .A1(n704), .A2(G472), .ZN(n650) );
  XNOR2_X1 U707 ( .A(n648), .B(KEYINPUT62), .ZN(n649) );
  XNOR2_X1 U708 ( .A(n650), .B(n649), .ZN(n651) );
  INV_X1 U709 ( .A(n651), .ZN(n655) );
  INV_X1 U710 ( .A(G952), .ZN(n652) );
  NAND2_X1 U711 ( .A1(n652), .A2(G953), .ZN(n653) );
  NAND2_X1 U712 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U713 ( .A(n656), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U714 ( .A(G110), .B(n657), .Z(G12) );
  XOR2_X1 U715 ( .A(G101), .B(n658), .Z(G3) );
  XNOR2_X1 U716 ( .A(G122), .B(KEYINPUT126), .ZN(n659) );
  XNOR2_X1 U717 ( .A(n660), .B(n659), .ZN(G24) );
  NAND2_X1 U718 ( .A1(n704), .A2(G475), .ZN(n663) );
  XNOR2_X1 U719 ( .A(n663), .B(n662), .ZN(n664) );
  NOR2_X2 U720 ( .A1(n664), .A2(n711), .ZN(n666) );
  XOR2_X1 U721 ( .A(KEYINPUT119), .B(KEYINPUT60), .Z(n665) );
  XNOR2_X1 U722 ( .A(n666), .B(n665), .ZN(G60) );
  NAND2_X1 U723 ( .A1(n704), .A2(G469), .ZN(n670) );
  XOR2_X1 U724 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n667) );
  XNOR2_X1 U725 ( .A(n670), .B(n669), .ZN(n671) );
  NOR2_X2 U726 ( .A1(n671), .A2(n711), .ZN(n672) );
  XNOR2_X1 U727 ( .A(n672), .B(KEYINPUT118), .ZN(G54) );
  NAND2_X1 U728 ( .A1(n704), .A2(G210), .ZN(n677) );
  XNOR2_X1 U729 ( .A(KEYINPUT72), .B(KEYINPUT54), .ZN(n674) );
  XNOR2_X1 U730 ( .A(n674), .B(KEYINPUT55), .ZN(n675) );
  XNOR2_X1 U731 ( .A(n673), .B(n675), .ZN(n676) );
  XNOR2_X1 U732 ( .A(n677), .B(n676), .ZN(n678) );
  NOR2_X2 U733 ( .A1(n678), .A2(n711), .ZN(n679) );
  XNOR2_X1 U734 ( .A(n679), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U735 ( .A(G104), .B(KEYINPUT111), .Z(n682) );
  NAND2_X1 U736 ( .A1(n680), .A2(n695), .ZN(n681) );
  XNOR2_X1 U737 ( .A(n682), .B(n681), .ZN(G6) );
  XNOR2_X1 U738 ( .A(KEYINPUT26), .B(KEYINPUT112), .ZN(n686) );
  XOR2_X1 U739 ( .A(G107), .B(KEYINPUT27), .Z(n684) );
  NAND2_X1 U740 ( .A1(n680), .A2(n697), .ZN(n683) );
  XNOR2_X1 U741 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U742 ( .A(n686), .B(n685), .ZN(G9) );
  NOR2_X1 U743 ( .A1(n687), .A2(n692), .ZN(n689) );
  XNOR2_X1 U744 ( .A(KEYINPUT113), .B(KEYINPUT29), .ZN(n688) );
  XNOR2_X1 U745 ( .A(n689), .B(n688), .ZN(n690) );
  XOR2_X1 U746 ( .A(G128), .B(n690), .Z(G30) );
  XOR2_X1 U747 ( .A(G143), .B(n691), .Z(G45) );
  NOR2_X1 U748 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U749 ( .A(G146), .B(n694), .Z(G48) );
  NAND2_X1 U750 ( .A1(n698), .A2(n695), .ZN(n696) );
  XNOR2_X1 U751 ( .A(n696), .B(G113), .ZN(G15) );
  NAND2_X1 U752 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U753 ( .A(n699), .B(G116), .ZN(G18) );
  XNOR2_X1 U754 ( .A(n700), .B(G125), .ZN(n701) );
  XNOR2_X1 U755 ( .A(n701), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U756 ( .A(G134), .B(n702), .Z(G36) );
  XNOR2_X1 U757 ( .A(G140), .B(n703), .ZN(G42) );
  NAND2_X1 U758 ( .A1(n704), .A2(G478), .ZN(n706) );
  XNOR2_X1 U759 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U760 ( .A1(n711), .A2(n707), .ZN(G63) );
  NAND2_X1 U761 ( .A1(n704), .A2(G217), .ZN(n709) );
  XNOR2_X1 U762 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U763 ( .A1(n711), .A2(n710), .ZN(G66) );
  NAND2_X1 U764 ( .A1(n712), .A2(n733), .ZN(n713) );
  XOR2_X1 U765 ( .A(KEYINPUT121), .B(n713), .Z(n718) );
  NAND2_X1 U766 ( .A1(G224), .A2(G953), .ZN(n714) );
  XNOR2_X1 U767 ( .A(n714), .B(KEYINPUT120), .ZN(n715) );
  XNOR2_X1 U768 ( .A(KEYINPUT61), .B(n715), .ZN(n716) );
  NAND2_X1 U769 ( .A1(n716), .A2(G898), .ZN(n717) );
  NAND2_X1 U770 ( .A1(n718), .A2(n717), .ZN(n723) );
  XNOR2_X1 U771 ( .A(KEYINPUT123), .B(n719), .ZN(n721) );
  NOR2_X1 U772 ( .A1(n733), .A2(G898), .ZN(n720) );
  NOR2_X1 U773 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U774 ( .A(n723), .B(n722), .ZN(n724) );
  XNOR2_X1 U775 ( .A(KEYINPUT122), .B(n724), .ZN(G69) );
  XOR2_X1 U776 ( .A(n725), .B(KEYINPUT124), .Z(n727) );
  XNOR2_X1 U777 ( .A(n726), .B(n727), .ZN(n731) );
  XOR2_X1 U778 ( .A(n731), .B(KEYINPUT125), .Z(n728) );
  XNOR2_X1 U779 ( .A(G227), .B(n728), .ZN(n729) );
  NAND2_X1 U780 ( .A1(G900), .A2(n729), .ZN(n730) );
  NAND2_X1 U781 ( .A1(n730), .A2(G953), .ZN(n736) );
  XNOR2_X1 U782 ( .A(n732), .B(n731), .ZN(n734) );
  NAND2_X1 U783 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U784 ( .A1(n736), .A2(n735), .ZN(G72) );
  XOR2_X1 U785 ( .A(G137), .B(n737), .Z(G39) );
  XNOR2_X1 U786 ( .A(n738), .B(G131), .ZN(n739) );
  XNOR2_X1 U787 ( .A(n739), .B(KEYINPUT127), .ZN(G33) );
  XOR2_X1 U788 ( .A(G119), .B(n740), .Z(G21) );
endmodule

