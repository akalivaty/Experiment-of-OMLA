//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G122), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT93), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT68), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G116), .ZN(new_n192));
  INV_X1    g006(.A(G116), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT68), .A3(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n193), .A2(G119), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G113), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT2), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G113), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(KEYINPUT69), .B1(new_n198), .B2(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n196), .B1(new_n192), .B2(new_n194), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT69), .ZN(new_n207));
  NOR3_X1   g021(.A1(new_n206), .A2(new_n207), .A3(new_n203), .ZN(new_n208));
  AND4_X1   g022(.A1(KEYINPUT70), .A2(new_n195), .A3(new_n197), .A4(new_n203), .ZN(new_n209));
  AOI21_X1  g023(.A(KEYINPUT70), .B1(new_n206), .B2(new_n203), .ZN(new_n210));
  OAI22_X1  g024(.A1(new_n205), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(KEYINPUT87), .A2(G107), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G104), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(KEYINPUT3), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT87), .A2(G107), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G107), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT88), .B1(new_n218), .B2(G104), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT88), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(new_n214), .A3(G107), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(G104), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT3), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n217), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G101), .ZN(new_n226));
  AND2_X1   g040(.A1(KEYINPUT87), .A2(G107), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(new_n212), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n228), .A2(new_n215), .B1(KEYINPUT3), .B2(new_n223), .ZN(new_n229));
  AOI21_X1  g043(.A(G101), .B1(new_n219), .B2(new_n221), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n226), .A2(new_n231), .A3(KEYINPUT4), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT4), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n225), .A2(new_n233), .A3(G101), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n211), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(new_n198), .B2(new_n204), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n206), .A2(KEYINPUT70), .A3(new_n203), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n223), .B1(new_n228), .B2(G104), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n229), .A2(new_n230), .B1(new_n240), .B2(G101), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n206), .A2(KEYINPUT5), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n242), .B(G113), .C1(KEYINPUT5), .C2(new_n197), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n239), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  AOI211_X1 g058(.A(KEYINPUT6), .B(new_n189), .C1(new_n235), .C2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G146), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G143), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT1), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G128), .ZN(new_n249));
  INV_X1    g063(.A(G143), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT64), .B1(new_n246), .B2(G143), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(new_n250), .A3(G146), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(KEYINPUT1), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n257), .A2(new_n247), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT66), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n250), .A2(G146), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n262), .B1(new_n254), .B2(new_n256), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT66), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(new_n259), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n253), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G125), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G224), .ZN(new_n270));
  AND2_X1   g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  NOR2_X1   g085(.A1(KEYINPUT0), .A2(G128), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n263), .A2(new_n271), .B1(new_n273), .B2(new_n252), .ZN(new_n274));
  OR2_X1    g088(.A1(new_n274), .A2(new_n267), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n268), .A2(new_n270), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n270), .B1(new_n268), .B2(new_n275), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n232), .A2(new_n234), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n198), .A2(KEYINPUT69), .A3(new_n204), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n207), .B1(new_n206), .B2(new_n203), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n237), .A2(new_n238), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n244), .B(new_n189), .C1(new_n279), .C2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT94), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n235), .A2(KEYINPUT94), .A3(new_n244), .A4(new_n189), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT6), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n235), .A2(new_n244), .ZN(new_n289));
  INV_X1    g103(.A(new_n189), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI211_X1 g105(.A(new_n245), .B(new_n278), .C1(new_n287), .C2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n285), .A2(new_n286), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n268), .A2(new_n275), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT7), .ZN(new_n296));
  INV_X1    g110(.A(new_n270), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n268), .A2(KEYINPUT7), .A3(new_n270), .A4(new_n275), .ZN(new_n299));
  INV_X1    g113(.A(new_n244), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n241), .B1(new_n239), .B2(new_n243), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XOR2_X1   g116(.A(new_n189), .B(KEYINPUT8), .Z(new_n303));
  OAI211_X1 g117(.A(new_n298), .B(new_n299), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n293), .B1(new_n294), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G210), .B1(G237), .B2(G902), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NOR3_X1   g121(.A1(new_n292), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n287), .A2(new_n291), .ZN(new_n309));
  INV_X1    g123(.A(new_n278), .ZN(new_n310));
  INV_X1    g124(.A(new_n245), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n301), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n303), .B1(new_n313), .B2(new_n244), .ZN(new_n314));
  INV_X1    g128(.A(new_n299), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n268), .A2(new_n275), .B1(KEYINPUT7), .B2(new_n270), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(G902), .B1(new_n317), .B2(new_n287), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n306), .B1(new_n312), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n187), .B1(new_n308), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT95), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G952), .ZN(new_n323));
  AOI211_X1 g137(.A(G953), .B(new_n323), .C1(G234), .C2(G237), .ZN(new_n324));
  XOR2_X1   g138(.A(KEYINPUT78), .B(G902), .Z(new_n325));
  AOI211_X1 g139(.A(new_n269), .B(new_n325), .C1(G234), .C2(G237), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT21), .B(G898), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n187), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n307), .B1(new_n292), .B2(new_n305), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n312), .A2(new_n318), .A3(new_n306), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT95), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n322), .A2(new_n329), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G469), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n269), .A2(G227), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(KEYINPUT86), .ZN(new_n338));
  XNOR2_X1  g152(.A(G110), .B(G140), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n338), .B(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n217), .A2(new_n224), .ZN(new_n341));
  INV_X1    g155(.A(G101), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n222), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT4), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n342), .B1(new_n229), .B2(new_n222), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n274), .B(new_n234), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT89), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n232), .A2(KEYINPUT89), .A3(new_n274), .A4(new_n234), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT11), .ZN(new_n351));
  INV_X1    g165(.A(G134), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n351), .B1(new_n352), .B2(G137), .ZN(new_n353));
  INV_X1    g167(.A(G137), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(KEYINPUT11), .A3(G134), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(G137), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n353), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G131), .ZN(new_n358));
  INV_X1    g172(.A(G131), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n353), .A2(new_n355), .A3(new_n359), .A4(new_n356), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n240), .A2(G101), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n231), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT10), .B1(new_n266), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n263), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT90), .ZN(new_n367));
  OAI21_X1  g181(.A(G128), .B1(new_n248), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(KEYINPUT90), .B1(new_n247), .B2(KEYINPUT1), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AND4_X1   g184(.A1(new_n264), .A2(new_n257), .A3(new_n247), .A4(new_n259), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n264), .B1(new_n263), .B2(new_n259), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(new_n241), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n365), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n350), .A2(new_n362), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT91), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n348), .A2(new_n349), .B1(new_n365), .B2(new_n375), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT91), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(new_n362), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n350), .A2(new_n376), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT92), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT92), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n379), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n361), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n340), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n340), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n249), .A2(new_n252), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n390), .B1(new_n371), .B2(new_n372), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(new_n241), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n261), .A2(new_n265), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n364), .B1(new_n393), .B2(new_n370), .ZN(new_n394));
  OAI211_X1 g208(.A(KEYINPUT12), .B(new_n361), .C1(new_n392), .C2(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n361), .B1(new_n392), .B2(new_n394), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT12), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI221_X4 g212(.A(new_n389), .B1(new_n395), .B2(new_n398), .C1(new_n378), .C2(new_n381), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n336), .B(new_n325), .C1(new_n388), .C2(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n336), .A2(new_n293), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n398), .A2(new_n395), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n382), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n389), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n389), .B1(new_n378), .B2(new_n381), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n387), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(G469), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n400), .A2(new_n402), .A3(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT9), .B(G234), .ZN(new_n410));
  OAI21_X1  g224(.A(G221), .B1(new_n410), .B2(G902), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT85), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n193), .A2(G122), .ZN(new_n414));
  INV_X1    g228(.A(G122), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(G116), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n417), .B(new_n228), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n250), .A2(G128), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT13), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n258), .A2(G143), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n419), .A2(new_n420), .ZN(new_n424));
  OAI21_X1  g238(.A(G134), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n419), .A2(new_n422), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n352), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n418), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n426), .B(new_n352), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n417), .A2(new_n228), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n193), .A2(G122), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT14), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(KEYINPUT100), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT14), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n414), .B1(new_n435), .B2(new_n416), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n218), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n428), .B1(new_n431), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G217), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n410), .A2(new_n439), .A3(G953), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n428), .B(new_n440), .C1(new_n431), .C2(new_n437), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n325), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT15), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n446), .A3(G478), .ZN(new_n447));
  INV_X1    g261(.A(G478), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n444), .B(new_n325), .C1(KEYINPUT15), .C2(new_n448), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(G237), .A2(G953), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G214), .ZN(new_n452));
  NOR2_X1   g266(.A1(KEYINPUT96), .A2(G143), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n451), .B(G214), .C1(KEYINPUT96), .C2(G143), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(KEYINPUT18), .A3(G131), .ZN(new_n457));
  XNOR2_X1  g271(.A(G125), .B(G140), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(new_n246), .ZN(new_n459));
  NAND2_X1  g273(.A1(KEYINPUT18), .A2(G131), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n454), .A2(new_n460), .A3(new_n455), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n457), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n456), .A2(G131), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n454), .A2(new_n359), .A3(new_n455), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n458), .B(KEYINPUT19), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n465), .B1(new_n467), .B2(G146), .ZN(new_n468));
  INV_X1    g282(.A(G140), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G125), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n267), .A2(G140), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT16), .ZN(new_n472));
  OR3_X1    g286(.A1(new_n267), .A2(KEYINPUT16), .A3(G140), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT82), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(new_n475), .A3(G146), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n472), .A2(new_n473), .A3(G146), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT82), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n462), .B1(new_n468), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G113), .B(G122), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(new_n214), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT17), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n463), .A2(new_n485), .A3(new_n464), .ZN(new_n486));
  AOI21_X1  g300(.A(G146), .B1(new_n472), .B2(new_n473), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT80), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n487), .B1(new_n488), .B2(new_n477), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n474), .A2(KEYINPUT80), .A3(G146), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n456), .A2(KEYINPUT17), .A3(G131), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n486), .A2(new_n489), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n482), .A3(new_n462), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n484), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(G475), .A2(G902), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT97), .B1(new_n484), .B2(new_n493), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n496), .B1(KEYINPUT20), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT20), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n494), .A2(KEYINPUT97), .A3(new_n499), .A4(new_n495), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n492), .A2(new_n462), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n483), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n493), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n293), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT99), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT99), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n504), .A2(new_n507), .A3(new_n293), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT98), .B(G475), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n501), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n409), .A2(new_n413), .A3(new_n450), .A4(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n335), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(G472), .A2(G902), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n514), .A2(KEYINPUT32), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT76), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT71), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n211), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n361), .A2(new_n274), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n352), .A2(G137), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n354), .A2(G134), .ZN(new_n521));
  OAI21_X1  g335(.A(G131), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n360), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n391), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n280), .A2(new_n281), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n239), .A2(KEYINPUT71), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n518), .A2(new_n519), .A3(new_n525), .A4(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT72), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT65), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n523), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n360), .A2(new_n522), .A3(KEYINPUT65), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT67), .B1(new_n266), .B2(new_n534), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n360), .A2(new_n522), .A3(KEYINPUT65), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT65), .B1(new_n360), .B2(new_n522), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT67), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n391), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n535), .A2(new_n540), .A3(new_n519), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n211), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n391), .A2(new_n524), .B1(new_n361), .B2(new_n274), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n543), .A2(KEYINPUT72), .A3(new_n518), .A4(new_n527), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n530), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT28), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT28), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n528), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(KEYINPUT74), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n451), .A2(G210), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT26), .B(G101), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n553), .B(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n516), .B1(new_n549), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n548), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n559), .B1(new_n545), .B2(KEYINPUT28), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n560), .A2(KEYINPUT76), .A3(new_n556), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n530), .A2(new_n544), .A3(new_n556), .ZN(new_n563));
  OAI211_X1 g377(.A(KEYINPUT30), .B(new_n519), .C1(new_n266), .C2(new_n523), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n211), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT30), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n565), .B1(new_n566), .B2(new_n541), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT31), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n563), .A2(KEYINPUT31), .A3(new_n567), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT75), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n530), .A2(new_n544), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n541), .A2(new_n566), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(new_n211), .A3(new_n564), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(new_n556), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(KEYINPUT75), .A3(KEYINPUT31), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n515), .B1(new_n562), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n572), .A2(new_n574), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT29), .B1(new_n579), .B2(new_n557), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n559), .A2(new_n557), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n546), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n325), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n530), .A2(new_n544), .A3(KEYINPUT77), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n518), .A2(new_n527), .ZN(new_n586));
  OR2_X1    g400(.A1(new_n586), .A2(new_n543), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT77), .B1(new_n530), .B2(new_n544), .ZN(new_n589));
  OAI21_X1  g403(.A(KEYINPUT28), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n590), .A2(KEYINPUT29), .A3(new_n581), .ZN(new_n591));
  OAI21_X1  g405(.A(G472), .B1(new_n584), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n514), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n571), .A2(new_n576), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n549), .A2(new_n516), .A3(new_n557), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT76), .B1(new_n560), .B2(new_n556), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n593), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n578), .B(new_n592), .C1(new_n598), .C2(KEYINPUT32), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n458), .A2(new_n246), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n476), .A2(new_n478), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT79), .B1(new_n191), .B2(G128), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT79), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n603), .A2(new_n258), .A3(G119), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n191), .A2(G128), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n602), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT24), .B(G110), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT81), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT23), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n610), .B1(new_n191), .B2(G128), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n258), .A2(KEYINPUT23), .A3(G119), .ZN(new_n612));
  INV_X1    g426(.A(G110), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n611), .A2(new_n612), .A3(new_n613), .A4(new_n605), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n608), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n608), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT81), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n601), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n611), .A2(new_n605), .A3(new_n612), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(G110), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n620), .B1(new_n607), .B2(new_n606), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n489), .B2(new_n490), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n269), .A2(G221), .A3(G234), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT83), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT22), .B(G137), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n618), .A2(new_n622), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n617), .A2(new_n615), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n629), .A2(new_n478), .A3(new_n476), .A4(new_n600), .ZN(new_n630));
  INV_X1    g444(.A(new_n622), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n626), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n325), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(KEYINPUT84), .A3(KEYINPUT25), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT25), .ZN(new_n635));
  INV_X1    g449(.A(new_n325), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n627), .B1(new_n618), .B2(new_n622), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n630), .A2(new_n631), .A3(new_n626), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT84), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n635), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n439), .B1(new_n325), .B2(G234), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n634), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n642), .A2(G902), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n637), .A2(new_n638), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n513), .A2(new_n599), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G101), .ZN(G3));
  AOI22_X1  g463(.A1(new_n404), .A2(new_n389), .B1(new_n406), .B2(new_n387), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n401), .B1(new_n650), .B2(G469), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n412), .B1(new_n651), .B2(new_n400), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n647), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n514), .B1(new_n562), .B2(new_n577), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n325), .B1(new_n562), .B2(new_n577), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(G472), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n654), .A2(KEYINPUT101), .A3(new_n655), .A4(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT101), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n655), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n659), .B1(new_n660), .B2(new_n653), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n444), .A2(KEYINPUT33), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT33), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n442), .A2(new_n664), .A3(new_n443), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n636), .A2(new_n448), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n445), .A2(new_n448), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n511), .A2(new_n328), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n662), .A2(new_n333), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT34), .B(G104), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G6));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n510), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT103), .A4(new_n509), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n496), .B1(KEYINPUT102), .B2(KEYINPUT20), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT102), .B(KEYINPUT20), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n494), .A2(new_n495), .A3(new_n680), .ZN(new_n681));
  AOI22_X1  g495(.A1(new_n679), .A2(new_n681), .B1(new_n447), .B2(new_n449), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n333), .A2(new_n678), .A3(new_n329), .A4(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n662), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT35), .B(G107), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G9));
  NAND2_X1  g501(.A1(new_n630), .A2(new_n631), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n626), .A2(KEYINPUT36), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n645), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n643), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n643), .A2(KEYINPUT104), .A3(new_n691), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n636), .B1(new_n594), .B2(new_n597), .ZN(new_n697));
  INV_X1    g511(.A(G472), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n655), .B(new_n696), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n657), .A2(KEYINPUT105), .A3(new_n655), .A4(new_n696), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n701), .A2(new_n513), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT37), .B(G110), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT106), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n703), .B(new_n705), .ZN(G12));
  AND3_X1   g520(.A1(new_n409), .A2(new_n413), .A3(new_n696), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n599), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(G900), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n324), .B1(new_n326), .B2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n676), .A2(new_n682), .A3(new_n677), .A4(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(KEYINPUT107), .A3(new_n333), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT107), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n320), .B2(new_n712), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n708), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G128), .ZN(G30));
  NAND2_X1  g533(.A1(new_n579), .A2(new_n556), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n293), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n588), .A2(new_n556), .A3(new_n589), .ZN(new_n722));
  OAI21_X1  g536(.A(G472), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n578), .B(new_n723), .C1(new_n598), .C2(KEYINPUT32), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(KEYINPUT108), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(new_n710), .B(KEYINPUT39), .Z(new_n727));
  NAND2_X1  g541(.A1(new_n652), .A2(new_n727), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n728), .A2(KEYINPUT40), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n331), .A2(new_n332), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT38), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n696), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n450), .B1(new_n501), .B2(new_n510), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n733), .A2(new_n187), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n728), .A2(KEYINPUT40), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n729), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n726), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT109), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n726), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(new_n250), .ZN(G45));
  NOR3_X1   g558(.A1(new_n511), .A2(new_n670), .A3(new_n710), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n333), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n708), .A2(new_n747), .ZN(new_n748));
  XOR2_X1   g562(.A(KEYINPUT110), .B(G146), .Z(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G48));
  NAND2_X1  g564(.A1(new_n382), .A2(new_n387), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n751), .A2(new_n389), .B1(new_n406), .B2(new_n403), .ZN(new_n752));
  OAI21_X1  g566(.A(G469), .B1(new_n752), .B2(new_n636), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n411), .A3(new_n400), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n754), .A2(new_n320), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n599), .A2(new_n755), .A3(new_n647), .A4(new_n671), .ZN(new_n756));
  XNOR2_X1  g570(.A(KEYINPUT41), .B(G113), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(G15));
  INV_X1    g572(.A(new_n754), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n599), .A2(new_n647), .A3(new_n684), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G116), .ZN(G18));
  AND4_X1   g575(.A1(new_n329), .A2(new_n696), .A3(new_n450), .A4(new_n511), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n599), .A2(new_n762), .A3(new_n755), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G119), .ZN(G21));
  NAND3_X1  g578(.A1(new_n333), .A2(new_n329), .A3(new_n735), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n754), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n590), .A2(new_n548), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n557), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n575), .A2(KEYINPUT31), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(new_n569), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n593), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n771), .B1(new_n656), .B2(G472), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n766), .A2(new_n772), .A3(new_n647), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G122), .ZN(G24));
  NAND4_X1  g588(.A1(new_n772), .A2(new_n696), .A3(new_n747), .A4(new_n759), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G125), .ZN(G27));
  AND4_X1   g590(.A1(new_n187), .A2(new_n331), .A3(new_n332), .A4(new_n411), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n409), .A2(new_n745), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n599), .A2(new_n647), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT42), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n599), .A2(new_n778), .A3(KEYINPUT42), .A4(new_n647), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G131), .ZN(G33));
  AND3_X1   g598(.A1(new_n409), .A2(new_n713), .A3(new_n777), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n599), .A2(new_n647), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G134), .ZN(G36));
  NAND2_X1  g601(.A1(new_n501), .A2(new_n510), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n788), .A2(new_n670), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT43), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n734), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(KEYINPUT44), .A3(new_n660), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT111), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n405), .A2(new_n407), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n336), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n650), .A2(KEYINPUT45), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n402), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT46), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n400), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n799), .A2(new_n800), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n411), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT44), .B1(new_n791), .B2(new_n660), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n331), .A2(new_n187), .A3(new_n332), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n793), .A2(new_n727), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G137), .ZN(G39));
  INV_X1    g624(.A(KEYINPUT47), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n804), .B(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n511), .A2(new_n670), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n711), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n599), .A2(new_n647), .A3(new_n814), .A4(new_n807), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  NOR2_X1   g631(.A1(new_n754), .A2(new_n807), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n725), .A2(new_n647), .A3(new_n324), .A4(new_n818), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n819), .A2(KEYINPUT115), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(KEYINPUT115), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(new_n511), .A3(new_n670), .A4(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n324), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n790), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n772), .A2(new_n647), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n807), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n753), .A2(new_n400), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n829), .A2(new_n412), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n828), .B1(new_n812), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT50), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n733), .A2(new_n187), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n759), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n832), .B1(new_n827), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n826), .A2(KEYINPUT50), .A3(new_n759), .A4(new_n833), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n772), .A2(new_n696), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n824), .A2(new_n754), .A3(new_n807), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n835), .A2(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n822), .A2(new_n831), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT51), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n826), .A2(new_n755), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(G952), .A3(new_n269), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n599), .A2(new_n647), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n839), .A2(new_n846), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n847), .B(KEYINPUT48), .Z(new_n848));
  AND2_X1   g662(.A1(new_n820), .A2(new_n821), .ZN(new_n849));
  AOI211_X1 g663(.A(new_n845), .B(new_n848), .C1(new_n849), .C2(new_n813), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n841), .A2(new_n842), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n843), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n679), .A2(new_n681), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n678), .A2(new_n450), .A3(new_n854), .A4(new_n711), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n855), .A2(new_n807), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n599), .A2(new_n707), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n772), .A2(new_n778), .A3(new_n696), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n786), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n781), .B2(new_n782), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n333), .B(new_n321), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n788), .A2(new_n450), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n861), .A2(KEYINPUT112), .A3(new_n329), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n861), .A2(new_n671), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n322), .A2(new_n334), .A3(new_n329), .A4(new_n862), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT112), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n863), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(new_n661), .A3(new_n658), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n703), .A2(new_n648), .ZN(new_n870));
  AND4_X1   g684(.A1(new_n756), .A2(new_n760), .A3(new_n763), .A4(new_n773), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n860), .A2(new_n869), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n599), .B(new_n707), .C1(new_n717), .C2(new_n747), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n333), .A2(new_n735), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n411), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n692), .A2(new_n876), .A3(new_n710), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n724), .A2(new_n409), .A3(new_n875), .A4(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n873), .A2(new_n878), .A3(new_n775), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT52), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n853), .B1(new_n872), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT113), .ZN(new_n882));
  INV_X1    g696(.A(new_n859), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n871), .A2(new_n783), .A3(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT52), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n879), .B(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n869), .A2(new_n648), .A3(new_n703), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n884), .A2(new_n886), .A3(KEYINPUT53), .A4(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n881), .A2(new_n882), .A3(new_n888), .ZN(new_n889));
  OAI211_X1 g703(.A(KEYINPUT113), .B(new_n853), .C1(new_n872), .C2(new_n880), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(KEYINPUT54), .A3(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n881), .A2(new_n892), .A3(new_n888), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT114), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT114), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n881), .A2(new_n888), .A3(new_n895), .A4(new_n892), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n891), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  OAI22_X1  g711(.A1(new_n852), .A2(new_n897), .B1(G952), .B2(G953), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n647), .A2(new_n187), .A3(new_n413), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n733), .A2(new_n789), .A3(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT49), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n829), .A2(new_n901), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n829), .A2(new_n901), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n900), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n898), .B1(new_n726), .B2(new_n904), .ZN(G75));
  NOR2_X1   g719(.A1(new_n269), .A2(G952), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n881), .A2(new_n888), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n636), .A3(new_n307), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n309), .A2(new_n311), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n278), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n312), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT55), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n914), .A2(KEYINPUT56), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n907), .B1(new_n910), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT116), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT56), .B1(new_n909), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n918), .B1(new_n917), .B2(new_n909), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n916), .B1(new_n919), .B2(new_n914), .ZN(G51));
  AOI211_X1 g734(.A(new_n325), .B(new_n798), .C1(new_n881), .C2(new_n888), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n401), .B(KEYINPUT117), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT57), .Z(new_n923));
  AND3_X1   g737(.A1(new_n881), .A2(new_n892), .A3(new_n888), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n892), .B1(new_n881), .B2(new_n888), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n752), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n921), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT118), .ZN(new_n929));
  OR3_X1    g743(.A1(new_n928), .A2(new_n929), .A3(new_n906), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n929), .B1(new_n928), .B2(new_n906), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(G54));
  AND2_X1   g746(.A1(KEYINPUT58), .A2(G475), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n908), .A2(new_n636), .A3(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n494), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n906), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n935), .B2(new_n934), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT119), .ZN(G60));
  XNOR2_X1  g752(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n448), .A2(new_n293), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n897), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n666), .B(KEYINPUT120), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT122), .ZN(new_n945));
  INV_X1    g759(.A(new_n943), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n941), .B(new_n946), .C1(new_n924), .C2(new_n925), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n907), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n944), .A2(new_n945), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n946), .B1(new_n897), .B2(new_n941), .ZN(new_n951));
  OAI21_X1  g765(.A(KEYINPUT122), .B1(new_n951), .B2(new_n948), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(G63));
  NAND2_X1  g767(.A1(G217), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT60), .Z(new_n955));
  AND2_X1   g769(.A1(new_n908), .A2(new_n955), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n956), .A2(new_n646), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n690), .B(KEYINPUT123), .Z(new_n958));
  AOI21_X1  g772(.A(new_n906), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT124), .B1(new_n956), .B2(new_n958), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n961), .A2(KEYINPUT61), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n957), .B(new_n959), .C1(new_n961), .C2(KEYINPUT61), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(G66));
  INV_X1    g779(.A(new_n327), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n269), .B1(new_n966), .B2(G224), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n887), .A2(new_n871), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n967), .B1(new_n968), .B2(new_n269), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n911), .B1(G898), .B2(new_n269), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n969), .B(new_n970), .Z(G69));
  NAND2_X1  g785(.A1(new_n573), .A2(new_n564), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(new_n466), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n805), .A2(new_n727), .A3(new_n875), .ZN(new_n974));
  INV_X1    g788(.A(new_n785), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n846), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n873), .A2(new_n775), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(new_n781), .B2(new_n782), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n977), .A2(new_n816), .A3(new_n809), .A4(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n269), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n269), .A2(G900), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT125), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n973), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n813), .A2(new_n862), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n728), .A2(new_n807), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n846), .A2(new_n986), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n816), .A2(new_n809), .A3(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n978), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n740), .A2(new_n742), .A3(new_n989), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n990), .A2(KEYINPUT62), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(KEYINPUT62), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n988), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n269), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n984), .B1(new_n994), .B2(new_n973), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n269), .B1(G227), .B2(G900), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n995), .B(new_n997), .ZN(G72));
  INV_X1    g812(.A(new_n968), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n988), .A2(new_n991), .A3(new_n999), .A4(new_n992), .ZN(new_n1000));
  NAND2_X1  g814(.A1(G472), .A2(G902), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT63), .Z(new_n1002));
  NAND2_X1  g816(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n720), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n579), .A2(new_n556), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1002), .ZN(new_n1007));
  NOR3_X1   g821(.A1(new_n1004), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n889), .A2(new_n890), .A3(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1002), .B1(new_n980), .B2(new_n968), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n906), .B1(new_n1010), .B2(new_n1006), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1005), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(KEYINPUT126), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT126), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1005), .A2(new_n1014), .A3(new_n1009), .A4(new_n1011), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1013), .A2(new_n1015), .ZN(G57));
endmodule


