//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n991, new_n992, new_n993, new_n994, new_n995;
  INV_X1    g000(.A(G134gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G127gat), .ZN(new_n203));
  INV_X1    g002(.A(G127gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G134gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G113gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G120gat), .ZN(new_n209));
  OR2_X1    g008(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(G113gat), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n207), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G120gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G113gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n216), .A2(new_n206), .B1(new_n203), .B2(new_n205), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n220), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223));
  INV_X1    g022(.A(G183gat), .ZN(new_n224));
  INV_X1    g023(.A(G190gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n225), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n221), .A2(new_n222), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G169gat), .ZN(new_n229));
  INV_X1    g028(.A(G176gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n233), .A2(KEYINPUT23), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(KEYINPUT23), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n228), .A2(new_n232), .A3(new_n234), .A4(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AND4_X1   g037(.A1(KEYINPUT25), .A2(new_n234), .A3(new_n232), .A4(new_n235), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n223), .A2(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(KEYINPUT66), .B2(new_n223), .ZN(new_n241));
  OR2_X1    g040(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n241), .B(new_n219), .C1(G183gat), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n239), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n238), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n233), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n231), .B1(KEYINPUT26), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT26), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n250), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n249), .A2(new_n251), .B1(G183gat), .B2(G190gat), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT27), .B1(new_n254), .B2(new_n224), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT27), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n256), .A2(KEYINPUT68), .A3(G183gat), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n255), .A2(new_n257), .A3(new_n242), .A4(new_n243), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT28), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT27), .B(G183gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n244), .A2(new_n259), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n260), .A2(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n258), .A2(KEYINPUT69), .A3(new_n259), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n253), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n247), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n258), .A2(KEYINPUT69), .A3(new_n259), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT69), .B1(new_n258), .B2(new_n259), .ZN(new_n270));
  AND4_X1   g069(.A1(KEYINPUT28), .A2(new_n262), .A3(new_n242), .A4(new_n243), .ZN(new_n271));
  NOR3_X1   g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n272), .A2(KEYINPUT70), .A3(new_n253), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n218), .B1(new_n268), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT70), .B1(new_n272), .B2(new_n253), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n264), .A2(new_n265), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n276), .A2(new_n267), .A3(new_n252), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n216), .A2(new_n206), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n203), .A2(new_n205), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n212), .A2(new_n209), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n280), .B1(new_n281), .B2(new_n207), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n275), .A2(new_n277), .A3(new_n282), .A4(new_n247), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n274), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G227gat), .ZN(new_n285));
  INV_X1    g084(.A(G233gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT74), .B1(new_n289), .B2(KEYINPUT34), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(KEYINPUT34), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT74), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT34), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n284), .A2(new_n292), .A3(new_n293), .A4(new_n288), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n290), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n274), .A2(new_n287), .A3(new_n283), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT32), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT33), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT72), .B(G71gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(G99gat), .ZN(new_n301));
  XOR2_X1   g100(.A(G15gat), .B(G43gat), .Z(new_n302));
  XOR2_X1   g101(.A(new_n301), .B(new_n302), .Z(new_n303));
  NAND3_X1  g102(.A1(new_n297), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n303), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n296), .B(KEYINPUT32), .C1(new_n298), .C2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n295), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT36), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n304), .A2(KEYINPUT73), .A3(new_n306), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT73), .B1(new_n304), .B2(new_n306), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n295), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n295), .A2(new_n307), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n309), .B1(new_n316), .B2(new_n308), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT85), .ZN(new_n319));
  INV_X1    g118(.A(G155gat), .ZN(new_n320));
  INV_X1    g119(.A(G162gat), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT2), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT79), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XOR2_X1   g123(.A(G141gat), .B(G148gat), .Z(new_n325));
  XNOR2_X1  g124(.A(G155gat), .B(G162gat), .ZN(new_n326));
  OAI211_X1 g125(.A(KEYINPUT79), .B(KEYINPUT2), .C1(new_n320), .C2(new_n321), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n326), .ZN(new_n329));
  XNOR2_X1  g128(.A(G141gat), .B(G148gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n329), .B1(KEYINPUT2), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT4), .B1(new_n282), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT4), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n218), .A2(new_n334), .A3(new_n331), .A4(new_n328), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G225gat), .A2(G233gat), .ZN(new_n337));
  AND3_X1   g136(.A1(new_n328), .A2(new_n331), .A3(KEYINPUT80), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT80), .B1(new_n328), .B2(new_n331), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340));
  NOR3_X1   g139(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n280), .B(KEYINPUT81), .C1(new_n281), .C2(new_n207), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT81), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(new_n213), .B2(new_n217), .ZN(new_n344));
  XOR2_X1   g143(.A(KEYINPUT82), .B(KEYINPUT3), .Z(new_n345));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n331), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n342), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n336), .B(new_n337), .C1(new_n341), .C2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n319), .B1(new_n348), .B2(KEYINPUT5), .ZN(new_n349));
  INV_X1    g148(.A(new_n347), .ZN(new_n350));
  INV_X1    g149(.A(new_n339), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n328), .A2(new_n331), .A3(KEYINPUT80), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(KEYINPUT3), .A3(new_n352), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n350), .A2(new_n353), .B1(new_n333), .B2(new_n335), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT5), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n354), .A2(KEYINPUT85), .A3(new_n355), .A4(new_n337), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n342), .A2(new_n344), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n338), .A2(new_n339), .ZN(new_n359));
  INV_X1    g158(.A(new_n332), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n358), .A2(new_n359), .B1(new_n360), .B2(new_n218), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n348), .B(KEYINPUT5), .C1(new_n337), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  XOR2_X1   g162(.A(KEYINPUT83), .B(KEYINPUT0), .Z(new_n364));
  XNOR2_X1  g163(.A(G57gat), .B(G85gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G1gat), .B(G29gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(KEYINPUT84), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n366), .B(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n363), .A2(KEYINPUT6), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n357), .A2(new_n369), .A3(new_n362), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT6), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n369), .B1(new_n357), .B2(new_n362), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n371), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G226gat), .A2(G233gat), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n275), .A2(new_n277), .A3(new_n247), .A4(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(KEYINPUT29), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n236), .A2(new_n237), .B1(new_n245), .B2(new_n239), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n380), .B1(new_n266), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT75), .B(G211gat), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT22), .B1(new_n384), .B2(G218gat), .ZN(new_n385));
  XOR2_X1   g184(.A(G197gat), .B(G204gat), .Z(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G211gat), .B(G218gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n388), .A2(KEYINPUT76), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n387), .B(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n383), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n380), .B1(new_n268), .B2(new_n273), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n247), .B(new_n378), .C1(new_n272), .C2(new_n253), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(new_n390), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G64gat), .B(G92gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT77), .ZN(new_n398));
  XNOR2_X1  g197(.A(G8gat), .B(G36gat), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n398), .B(new_n399), .Z(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT78), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n400), .B1(new_n392), .B2(new_n395), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT78), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n395), .A3(new_n400), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(KEYINPUT30), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n376), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT29), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n346), .A2(new_n411), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n390), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G228gat), .A2(G233gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n340), .B1(new_n390), .B2(KEYINPUT29), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n359), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  OR2_X1    g217(.A1(new_n385), .A2(new_n386), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT29), .B1(new_n419), .B2(new_n388), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n420), .B1(new_n388), .B2(new_n419), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n360), .B1(new_n421), .B2(new_n345), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n414), .B1(new_n422), .B2(new_n413), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT86), .B(KEYINPUT31), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(G50gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(G78gat), .B(G106gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(G22gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(KEYINPUT87), .A2(G22gat), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n430), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n424), .B(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n410), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT40), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT89), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n436), .B1(new_n354), .B2(new_n337), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n336), .B1(new_n341), .B2(new_n347), .ZN(new_n438));
  INV_X1    g237(.A(new_n337), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(KEYINPUT89), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n361), .A2(new_n337), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n437), .A2(KEYINPUT39), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n369), .B(KEYINPUT88), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT39), .B1(new_n437), .B2(new_n440), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n435), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n443), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n363), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n445), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n449), .A2(KEYINPUT40), .A3(new_n443), .A4(new_n442), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n446), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n407), .A2(new_n409), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n433), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n372), .A2(new_n373), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n454), .A2(new_n448), .B1(KEYINPUT6), .B2(new_n375), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT37), .B1(new_n392), .B2(new_n395), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n393), .A2(new_n394), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT37), .B1(new_n458), .B2(new_n390), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n383), .A2(new_n391), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n400), .A2(KEYINPUT38), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n392), .A2(KEYINPUT37), .A3(new_n395), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n401), .B1(new_n464), .B2(new_n456), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT38), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n455), .A2(new_n408), .A3(new_n463), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n453), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n318), .A2(new_n434), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n433), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n470), .B1(new_n295), .B2(new_n307), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(new_n316), .ZN(new_n472));
  INV_X1    g271(.A(new_n455), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n405), .B(new_n403), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT30), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n408), .B(new_n475), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n474), .A2(new_n476), .A3(KEYINPUT35), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n472), .A2(new_n473), .A3(new_n477), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n290), .A2(new_n291), .A3(new_n294), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT73), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n307), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n479), .B1(new_n481), .B2(new_n311), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n482), .A2(new_n410), .A3(new_n471), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT35), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n478), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n485), .ZN(new_n486));
  XOR2_X1   g285(.A(G169gat), .B(G197gat), .Z(new_n487));
  XNOR2_X1  g286(.A(G113gat), .B(G141gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT12), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(G29gat), .ZN(new_n494));
  INV_X1    g293(.A(G36gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT14), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT14), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n497), .B1(G29gat), .B2(G36gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(G29gat), .A2(G36gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(G50gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(G43gat), .ZN(new_n502));
  INV_X1    g301(.A(G43gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(G50gat), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n502), .A2(new_n504), .A3(KEYINPUT15), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n500), .B(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(KEYINPUT91), .B(G50gat), .Z(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n503), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT15), .B1(new_n508), .B2(new_n502), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT17), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n505), .A2(new_n498), .A3(new_n499), .A4(new_n496), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT15), .B1(new_n503), .B2(G50gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n501), .A2(G43gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n500), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT91), .B(G50gat), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n502), .B1(new_n516), .B2(G43gat), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT15), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n511), .A2(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT17), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(G1gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT16), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n429), .A2(G15gat), .ZN(new_n524));
  INV_X1    g323(.A(G15gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(G22gat), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(G1gat), .B1(new_n524), .B2(new_n526), .ZN(new_n528));
  OAI21_X1  g327(.A(G8gat), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n530));
  INV_X1    g329(.A(G8gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(G15gat), .B(G22gat), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n530), .B(new_n531), .C1(G1gat), .C2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n510), .A2(new_n521), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT92), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT92), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n510), .A2(new_n521), .A3(new_n538), .A4(new_n535), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G229gat), .A2(G233gat), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n519), .A2(new_n534), .A3(KEYINPUT93), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT93), .B1(new_n519), .B2(new_n534), .ZN(new_n543));
  OAI211_X1 g342(.A(KEYINPUT18), .B(new_n541), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  OAI22_X1  g345(.A1(new_n542), .A2(new_n543), .B1(new_n519), .B2(new_n534), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n541), .B(KEYINPUT94), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT13), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n543), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n519), .A2(new_n534), .A3(KEYINPUT93), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n552), .A2(new_n553), .B1(G229gat), .B2(G233gat), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT18), .B1(new_n540), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n493), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n511), .A2(new_n515), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n517), .A2(new_n518), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n557), .A2(new_n520), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n520), .B1(new_n557), .B2(new_n558), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n538), .B1(new_n561), .B2(new_n535), .ZN(new_n562));
  INV_X1    g361(.A(new_n539), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n554), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT18), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n540), .A2(new_n545), .B1(new_n547), .B2(new_n549), .ZN(new_n567));
  INV_X1    g366(.A(new_n493), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n556), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n486), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(G57gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(G64gat), .ZN(new_n573));
  INV_X1    g372(.A(G64gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(G57gat), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT9), .ZN(new_n576));
  NAND2_X1  g375(.A1(G71gat), .A2(G78gat), .ZN(new_n577));
  AOI22_X1  g376(.A1(new_n573), .A2(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(G71gat), .A2(G78gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n577), .B(KEYINPUT95), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n577), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT96), .ZN(new_n584));
  NOR3_X1   g383(.A1(new_n583), .A2(new_n579), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n579), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT96), .B1(new_n586), .B2(new_n577), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n578), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT21), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n535), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(new_n224), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n590), .ZN(new_n593));
  XNOR2_X1  g392(.A(G127gat), .B(G155gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n592), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n597));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT97), .B(G211gat), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n599), .B(new_n600), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n596), .B(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AND2_X1   g402(.A1(G232gat), .A2(G233gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n604), .A2(KEYINPUT41), .ZN(new_n605));
  XNOR2_X1  g404(.A(G190gat), .B(G218gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G99gat), .A2(G106gat), .ZN(new_n609));
  INV_X1    g408(.A(G85gat), .ZN(new_n610));
  INV_X1    g409(.A(G92gat), .ZN(new_n611));
  AOI22_X1  g410(.A1(KEYINPUT8), .A2(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g411(.A1(KEYINPUT98), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n613));
  NAND3_X1  g412(.A1(KEYINPUT98), .A2(G85gat), .A3(G92gat), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT7), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n612), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  OR2_X1    g416(.A1(G99gat), .A2(G106gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n609), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n612), .A2(new_n613), .A3(new_n616), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n621), .A2(new_n609), .A3(new_n618), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n561), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n623), .ZN(new_n627));
  AOI22_X1  g426(.A1(new_n627), .A2(new_n519), .B1(KEYINPUT41), .B2(new_n604), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n624), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n626), .B1(new_n624), .B2(new_n628), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n608), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n631), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n633), .A2(new_n607), .A3(new_n629), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT10), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n623), .A2(new_n589), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n621), .A2(KEYINPUT99), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n619), .A2(KEYINPUT100), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT100), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n618), .A2(new_n641), .A3(new_n609), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n612), .A2(new_n644), .A3(new_n613), .A4(new_n616), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n639), .A2(KEYINPUT101), .A3(new_n643), .A4(new_n645), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n646), .A2(new_n588), .A3(new_n582), .A4(new_n620), .ZN(new_n647));
  AOI22_X1  g446(.A1(new_n617), .A2(new_n644), .B1(new_n640), .B2(new_n642), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT101), .B1(new_n648), .B2(new_n639), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n637), .B(new_n638), .C1(new_n647), .C2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n589), .A2(new_n637), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n627), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G230gat), .A2(G233gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n638), .B1(new_n647), .B2(new_n649), .ZN(new_n656));
  INV_X1    g455(.A(new_n654), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G120gat), .B(G148gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G176gat), .ZN(new_n661));
  INV_X1    g460(.A(G204gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n655), .A2(new_n658), .A3(new_n663), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n603), .A2(new_n636), .A3(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n571), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n376), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n452), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT102), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n676), .B(KEYINPUT16), .Z(new_n677));
  OR2_X1    g476(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n678), .A2(G8gat), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n674), .A2(new_n675), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(G8gat), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(G1325gat));
  OR2_X1    g481(.A1(new_n316), .A2(new_n308), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n670), .A2(new_n525), .A3(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n571), .A2(new_n318), .A3(new_n669), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n685), .B1(new_n525), .B2(new_n686), .ZN(G1326gat));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n433), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT43), .B(G22gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  NAND2_X1  g489(.A1(new_n602), .A2(new_n668), .ZN(new_n691));
  INV_X1    g490(.A(new_n570), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n636), .A2(KEYINPUT44), .ZN(new_n695));
  INV_X1    g494(.A(new_n307), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n433), .B1(new_n696), .B2(new_n479), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n474), .A2(new_n476), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n314), .A2(new_n697), .A3(new_n698), .A4(new_n376), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n452), .A2(new_n455), .A3(KEYINPUT35), .ZN(new_n700));
  AOI22_X1  g499(.A1(new_n699), .A2(KEYINPUT35), .B1(new_n700), .B2(new_n472), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n469), .B1(new_n701), .B2(KEYINPUT103), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n485), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n695), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n453), .A2(new_n467), .B1(new_n410), .B2(new_n433), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n699), .A2(KEYINPUT35), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n318), .A2(new_n706), .B1(new_n707), .B2(new_n478), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT44), .B1(new_n708), .B2(new_n636), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n694), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(G29gat), .B1(new_n711), .B2(new_n376), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n708), .A2(new_n692), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n691), .A2(new_n636), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n713), .A2(new_n494), .A3(new_n671), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT45), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n712), .A2(new_n716), .ZN(G1328gat));
  INV_X1    g516(.A(new_n714), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n495), .B1(new_n719), .B2(KEYINPUT104), .ZN(new_n720));
  NOR4_X1   g519(.A1(new_n571), .A2(new_n698), .A3(new_n718), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(KEYINPUT104), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G36gat), .B1(new_n711), .B2(new_n698), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(G1329gat));
  XNOR2_X1  g524(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n684), .A2(new_n503), .A3(new_n714), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n713), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT107), .B1(new_n571), .B2(new_n728), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n318), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n503), .B1(new_n710), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n732), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n695), .ZN(new_n737));
  AOI22_X1  g536(.A1(new_n485), .A2(new_n703), .B1(new_n318), .B2(new_n706), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n701), .A2(KEYINPUT103), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n741), .B1(new_n486), .B2(new_n635), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n733), .B(new_n693), .C1(new_n740), .C2(new_n742), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n743), .A2(new_n735), .A3(G43gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n726), .B1(new_n736), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n732), .A2(KEYINPUT47), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n503), .B1(new_n743), .B2(KEYINPUT108), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n705), .A2(new_n709), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n749), .A2(new_n750), .A3(new_n733), .A4(new_n693), .ZN(new_n751));
  AOI211_X1 g550(.A(new_n746), .B(new_n747), .C1(new_n748), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n743), .A2(KEYINPUT108), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n753), .A2(G43gat), .A3(new_n751), .ZN(new_n754));
  INV_X1    g553(.A(new_n747), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT109), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n745), .B1(new_n752), .B2(new_n756), .ZN(G1330gat));
  NAND3_X1  g556(.A1(new_n714), .A2(new_n433), .A3(new_n516), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n759));
  OAI22_X1  g558(.A1(new_n571), .A2(new_n758), .B1(new_n759), .B2(KEYINPUT48), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n710), .A2(new_n433), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n760), .B1(new_n761), .B2(new_n507), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n759), .A2(KEYINPUT48), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n762), .B(new_n763), .Z(G1331gat));
  NAND2_X1  g563(.A1(new_n738), .A2(new_n739), .ZN(new_n765));
  NOR4_X1   g564(.A1(new_n602), .A2(new_n668), .A3(new_n570), .A4(new_n635), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n671), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n452), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n771));
  XOR2_X1   g570(.A(KEYINPUT49), .B(G64gat), .Z(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n770), .B2(new_n772), .ZN(G1333gat));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n774));
  INV_X1    g573(.A(G71gat), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n767), .A2(new_n775), .A3(new_n684), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n765), .A2(new_n766), .ZN(new_n777));
  OAI21_X1  g576(.A(G71gat), .B1(new_n777), .B2(new_n318), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT111), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n779), .B1(new_n776), .B2(new_n778), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n774), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n782), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n784), .A2(KEYINPUT50), .A3(new_n780), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(G1334gat));
  NAND2_X1  g585(.A1(new_n767), .A2(new_n433), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g587(.A1(new_n603), .A2(new_n570), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n749), .A2(new_n667), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(G85gat), .B1(new_n790), .B2(new_n376), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n603), .A2(new_n570), .A3(new_n636), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n702), .B2(new_n704), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n765), .A2(KEYINPUT51), .A3(new_n792), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n671), .A2(new_n610), .A3(new_n667), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n799), .B(KEYINPUT112), .Z(new_n800));
  OAI21_X1  g599(.A(new_n791), .B1(new_n798), .B2(new_n800), .ZN(G1336gat));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n668), .B1(new_n795), .B2(new_n796), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n803), .A2(new_n611), .A3(new_n452), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n802), .B1(new_n804), .B2(KEYINPUT113), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n698), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n806), .B2(new_n611), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  OAI221_X1 g607(.A(new_n804), .B1(KEYINPUT113), .B2(new_n802), .C1(new_n806), .C2(new_n611), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(G1337gat));
  INV_X1    g609(.A(G99gat), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n803), .A2(new_n811), .A3(new_n684), .ZN(new_n812));
  OAI21_X1  g611(.A(G99gat), .B1(new_n790), .B2(new_n318), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(G1338gat));
  NOR2_X1   g613(.A1(new_n470), .A2(G106gat), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n803), .A2(KEYINPUT114), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(G106gat), .B1(new_n790), .B2(new_n470), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n816), .A2(new_n817), .A3(KEYINPUT115), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n819));
  NAND2_X1  g618(.A1(KEYINPUT115), .A2(KEYINPUT53), .ZN(new_n820));
  AOI22_X1  g619(.A1(new_n803), .A2(new_n815), .B1(KEYINPUT114), .B2(new_n820), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n818), .A2(new_n819), .B1(new_n817), .B2(new_n821), .ZN(G1339gat));
  NAND4_X1  g621(.A1(new_n603), .A2(new_n692), .A3(new_n636), .A4(new_n668), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n552), .A2(new_n553), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n541), .B1(new_n540), .B2(new_n825), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n547), .A2(new_n549), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n491), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n635), .A2(new_n569), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n654), .B1(new_n651), .B2(new_n627), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n650), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT54), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n657), .B1(new_n650), .B2(new_n652), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT55), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n653), .A2(new_n836), .A3(new_n654), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n664), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n666), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n655), .A2(KEYINPUT54), .A3(new_n832), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n663), .B1(new_n834), .B2(new_n836), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT55), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT116), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n837), .B(new_n664), .C1(new_n833), .C2(new_n834), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n840), .A2(new_n841), .A3(KEYINPUT55), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n846), .A2(new_n847), .A3(new_n666), .A4(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n830), .B1(new_n843), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n667), .A2(new_n569), .A3(new_n829), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n843), .A2(new_n849), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(new_n570), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n851), .B1(new_n855), .B2(new_n635), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n824), .B1(new_n856), .B2(new_n602), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n698), .A2(new_n671), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n472), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n860), .A2(new_n208), .A3(new_n692), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n482), .A2(new_n471), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n570), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n861), .B1(new_n208), .B2(new_n865), .ZN(G1340gat));
  OAI21_X1  g665(.A(G120gat), .B1(new_n860), .B2(new_n668), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n667), .A2(new_n210), .A3(new_n211), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n867), .B1(new_n863), .B2(new_n868), .ZN(G1341gat));
  OAI21_X1  g668(.A(G127gat), .B1(new_n860), .B2(new_n602), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n603), .A2(new_n204), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n863), .B2(new_n871), .ZN(G1342gat));
  NOR3_X1   g671(.A1(new_n863), .A2(G134gat), .A3(new_n636), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n875));
  OAI21_X1  g674(.A(G134gat), .B1(new_n860), .B2(new_n636), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(G1343gat));
  NAND2_X1  g677(.A1(new_n856), .A2(new_n602), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n823), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n318), .A2(new_n671), .A3(new_n698), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n880), .A2(new_n433), .A3(new_n882), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n883), .A2(G141gat), .A3(new_n692), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n885), .B1(new_n857), .B2(new_n470), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n470), .A2(new_n885), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n570), .A2(new_n666), .A3(new_n846), .A4(new_n848), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n635), .B1(new_n888), .B2(new_n852), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n602), .B1(new_n889), .B2(new_n850), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n890), .A2(KEYINPUT117), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n823), .B1(new_n890), .B2(KEYINPUT117), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n887), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n881), .B1(new_n886), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n570), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n884), .B1(new_n895), .B2(G141gat), .ZN(new_n896));
  XOR2_X1   g695(.A(new_n896), .B(KEYINPUT58), .Z(G1344gat));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n830), .A2(new_n842), .A3(new_n839), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n544), .B1(new_n537), .B2(new_n539), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n547), .A2(new_n549), .ZN(new_n901));
  NOR4_X1   g700(.A1(new_n555), .A2(new_n900), .A3(new_n901), .A4(new_n493), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n568), .B1(new_n566), .B2(new_n567), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n666), .B(new_n848), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n852), .B1(new_n904), .B2(new_n842), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n899), .B1(new_n905), .B2(new_n636), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n823), .B1(new_n906), .B2(new_n603), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n470), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n602), .B1(new_n889), .B2(new_n899), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(KEYINPUT119), .A3(new_n823), .ZN(new_n911));
  AOI21_X1  g710(.A(KEYINPUT57), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n887), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n857), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n667), .B(new_n882), .C1(new_n912), .C2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT120), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n880), .A2(new_n887), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n910), .A2(KEYINPUT119), .A3(new_n823), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT119), .B1(new_n910), .B2(new_n823), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n918), .A2(new_n919), .A3(new_n470), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n917), .B1(new_n920), .B2(KEYINPUT57), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n921), .A2(new_n922), .A3(new_n667), .A4(new_n882), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n916), .A2(new_n923), .A3(G148gat), .ZN(new_n924));
  AOI211_X1 g723(.A(new_n668), .B(new_n881), .C1(new_n886), .C2(new_n893), .ZN(new_n925));
  INV_X1    g724(.A(G148gat), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n926), .A2(KEYINPUT59), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT118), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n886), .A2(new_n893), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(new_n667), .A3(new_n882), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT118), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n931), .A2(new_n932), .A3(new_n927), .ZN(new_n933));
  AOI22_X1  g732(.A1(new_n924), .A2(KEYINPUT59), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n883), .A2(G148gat), .A3(new_n668), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n898), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(new_n935), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n929), .A2(new_n933), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT59), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n926), .B1(new_n915), .B2(KEYINPUT120), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(new_n923), .ZN(new_n941));
  OAI211_X1 g740(.A(KEYINPUT121), .B(new_n937), .C1(new_n938), .C2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n936), .A2(new_n942), .ZN(G1345gat));
  NOR3_X1   g742(.A1(new_n883), .A2(G155gat), .A3(new_n602), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n894), .A2(new_n603), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(G155gat), .ZN(new_n946));
  XOR2_X1   g745(.A(new_n946), .B(KEYINPUT122), .Z(G1346gat));
  AND2_X1   g746(.A1(new_n894), .A2(new_n635), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n635), .A2(new_n321), .ZN(new_n949));
  OAI22_X1  g748(.A1(new_n948), .A2(new_n321), .B1(new_n883), .B2(new_n949), .ZN(G1347gat));
  NOR2_X1   g749(.A1(new_n857), .A2(new_n671), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n951), .A2(new_n452), .A3(new_n472), .ZN(new_n952));
  OAI21_X1  g751(.A(G169gat), .B1(new_n952), .B2(new_n692), .ZN(new_n953));
  XOR2_X1   g752(.A(new_n953), .B(KEYINPUT123), .Z(new_n954));
  NAND3_X1  g753(.A1(new_n951), .A2(new_n452), .A3(new_n862), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n570), .A2(new_n229), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(G1348gat));
  OAI21_X1  g756(.A(G176gat), .B1(new_n952), .B2(new_n668), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n667), .A2(new_n230), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n955), .B2(new_n959), .ZN(G1349gat));
  OAI21_X1  g759(.A(G183gat), .B1(new_n952), .B2(new_n602), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n603), .A2(new_n262), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n955), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g763(.A(G190gat), .B1(new_n952), .B2(new_n636), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT61), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n635), .A2(new_n242), .A3(new_n243), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n955), .B2(new_n967), .ZN(G1351gat));
  INV_X1    g767(.A(G197gat), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n733), .A2(new_n698), .A3(new_n470), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n951), .A2(new_n969), .A3(new_n570), .A4(new_n970), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT124), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n733), .A2(new_n671), .A3(new_n698), .ZN(new_n973));
  XOR2_X1   g772(.A(new_n973), .B(KEYINPUT125), .Z(new_n974));
  INV_X1    g773(.A(new_n921), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n974), .A2(new_n975), .A3(new_n692), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n972), .B1(new_n976), .B2(new_n969), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n977), .B(new_n978), .ZN(G1352gat));
  NAND2_X1  g778(.A1(new_n951), .A2(new_n970), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n980), .A2(G204gat), .A3(new_n668), .ZN(new_n981));
  XNOR2_X1  g780(.A(new_n981), .B(KEYINPUT62), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n921), .A2(new_n667), .ZN(new_n983));
  OAI21_X1  g782(.A(G204gat), .B1(new_n974), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(new_n984), .ZN(G1353gat));
  NAND2_X1  g784(.A1(new_n973), .A2(new_n603), .ZN(new_n986));
  OAI21_X1  g785(.A(G211gat), .B1(new_n975), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g786(.A(new_n987), .B(KEYINPUT63), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n980), .A2(new_n384), .A3(new_n602), .ZN(new_n989));
  OR2_X1    g788(.A1(new_n988), .A2(new_n989), .ZN(G1354gat));
  INV_X1    g789(.A(new_n980), .ZN(new_n991));
  AOI21_X1  g790(.A(G218gat), .B1(new_n991), .B2(new_n635), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n635), .A2(G218gat), .ZN(new_n993));
  XNOR2_X1  g792(.A(new_n993), .B(KEYINPUT127), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n974), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n992), .B1(new_n995), .B2(new_n921), .ZN(G1355gat));
endmodule


