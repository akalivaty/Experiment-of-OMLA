//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 0 0 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n544,
    new_n546, new_n547, new_n548, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n599, new_n601, new_n602, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT64), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT65), .Z(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n460), .A2(new_n461), .A3(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(KEYINPUT66), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n465));
  OAI211_X1 g040(.A(new_n459), .B(new_n462), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G137), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n463), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  XNOR2_X1  g045(.A(new_n470), .B(KEYINPUT67), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n461), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n468), .A2(new_n471), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n482));
  INV_X1    g057(.A(G136), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n482), .B1(new_n466), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g059(.A(G2105), .B(new_n462), .C1(new_n464), .C2(new_n465), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n484), .B1(G124), .B2(new_n486), .ZN(G162));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT4), .B1(new_n466), .B2(new_n488), .ZN(new_n489));
  OR3_X1    g064(.A1(new_n488), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(new_n475), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n459), .A2(G114), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(new_n486), .B2(G126), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT68), .B(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n508), .A2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XOR2_X1   g092(.A(new_n517), .B(KEYINPUT7), .Z(new_n518));
  AND2_X1   g093(.A1(new_n505), .A2(new_n509), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n518), .B1(new_n519), .B2(G89), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n521));
  INV_X1    g096(.A(G51), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n512), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT69), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n523), .A2(new_n524), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n520), .B1(new_n525), .B2(new_n526), .ZN(G286));
  INV_X1    g102(.A(G286), .ZN(G168));
  AOI22_X1  g103(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n507), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n510), .A2(new_n531), .B1(new_n512), .B2(new_n532), .ZN(new_n533));
  OR3_X1    g108(.A1(new_n530), .A2(new_n533), .A3(KEYINPUT70), .ZN(new_n534));
  OAI21_X1  g109(.A(KEYINPUT70), .B1(new_n530), .B2(new_n533), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(G171));
  AOI22_X1  g111(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n507), .ZN(new_n538));
  INV_X1    g113(.A(G81), .ZN(new_n539));
  INV_X1    g114(.A(G43), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n510), .A2(new_n539), .B1(new_n512), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  AND3_X1   g118(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G36), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT71), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n544), .A2(new_n548), .ZN(G188));
  NAND2_X1  g124(.A1(new_n519), .A2(G91), .ZN(new_n550));
  INV_X1    g125(.A(new_n512), .ZN(new_n551));
  XNOR2_X1  g126(.A(KEYINPUT72), .B(KEYINPUT9), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n551), .A2(G53), .A3(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  INV_X1    g129(.A(G53), .ZN(new_n555));
  OAI211_X1 g130(.A(KEYINPUT72), .B(new_n554), .C1(new_n512), .C2(new_n555), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n550), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  XNOR2_X1  g133(.A(KEYINPUT73), .B(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n504), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n507), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n562), .B1(new_n561), .B2(new_n560), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n557), .A2(new_n563), .ZN(G299));
  INV_X1    g139(.A(G171), .ZN(G301));
  NAND2_X1  g140(.A1(new_n519), .A2(G87), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n551), .A2(G49), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  AOI22_X1  g144(.A1(new_n505), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n570), .A2(new_n507), .ZN(new_n571));
  INV_X1    g146(.A(G86), .ZN(new_n572));
  INV_X1    g147(.A(G48), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n510), .A2(new_n572), .B1(new_n512), .B2(new_n573), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n571), .A2(new_n574), .ZN(G305));
  AOI22_X1  g150(.A1(new_n519), .A2(G85), .B1(G47), .B2(new_n551), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n576), .B(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n579), .A2(new_n507), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(G290));
  NAND2_X1  g156(.A1(G301), .A2(G868), .ZN(new_n582));
  AND3_X1   g157(.A1(new_n505), .A2(G92), .A3(new_n509), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT76), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT10), .ZN(new_n585));
  NAND2_X1  g160(.A1(G79), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G66), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n504), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(G54), .A2(new_n551), .B1(new_n588), .B2(G651), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n584), .A2(KEYINPUT10), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n582), .B1(new_n592), .B2(G868), .ZN(G284));
  OAI21_X1  g168(.A(new_n582), .B1(new_n592), .B2(G868), .ZN(G321));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(G299), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n596), .B1(G168), .B2(new_n595), .ZN(G297));
  OAI21_X1  g172(.A(new_n596), .B1(G168), .B2(new_n595), .ZN(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n592), .B1(new_n599), .B2(G860), .ZN(G148));
  INV_X1    g175(.A(new_n542), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(new_n595), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n590), .A2(new_n591), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n602), .B1(new_n604), .B2(new_n595), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g181(.A(new_n475), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(new_n469), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT13), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(G2100), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n486), .A2(G123), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n467), .A2(G135), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n459), .A2(G111), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n612), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(G2096), .Z(new_n617));
  NAND2_X1  g192(.A1(new_n611), .A2(new_n617), .ZN(G156));
  XNOR2_X1  g193(.A(KEYINPUT15), .B(G2430), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2435), .ZN(new_n620));
  XNOR2_X1  g195(.A(G2427), .B(G2438), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n622), .A2(KEYINPUT14), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2443), .B(G2446), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2451), .B(G2454), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n626), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G1341), .B(G1348), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(KEYINPUT78), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(KEYINPUT78), .ZN(new_n634));
  INV_X1    g209(.A(G14), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n630), .B2(new_n631), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(G401));
  XNOR2_X1  g213(.A(G2067), .B(G2678), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT79), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g216(.A1(G2072), .A2(G2078), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n442), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT17), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2084), .B(G2090), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n643), .B(KEYINPUT80), .Z(new_n647));
  OAI211_X1 g222(.A(new_n645), .B(new_n646), .C1(new_n641), .C2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT81), .ZN(new_n649));
  NOR3_X1   g224(.A1(new_n640), .A2(new_n643), .A3(new_n646), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT18), .ZN(new_n651));
  OR3_X1    g226(.A1(new_n641), .A2(new_n644), .A3(new_n646), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n649), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(G2100), .Z(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT82), .B(G2096), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G227));
  XNOR2_X1  g232(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT84), .ZN(new_n661));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1956), .B(G2474), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1961), .B(G1966), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT85), .B(KEYINPUT20), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n664), .A2(new_n665), .ZN(new_n671));
  OR3_X1    g246(.A1(new_n663), .A2(new_n666), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n669), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(G1991), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n675), .A2(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(G1996), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n676), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n678), .B1(new_n676), .B2(new_n679), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n659), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n682), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n684), .A2(new_n680), .A3(new_n658), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(G229));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G22), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G166), .B2(new_n688), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1971), .ZN(new_n691));
  NOR2_X1   g266(.A1(G16), .A2(G23), .ZN(new_n692));
  INV_X1    g267(.A(G288), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n692), .B1(new_n693), .B2(G16), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT33), .B(G1976), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n694), .B(new_n695), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n688), .A2(G6), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n571), .A2(new_n574), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(new_n688), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT32), .B(G1981), .Z(new_n700));
  XOR2_X1   g275(.A(new_n699), .B(new_n700), .Z(new_n701));
  NOR3_X1   g276(.A1(new_n691), .A2(new_n696), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT34), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G25), .ZN(new_n705));
  OR2_X1    g280(.A1(G95), .A2(G2105), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n706), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n707));
  INV_X1    g282(.A(G131), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n466), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G119), .B2(new_n486), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n705), .B1(new_n710), .B2(new_n704), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT35), .B(G1991), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT88), .ZN(new_n716));
  MUX2_X1   g291(.A(G24), .B(G290), .S(G16), .Z(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n717), .B2(G1986), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G1986), .B2(new_n717), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n703), .A2(new_n715), .A3(new_n719), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT36), .Z(new_n721));
  INV_X1    g296(.A(G299), .ZN(new_n722));
  OAI21_X1  g297(.A(KEYINPUT23), .B1(new_n722), .B2(new_n688), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n688), .A2(G20), .ZN(new_n724));
  MUX2_X1   g299(.A(new_n723), .B(KEYINPUT23), .S(new_n724), .Z(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(G1956), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(G1956), .ZN(new_n727));
  INV_X1    g302(.A(G2090), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n704), .A2(G35), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G162), .B2(new_n704), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT29), .Z(new_n731));
  OAI211_X1 g306(.A(new_n726), .B(new_n727), .C1(new_n728), .C2(new_n731), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT96), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n704), .A2(G26), .ZN(new_n734));
  OR2_X1    g309(.A1(G104), .A2(G2105), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n735), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT90), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n486), .A2(G128), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n467), .A2(G140), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n734), .B1(new_n741), .B2(new_n704), .ZN(new_n742));
  MUX2_X1   g317(.A(new_n734), .B(new_n742), .S(KEYINPUT28), .Z(new_n743));
  INV_X1    g318(.A(G2067), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n688), .A2(G19), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n542), .B2(new_n688), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1341), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n688), .A2(G4), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n592), .B2(new_n688), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT89), .B(G1348), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n748), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n745), .B(new_n753), .C1(new_n751), .C2(new_n752), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT91), .ZN(new_n755));
  NOR2_X1   g330(.A1(G16), .A2(G21), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G168), .B2(G16), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT95), .B(G1966), .Z(new_n758));
  XOR2_X1   g333(.A(KEYINPUT27), .B(G1996), .Z(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT94), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  OR2_X1    g336(.A1(G29), .A2(G32), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT26), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n765), .A2(new_n766), .B1(G105), .B2(new_n469), .ZN(new_n767));
  INV_X1    g342(.A(G141), .ZN(new_n768));
  INV_X1    g343(.A(G129), .ZN(new_n769));
  OAI221_X1 g344(.A(new_n767), .B1(new_n466), .B2(new_n768), .C1(new_n769), .C2(new_n485), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n762), .B1(new_n770), .B2(new_n704), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n757), .A2(new_n758), .B1(new_n761), .B2(new_n771), .ZN(new_n772));
  AND2_X1   g347(.A1(KEYINPUT24), .A2(G34), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n704), .B1(KEYINPUT24), .B2(G34), .ZN(new_n774));
  OAI22_X1  g349(.A1(G160), .A2(new_n704), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n775), .A2(G2084), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(G2084), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT31), .B(G11), .ZN(new_n778));
  INV_X1    g353(.A(G28), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n779), .A2(KEYINPUT30), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT30), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n704), .B1(new_n781), .B2(G28), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n778), .B1(new_n780), .B2(new_n782), .C1(new_n616), .C2(new_n704), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n776), .A2(new_n777), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n704), .A2(G27), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G164), .B2(new_n704), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(G2078), .Z(new_n787));
  NAND3_X1  g362(.A1(new_n772), .A2(new_n784), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n757), .A2(new_n758), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n688), .A2(G5), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G171), .B2(new_n688), .ZN(new_n791));
  OAI22_X1  g366(.A1(new_n791), .A2(G1961), .B1(new_n761), .B2(new_n771), .ZN(new_n792));
  AOI211_X1 g367(.A(new_n789), .B(new_n792), .C1(G1961), .C2(new_n791), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT93), .ZN(new_n794));
  OAI22_X1  g369(.A1(new_n794), .A2(G2072), .B1(G29), .B2(G33), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n469), .A2(G103), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT25), .Z(new_n797));
  NAND2_X1  g372(.A1(new_n467), .A2(G139), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n607), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n797), .B(new_n798), .C1(new_n459), .C2(new_n799), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT92), .Z(new_n801));
  AOI21_X1  g376(.A(new_n795), .B1(new_n801), .B2(G29), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n794), .A2(G2072), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n793), .A2(new_n804), .ZN(new_n805));
  AOI211_X1 g380(.A(new_n788), .B(new_n805), .C1(new_n728), .C2(new_n731), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n733), .A2(new_n755), .A3(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(KEYINPUT97), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(KEYINPUT97), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n721), .B1(new_n808), .B2(new_n809), .ZN(G311));
  INV_X1    g385(.A(G311), .ZN(G150));
  NAND2_X1  g386(.A1(new_n519), .A2(G93), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT98), .B(G55), .Z(new_n814));
  OAI221_X1 g389(.A(new_n812), .B1(new_n507), .B2(new_n813), .C1(new_n512), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G860), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT37), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n592), .A2(G559), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT38), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n601), .B(new_n815), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT39), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(KEYINPUT99), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(G860), .B1(new_n821), .B2(new_n822), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n823), .B2(KEYINPUT99), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n817), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT100), .Z(G145));
  XOR2_X1   g404(.A(new_n616), .B(G162), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n479), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n498), .B(new_n770), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n740), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(new_n800), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT101), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT101), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n833), .A2(new_n836), .A3(new_n800), .ZN(new_n837));
  INV_X1    g412(.A(new_n833), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(new_n801), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n835), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n486), .A2(G130), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n467), .A2(G142), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT102), .ZN(new_n844));
  INV_X1    g419(.A(G118), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n843), .A2(new_n844), .B1(new_n845), .B2(G2105), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n844), .B2(new_n843), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n841), .A2(new_n842), .A3(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n840), .A2(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n710), .B(new_n609), .Z(new_n851));
  NAND4_X1  g426(.A1(new_n835), .A2(new_n839), .A3(new_n848), .A4(new_n837), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n851), .B1(new_n850), .B2(new_n852), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n831), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(G37), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n850), .A2(new_n852), .ZN(new_n858));
  INV_X1    g433(.A(new_n851), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n831), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT103), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT103), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n860), .A2(new_n865), .A3(new_n861), .A4(new_n862), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n857), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT40), .Z(G395));
  INV_X1    g443(.A(KEYINPUT104), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n820), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n604), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n603), .A2(new_n722), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n592), .A2(G299), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT41), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n872), .A2(KEYINPUT41), .A3(new_n873), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n871), .A2(new_n878), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n879), .A2(KEYINPUT105), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(KEYINPUT105), .ZN(new_n881));
  INV_X1    g456(.A(new_n874), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n871), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT107), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(G303), .B(new_n698), .ZN(new_n888));
  XNOR2_X1  g463(.A(G290), .B(G288), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n889), .A2(KEYINPUT106), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(KEYINPUT106), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n891), .A2(new_n888), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n895), .B1(KEYINPUT107), .B2(KEYINPUT42), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n885), .A2(new_n886), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n880), .A2(new_n897), .A3(new_n881), .A4(new_n883), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n887), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n896), .B1(new_n887), .B2(new_n898), .ZN(new_n900));
  OAI21_X1  g475(.A(G868), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n815), .A2(new_n595), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(G295));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n902), .ZN(G331));
  NAND3_X1  g479(.A1(new_n876), .A2(KEYINPUT109), .A3(new_n877), .ZN(new_n905));
  XNOR2_X1  g480(.A(G171), .B(G286), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(new_n820), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT109), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n874), .A2(new_n909), .A3(new_n875), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n905), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n907), .A2(new_n874), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(KEYINPUT110), .A3(new_n912), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n913), .B(new_n894), .C1(KEYINPUT110), .C2(new_n911), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n878), .A2(new_n908), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n912), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n856), .B1(new_n916), .B2(new_n894), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  XOR2_X1   g493(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n914), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n916), .A2(new_n894), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n919), .B1(new_n922), .B2(new_n917), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n922), .A2(new_n917), .A3(new_n919), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n914), .A2(new_n918), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n925), .B1(KEYINPUT43), .B2(new_n926), .ZN(new_n927));
  MUX2_X1   g502(.A(new_n924), .B(new_n927), .S(KEYINPUT44), .Z(G397));
  INV_X1    g503(.A(KEYINPUT126), .ZN(new_n929));
  INV_X1    g504(.A(G1384), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n460), .B1(new_n461), .B2(G2104), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n473), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n932), .A2(G138), .A3(new_n459), .A4(new_n462), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n491), .B1(new_n933), .B2(KEYINPUT4), .ZN(new_n934));
  INV_X1    g509(.A(G126), .ZN(new_n935));
  OAI22_X1  g510(.A1(new_n485), .A2(new_n935), .B1(new_n494), .B2(new_n495), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n930), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n468), .A2(new_n471), .A3(new_n478), .A4(G40), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n740), .B(G2067), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n770), .B(G1996), .ZN(new_n944));
  OR2_X1    g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n710), .B(new_n712), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G1986), .ZN(new_n948));
  XNOR2_X1  g523(.A(G290), .B(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n942), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n940), .B1(new_n937), .B2(KEYINPUT50), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT50), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n952), .B(new_n930), .C1(new_n934), .C2(new_n936), .ZN(new_n953));
  XNOR2_X1  g528(.A(KEYINPUT116), .B(G2084), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT117), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT117), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n951), .A2(new_n957), .A3(new_n953), .A4(new_n954), .ZN(new_n958));
  AOI21_X1  g533(.A(G1384), .B1(new_n493), .B2(new_n497), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT45), .ZN(new_n960));
  INV_X1    g535(.A(new_n940), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(new_n939), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n758), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n956), .A2(new_n958), .A3(new_n964), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n965), .A2(G8), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(G286), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n956), .A2(new_n964), .A3(G168), .A4(new_n958), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT51), .B1(new_n968), .B2(G8), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT122), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n968), .A2(G8), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n969), .A2(KEYINPUT122), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n967), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n962), .A2(G2078), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT53), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n961), .B1(new_n959), .B2(new_n952), .ZN(new_n978));
  INV_X1    g553(.A(new_n953), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT118), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT118), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n951), .A2(new_n981), .A3(new_n953), .ZN(new_n982));
  AOI21_X1  g557(.A(G1961), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(G171), .B1(new_n977), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT54), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n977), .A2(G171), .A3(new_n983), .ZN(new_n987));
  OR3_X1    g562(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G1971), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n962), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n951), .A2(new_n953), .ZN(new_n991));
  XNOR2_X1  g566(.A(KEYINPUT111), .B(G2090), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n996));
  INV_X1    g571(.A(G8), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n996), .B1(G166), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(G303), .A2(G8), .A3(new_n1000), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n990), .B(KEYINPUT112), .C1(new_n991), .C2(new_n992), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n995), .A2(G8), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT49), .ZN(new_n1005));
  NAND3_X1  g580(.A1(G305), .A2(new_n1005), .A3(G1981), .ZN(new_n1006));
  INV_X1    g581(.A(G1981), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT49), .B1(new_n698), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n1010));
  NOR2_X1   g585(.A1(G305), .A2(G1981), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1009), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n937), .A2(new_n940), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1014), .A2(new_n997), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1008), .B(new_n1006), .C1(new_n1011), .C2(KEYINPUT114), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n693), .A2(G1976), .ZN(new_n1018));
  INV_X1    g593(.A(G1976), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT52), .B1(G288), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1015), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT52), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1017), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n953), .B1(new_n951), .B2(KEYINPUT115), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n1026));
  AOI211_X1 g601(.A(new_n1026), .B(new_n940), .C1(new_n937), .C2(KEYINPUT50), .ZN(new_n1027));
  OR3_X1    g602(.A1(new_n1025), .A2(new_n1027), .A3(new_n992), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n997), .B1(new_n1028), .B2(new_n990), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1004), .B(new_n1024), .C1(new_n1002), .C2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n986), .B1(new_n985), .B2(new_n987), .ZN(new_n1032));
  AND4_X1   g607(.A1(new_n975), .A2(new_n988), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1348), .B1(new_n980), .B2(new_n982), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1014), .A2(new_n744), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1034), .A2(KEYINPUT119), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n1038));
  INV_X1    g613(.A(G1348), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n951), .A2(new_n981), .A3(new_n953), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n981), .B1(new_n951), .B2(new_n953), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1038), .B1(new_n1042), .B2(new_n1035), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1037), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT60), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT119), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1042), .A2(new_n1038), .A3(new_n1035), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n603), .B1(new_n1049), .B2(KEYINPUT60), .ZN(new_n1050));
  AOI211_X1 g625(.A(new_n1045), .B(new_n592), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1046), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT58), .B(G1341), .ZN(new_n1053));
  OAI22_X1  g628(.A1(new_n962), .A2(G1996), .B1(new_n1014), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n542), .ZN(new_n1055));
  XOR2_X1   g630(.A(new_n1055), .B(KEYINPUT59), .Z(new_n1056));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n1058));
  XNOR2_X1  g633(.A(G299), .B(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1956), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT56), .B(G2072), .Z(new_n1062));
  OR2_X1    g637(.A1(new_n962), .A2(new_n1062), .ZN(new_n1063));
  AOI211_X1 g638(.A(new_n1057), .B(new_n1059), .C1(new_n1061), .C2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(G299), .B(KEYINPUT57), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n979), .B1(new_n978), .B2(new_n1026), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n951), .A2(KEYINPUT115), .ZN(new_n1067));
  AOI21_X1  g642(.A(G1956), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n962), .A2(new_n1062), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1065), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1061), .A2(new_n1059), .A3(new_n1063), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1064), .B1(new_n1072), .B2(KEYINPUT61), .ZN(new_n1073));
  NOR2_X1   g648(.A1(KEYINPUT120), .A2(KEYINPUT61), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1070), .A2(new_n1071), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1056), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1052), .A2(new_n1076), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1068), .A2(new_n1065), .A3(new_n1069), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(new_n603), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1044), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1070), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT121), .B1(new_n1077), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n1084));
  AOI211_X1 g659(.A(new_n1084), .B(new_n1081), .C1(new_n1052), .C2(new_n1076), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1033), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT63), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n966), .A2(G168), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1087), .B1(new_n1030), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1088), .A2(new_n1087), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n995), .A2(G8), .A3(new_n1003), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1002), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1090), .A2(new_n1004), .A3(new_n1024), .A4(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1089), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1004), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n1024), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1017), .A2(new_n1019), .A3(new_n693), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1015), .B1(new_n1098), .B2(new_n1011), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1095), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1031), .A2(new_n985), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n972), .A2(new_n971), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(KEYINPUT122), .B2(new_n969), .ZN(new_n1105));
  INV_X1    g680(.A(new_n974), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1105), .A2(new_n1106), .B1(G286), .B2(new_n966), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1103), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n975), .A2(KEYINPUT62), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1102), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n950), .B1(new_n1086), .B2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n947), .A2(new_n942), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n941), .A2(new_n948), .A3(new_n580), .A4(new_n578), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1114), .B(KEYINPUT124), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1113), .B1(KEYINPUT48), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(KEYINPUT48), .B2(new_n1116), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT46), .ZN(new_n1119));
  OR3_X1    g694(.A1(new_n942), .A2(new_n1119), .A3(G1996), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n941), .B1(new_n943), .B2(new_n770), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1119), .B1(new_n942), .B2(G1996), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  XOR2_X1   g699(.A(KEYINPUT123), .B(KEYINPUT47), .Z(new_n1125));
  OR2_X1    g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n710), .A2(new_n712), .ZN(new_n1127));
  OAI22_X1  g702(.A1(new_n945), .A2(new_n1127), .B1(G2067), .B2(new_n740), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n941), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1118), .A2(new_n1126), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  XOR2_X1   g706(.A(new_n1131), .B(KEYINPUT125), .Z(new_n1132));
  OAI21_X1  g707(.A(new_n929), .B1(new_n1112), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1132), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1100), .B1(new_n1089), .B2(new_n1094), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1031), .B(new_n985), .C1(new_n975), .C2(KEYINPUT62), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1049), .A2(KEYINPUT60), .ZN(new_n1139));
  OAI21_X1  g714(.A(KEYINPUT60), .B1(new_n1037), .B2(new_n1043), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n592), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1049), .A2(KEYINPUT60), .A3(new_n603), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1139), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1059), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT61), .B1(new_n1078), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1064), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1145), .A2(new_n1075), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1056), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1082), .B1(new_n1143), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n1084), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1077), .A2(KEYINPUT121), .A3(new_n1082), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1138), .B1(new_n1153), .B2(new_n1033), .ZN(new_n1154));
  OAI211_X1 g729(.A(KEYINPUT126), .B(new_n1134), .C1(new_n1154), .C2(new_n950), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1133), .A2(new_n1155), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g731(.A1(new_n656), .A2(new_n637), .A3(G319), .ZN(new_n1158));
  NAND3_X1  g732(.A1(new_n683), .A2(new_n685), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g733(.A(new_n1159), .B1(new_n923), .B2(new_n921), .ZN(new_n1160));
  INV_X1    g734(.A(new_n867), .ZN(new_n1161));
  INV_X1    g735(.A(KEYINPUT127), .ZN(new_n1162));
  NAND3_X1  g736(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  AND3_X1   g737(.A1(new_n683), .A2(new_n685), .A3(new_n1158), .ZN(new_n1164));
  NAND2_X1  g738(.A1(new_n1164), .A2(new_n924), .ZN(new_n1165));
  OAI21_X1  g739(.A(KEYINPUT127), .B1(new_n1165), .B2(new_n867), .ZN(new_n1166));
  NAND2_X1  g740(.A1(new_n1163), .A2(new_n1166), .ZN(G308));
  NAND2_X1  g741(.A1(new_n1160), .A2(new_n1161), .ZN(G225));
endmodule


