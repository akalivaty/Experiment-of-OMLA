//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT12), .ZN(new_n206));
  NAND2_X1  g005(.A1(G229gat), .A2(G233gat), .ZN(new_n207));
  XOR2_X1   g006(.A(new_n207), .B(KEYINPUT13), .Z(new_n208));
  INV_X1    g007(.A(KEYINPUT91), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT14), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(KEYINPUT91), .A2(KEYINPUT14), .ZN(new_n212));
  OAI22_X1  g011(.A1(new_n211), .A2(new_n212), .B1(G29gat), .B2(G36gat), .ZN(new_n213));
  INV_X1    g012(.A(G29gat), .ZN(new_n214));
  INV_X1    g013(.A(G36gat), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n214), .B(new_n215), .C1(new_n209), .C2(new_n210), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT92), .ZN(new_n218));
  AOI22_X1  g017(.A1(new_n217), .A2(new_n218), .B1(G29gat), .B2(G36gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(new_n218), .B2(new_n217), .ZN(new_n220));
  INV_X1    g019(.A(G50gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G43gat), .ZN(new_n222));
  INV_X1    g021(.A(G43gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G50gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n224), .A3(KEYINPUT15), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n220), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n225), .B(KEYINPUT93), .ZN(new_n228));
  NAND2_X1  g027(.A1(G29gat), .A2(G36gat), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n228), .A2(new_n217), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT94), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n222), .A2(new_n224), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT15), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n232), .B(new_n233), .C1(new_n231), .C2(new_n222), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT95), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n234), .B(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n230), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n227), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G15gat), .B(G22gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT16), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(G1gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(G1gat), .B2(new_n239), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(G8gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n226), .A2(new_n220), .B1(new_n230), .B2(new_n236), .ZN(new_n245));
  INV_X1    g044(.A(new_n243), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n208), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n207), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT17), .B1(new_n227), .B2(new_n237), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n246), .B1(new_n250), .B2(KEYINPUT96), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT96), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT17), .B1(new_n243), .B2(new_n252), .ZN(new_n253));
  OR2_X1    g052(.A1(new_n238), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n249), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n248), .B1(new_n255), .B2(KEYINPUT18), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n238), .A2(new_n253), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n252), .B1(new_n245), .B2(KEYINPUT17), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n257), .B1(new_n258), .B2(new_n246), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT18), .ZN(new_n260));
  NOR3_X1   g059(.A1(new_n259), .A2(new_n260), .A3(new_n249), .ZN(new_n261));
  OAI211_X1 g060(.A(KEYINPUT90), .B(new_n206), .C1(new_n256), .C2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n260), .B1(new_n259), .B2(new_n249), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n255), .A2(KEYINPUT18), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n265), .A3(new_n248), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n206), .B1(new_n266), .B2(KEYINPUT90), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT85), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT36), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT34), .ZN(new_n272));
  NOR2_X1   g071(.A1(KEYINPUT69), .A2(KEYINPUT28), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT27), .B(G183gat), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n275), .B2(G190gat), .ZN(new_n276));
  INV_X1    g075(.A(G190gat), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n274), .B(new_n277), .C1(KEYINPUT69), .C2(KEYINPUT28), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G169gat), .A2(G176gat), .ZN(new_n280));
  INV_X1    g079(.A(G169gat), .ZN(new_n281));
  INV_X1    g080(.A(G176gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT26), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n283), .B1(KEYINPUT65), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT26), .B1(new_n287), .B2(new_n284), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n280), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n279), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT23), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n283), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT23), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n293), .A2(new_n280), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT24), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n290), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT64), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n301));
  OR2_X1    g100(.A1(G183gat), .A2(G190gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n290), .A2(KEYINPUT64), .A3(new_n297), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n300), .A2(new_n301), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT25), .B1(new_n296), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT25), .B1(new_n294), .B2(KEYINPUT23), .ZN(new_n306));
  NAND4_X1  g105(.A1(KEYINPUT67), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n298), .A2(new_n307), .A3(new_n302), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT67), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n301), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n306), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT66), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n287), .A2(KEYINPUT23), .ZN(new_n314));
  NOR3_X1   g113(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n313), .B(new_n280), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT65), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n318), .A2(new_n281), .A3(new_n282), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n319), .A2(KEYINPUT23), .A3(new_n287), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n313), .B1(new_n320), .B2(new_n280), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n312), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT68), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n305), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT25), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n325), .B1(new_n283), .B2(new_n292), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n298), .A2(new_n302), .A3(new_n307), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n326), .B1(new_n327), .B2(new_n310), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n280), .B1(new_n314), .B2(new_n315), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT66), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n328), .B1(new_n330), .B2(new_n316), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT68), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n291), .B1(new_n324), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n334));
  OR2_X1    g133(.A1(KEYINPUT72), .A2(G127gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(KEYINPUT72), .A2(G127gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(G134gat), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G127gat), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT71), .B1(new_n338), .B2(G134gat), .ZN(new_n339));
  OR3_X1    g138(.A1(new_n338), .A2(KEYINPUT71), .A3(G134gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n337), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G113gat), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n344), .A2(G120gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(G120gat), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT1), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n337), .A2(new_n340), .A3(KEYINPUT73), .A4(new_n339), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n343), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G127gat), .B(G134gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n333), .A2(new_n334), .A3(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n279), .A2(new_n289), .A3(new_n290), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n296), .A2(new_n304), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n325), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n357), .B1(new_n331), .B2(KEYINPUT68), .ZN(new_n358));
  AOI211_X1 g157(.A(new_n323), .B(new_n328), .C1(new_n316), .C2(new_n330), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n355), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n347), .B1(new_n341), .B2(new_n342), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n361), .A2(new_n349), .B1(new_n347), .B2(new_n351), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT74), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n353), .A2(new_n334), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n360), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n354), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G227gat), .A2(G233gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n272), .B1(new_n368), .B2(KEYINPUT77), .ZN(new_n369));
  INV_X1    g168(.A(new_n367), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n370), .B1(new_n354), .B2(new_n365), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT77), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT34), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n354), .A2(new_n365), .A3(new_n370), .ZN(new_n375));
  XNOR2_X1  g174(.A(G15gat), .B(G43gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(KEYINPUT75), .ZN(new_n377));
  XNOR2_X1  g176(.A(G71gat), .B(G99gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT33), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n375), .A2(KEYINPUT32), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT76), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT76), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n375), .A2(new_n383), .A3(KEYINPUT32), .A4(new_n380), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n375), .A2(KEYINPUT32), .ZN(new_n386));
  INV_X1    g185(.A(new_n375), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n386), .B(new_n379), .C1(new_n387), .C2(KEYINPUT33), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n374), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n369), .ZN(new_n390));
  INV_X1    g189(.A(new_n373), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n385), .A2(new_n388), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n271), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n385), .A2(new_n388), .ZN(new_n394));
  INV_X1    g193(.A(new_n374), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n374), .A2(new_n385), .A3(new_n388), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(KEYINPUT36), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G78gat), .B(G106gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(G22gat), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G197gat), .B(G204gat), .ZN(new_n403));
  INV_X1    g202(.A(G211gat), .ZN(new_n404));
  INV_X1    g203(.A(G218gat), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n403), .B1(KEYINPUT22), .B2(new_n406), .ZN(new_n407));
  XOR2_X1   g206(.A(G211gat), .B(G218gat), .Z(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT29), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT3), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OR2_X1    g211(.A1(KEYINPUT81), .A2(G141gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(KEYINPUT81), .A2(G141gat), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n413), .A2(G148gat), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G148gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(G141gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(G155gat), .A2(G162gat), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT2), .ZN(new_n419));
  INV_X1    g218(.A(G155gat), .ZN(new_n420));
  INV_X1    g219(.A(G162gat), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n415), .A2(new_n417), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n420), .A2(new_n421), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n418), .ZN(new_n425));
  XOR2_X1   g224(.A(G141gat), .B(G148gat), .Z(new_n426));
  AOI21_X1  g225(.A(new_n425), .B1(new_n426), .B2(new_n419), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n412), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT3), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n410), .B1(new_n431), .B2(new_n411), .ZN(new_n432));
  OAI211_X1 g231(.A(G228gat), .B(G233gat), .C1(new_n429), .C2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n432), .ZN(new_n434));
  NAND2_X1  g233(.A1(G228gat), .A2(G233gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n426), .A2(new_n419), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n424), .A2(new_n418), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n415), .A2(new_n417), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n422), .A2(new_n418), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT82), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT82), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n434), .B(new_n435), .C1(new_n445), .C2(new_n412), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT31), .B(G50gat), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n448), .B1(new_n433), .B2(new_n446), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n402), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n451), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(new_n401), .A3(new_n449), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(G8gat), .B(G36gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(G64gat), .B(G92gat), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n457), .B(new_n458), .Z(new_n459));
  NAND2_X1  g258(.A1(G226gat), .A2(G233gat), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n360), .B2(new_n411), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n333), .A2(new_n460), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT78), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n460), .B1(new_n333), .B2(KEYINPUT29), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT78), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n410), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT79), .B1(new_n333), .B2(new_n460), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT79), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n360), .A2(new_n470), .A3(new_n461), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n465), .A2(new_n469), .A3(new_n410), .A4(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT80), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(new_n473), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n459), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n360), .A2(new_n461), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n466), .B1(new_n465), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n462), .A2(KEYINPUT78), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n409), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n470), .B1(new_n360), .B2(new_n461), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n462), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n483), .A2(KEYINPUT80), .A3(new_n410), .A4(new_n471), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n481), .A2(new_n484), .A3(new_n476), .A4(new_n459), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT30), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n477), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n442), .A2(new_n362), .A3(KEYINPUT4), .A4(new_n444), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT3), .B1(new_n423), .B2(new_n427), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n353), .A2(new_n431), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n350), .A2(new_n352), .A3(new_n428), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G225gat), .A2(G233gat), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n489), .A2(new_n491), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT5), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n353), .A2(new_n441), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n492), .ZN(new_n499));
  INV_X1    g298(.A(new_n495), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n491), .A2(new_n497), .A3(new_n495), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n442), .A2(new_n362), .A3(new_n493), .A4(new_n444), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n496), .A2(new_n501), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  XOR2_X1   g306(.A(G1gat), .B(G29gat), .Z(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G57gat), .B(G85gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT6), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT84), .B1(new_n507), .B2(new_n512), .ZN(new_n515));
  AOI21_X1  g314(.A(KEYINPUT6), .B1(new_n507), .B2(new_n512), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n496), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n503), .A2(new_n506), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT84), .ZN(new_n520));
  INV_X1    g319(.A(new_n512), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n515), .A2(new_n516), .A3(new_n522), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n514), .A2(new_n523), .B1(new_n485), .B2(new_n486), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n456), .B1(new_n488), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n270), .B1(new_n399), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n514), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n485), .A2(new_n486), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n481), .A2(new_n484), .A3(new_n476), .ZN(new_n530));
  INV_X1    g329(.A(new_n459), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(new_n486), .B2(new_n485), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n455), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n534), .A2(KEYINPUT85), .A3(new_n398), .A4(new_n393), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n506), .A2(new_n491), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n536), .A2(KEYINPUT86), .A3(new_n500), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT86), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n431), .A2(new_n490), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n504), .A2(new_n505), .B1(new_n539), .B2(new_n353), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n538), .B1(new_n540), .B2(new_n495), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT39), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n521), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n498), .A2(new_n495), .A3(new_n492), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n537), .A2(new_n541), .A3(KEYINPUT39), .A4(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(KEYINPUT40), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT87), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n519), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n507), .A2(KEYINPUT87), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n549), .A2(new_n550), .A3(new_n521), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT40), .B1(new_n544), .B2(new_n546), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n475), .A2(KEYINPUT30), .A3(new_n476), .A4(new_n459), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n555), .A2(new_n532), .A3(new_n528), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT38), .ZN(new_n558));
  XOR2_X1   g357(.A(KEYINPUT88), .B(KEYINPUT37), .Z(new_n559));
  NAND4_X1  g358(.A1(new_n481), .A2(new_n484), .A3(new_n476), .A4(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n560), .A2(new_n531), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n530), .A2(KEYINPUT37), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n465), .A2(new_n469), .A3(new_n409), .A4(new_n471), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n564), .A2(KEYINPUT37), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n410), .B1(new_n479), .B2(new_n480), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT38), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n567), .A2(new_n560), .A3(new_n531), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n551), .A2(new_n516), .B1(KEYINPUT6), .B2(new_n513), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n569), .A3(new_n485), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n557), .B(new_n456), .C1(new_n563), .C2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n526), .A2(new_n535), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n529), .A2(new_n533), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n455), .B1(new_n396), .B2(new_n397), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT35), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT89), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n389), .A2(new_n392), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT89), .B1(new_n396), .B2(new_n397), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n556), .ZN(new_n581));
  NOR3_X1   g380(.A1(new_n455), .A2(new_n569), .A3(KEYINPUT35), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI22_X1  g382(.A1(new_n575), .A2(new_n576), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n269), .B1(new_n572), .B2(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G183gat), .B(G211gat), .Z(new_n586));
  INV_X1    g385(.A(G71gat), .ZN(new_n587));
  INV_X1    g386(.A(G78gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(G71gat), .A2(G78gat), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n591));
  OAI22_X1  g390(.A1(new_n589), .A2(new_n590), .B1(new_n591), .B2(KEYINPUT97), .ZN(new_n592));
  INV_X1    g391(.A(G57gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(G64gat), .ZN(new_n594));
  INV_X1    g393(.A(G64gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(G57gat), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n591), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n592), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT98), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n599), .A2(KEYINPUT21), .ZN(new_n600));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n600), .A2(new_n601), .ZN(new_n603));
  OAI21_X1  g402(.A(G127gat), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NOR3_X1   g404(.A1(new_n602), .A2(new_n603), .A3(G127gat), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n586), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n606), .ZN(new_n608));
  INV_X1    g407(.A(new_n586), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n608), .A2(new_n609), .A3(new_n604), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n243), .B1(new_n599), .B2(KEYINPUT21), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n612), .B(KEYINPUT99), .Z(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(new_n420), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n611), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n607), .A2(new_n610), .A3(new_n616), .A4(new_n617), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G85gat), .A2(G92gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT7), .ZN(new_n624));
  NAND2_X1  g423(.A1(G99gat), .A2(G106gat), .ZN(new_n625));
  INV_X1    g424(.A(G85gat), .ZN(new_n626));
  INV_X1    g425(.A(G92gat), .ZN(new_n627));
  AOI22_X1  g426(.A1(KEYINPUT8), .A2(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G99gat), .B(G106gat), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n629), .B(new_n630), .Z(new_n631));
  AOI21_X1  g430(.A(new_n631), .B1(new_n227), .B2(new_n237), .ZN(new_n632));
  NAND3_X1  g431(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT100), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n636), .B(new_n633), .C1(new_n245), .C2(new_n631), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n629), .B(new_n630), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n250), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n245), .A2(KEYINPUT17), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n635), .A2(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G190gat), .B(G218gat), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT101), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(G134gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(new_n421), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT102), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n641), .B(new_n642), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n644), .A2(new_n651), .A3(new_n647), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n649), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n650), .ZN(new_n654));
  INV_X1    g453(.A(new_n652), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n651), .B1(new_n644), .B2(new_n647), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(G230gat), .A2(G233gat), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT103), .B(KEYINPUT10), .Z(new_n659));
  XOR2_X1   g458(.A(new_n592), .B(new_n597), .Z(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT98), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT98), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n598), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n661), .A2(new_n631), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n638), .A2(new_n660), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n659), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n638), .A2(KEYINPUT10), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n599), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n658), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n664), .A2(new_n665), .ZN(new_n671));
  INV_X1    g470(.A(new_n658), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(G120gat), .B(G148gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(G176gat), .B(G204gat), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n675), .B(new_n676), .Z(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n670), .A2(new_n673), .A3(new_n677), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n622), .A2(new_n653), .A3(new_n657), .A4(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n585), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(new_n527), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(G1gat), .Z(G1324gat));
  NAND3_X1  g486(.A1(new_n585), .A2(new_n556), .A3(new_n684), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n688), .A2(G8gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT16), .B(G8gat), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT42), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(KEYINPUT42), .B2(new_n691), .ZN(G1325gat));
  INV_X1    g492(.A(new_n399), .ZN(new_n694));
  OAI21_X1  g493(.A(G15gat), .B1(new_n685), .B2(new_n694), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n580), .A2(G15gat), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n695), .B1(new_n685), .B2(new_n696), .ZN(G1326gat));
  NOR2_X1   g496(.A1(new_n685), .A2(new_n456), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT43), .B(G22gat), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  NAND2_X1  g499(.A1(new_n657), .A2(new_n653), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n702), .A2(new_n622), .A3(new_n681), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n585), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n527), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n214), .ZN(new_n706));
  OR3_X1    g505(.A1(new_n704), .A2(KEYINPUT104), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT104), .B1(new_n704), .B2(new_n706), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n707), .A2(KEYINPUT45), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT45), .B1(new_n707), .B2(new_n708), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n621), .B(KEYINPUT105), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n712), .A2(new_n269), .A3(new_n681), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n701), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n456), .B1(new_n563), .B2(new_n570), .ZN(new_n716));
  INV_X1    g515(.A(new_n557), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n534), .A2(new_n398), .A3(new_n393), .ZN(new_n719));
  OAI21_X1  g518(.A(KEYINPUT106), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n719), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(new_n571), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n715), .B1(new_n724), .B2(new_n584), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n572), .A2(new_n584), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n714), .B1(new_n726), .B2(new_n701), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n713), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  OAI211_X1 g530(.A(KEYINPUT107), .B(new_n713), .C1(new_n725), .C2(new_n727), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n731), .A2(new_n733), .A3(new_n527), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n711), .B1(new_n734), .B2(new_n214), .ZN(G1328gat));
  NOR3_X1   g534(.A1(new_n704), .A2(G36gat), .A3(new_n581), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT46), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(KEYINPUT108), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n739));
  OR2_X1    g538(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n731), .A2(new_n733), .A3(new_n581), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n738), .B(new_n740), .C1(new_n741), .C2(new_n215), .ZN(G1329gat));
  OAI21_X1  g541(.A(G43gat), .B1(new_n728), .B2(new_n694), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n704), .A2(G43gat), .A3(new_n580), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n743), .A2(KEYINPUT47), .A3(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n730), .A2(new_n399), .A3(new_n732), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n744), .B1(new_n747), .B2(G43gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n748), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g548(.A(G50gat), .B1(new_n728), .B2(new_n456), .ZN(new_n750));
  AOI21_X1  g549(.A(KEYINPUT109), .B1(new_n585), .B2(new_n703), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n221), .B(new_n455), .C1(new_n704), .C2(new_n752), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n750), .B(KEYINPUT48), .C1(new_n751), .C2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n753), .A2(new_n751), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n730), .A2(new_n455), .A3(new_n732), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n755), .B1(new_n756), .B2(G50gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n754), .B1(new_n757), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g557(.A1(new_n718), .A2(KEYINPUT106), .A3(new_n719), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n722), .B1(new_n721), .B2(new_n571), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n584), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR4_X1   g560(.A1(new_n701), .A2(new_n621), .A3(new_n268), .A4(new_n682), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(new_n527), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(new_n593), .ZN(G1332gat));
  NOR2_X1   g564(.A1(new_n763), .A2(new_n581), .ZN(new_n766));
  NOR2_X1   g565(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n767));
  AND2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n766), .B2(new_n767), .ZN(G1333gat));
  XOR2_X1   g569(.A(new_n580), .B(KEYINPUT110), .Z(new_n771));
  OAI21_X1  g570(.A(new_n587), .B1(new_n763), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n399), .A2(G71gat), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n763), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g574(.A1(new_n763), .A2(new_n456), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(new_n588), .ZN(G1335gat));
  NOR2_X1   g576(.A1(new_n622), .A2(new_n268), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n681), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(new_n725), .B2(new_n727), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT111), .B1(new_n781), .B2(new_n527), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G85gat), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n781), .A2(KEYINPUT111), .A3(new_n527), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n778), .A2(new_n701), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n761), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n787), .B1(new_n761), .B2(new_n790), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n681), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n705), .A2(new_n626), .ZN(new_n795));
  OAI22_X1  g594(.A1(new_n783), .A2(new_n784), .B1(new_n794), .B2(new_n795), .ZN(G1336gat));
  OAI211_X1 g595(.A(new_n556), .B(new_n780), .C1(new_n725), .C2(new_n727), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(G92gat), .ZN(new_n798));
  XOR2_X1   g597(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n799));
  NAND2_X1  g598(.A1(new_n556), .A2(new_n627), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n798), .B(new_n799), .C1(new_n794), .C2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n797), .A2(new_n802), .A3(G92gat), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n802), .B1(new_n797), .B2(G92gat), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n575), .A2(new_n576), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n580), .A2(new_n583), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n720), .A2(new_n723), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI22_X1  g606(.A1(new_n807), .A2(new_n789), .B1(new_n785), .B2(new_n786), .ZN(new_n808));
  AOI211_X1 g607(.A(new_n682), .B(new_n800), .C1(new_n808), .C2(new_n791), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n803), .A2(new_n804), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n801), .B1(new_n810), .B2(new_n811), .ZN(G1337gat));
  OAI21_X1  g611(.A(G99gat), .B1(new_n781), .B2(new_n694), .ZN(new_n813));
  OR2_X1    g612(.A1(new_n580), .A2(G99gat), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n794), .B2(new_n814), .ZN(G1338gat));
  OAI21_X1  g614(.A(G106gat), .B1(new_n781), .B2(new_n456), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n456), .A2(G106gat), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n681), .B(new_n817), .C1(new_n792), .C2(new_n793), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g619(.A(new_n712), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822));
  XOR2_X1   g621(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n678), .B1(new_n670), .B2(new_n824), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n672), .B(new_n668), .C1(new_n671), .C2(new_n659), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(new_n670), .A3(KEYINPUT54), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT115), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n826), .A2(new_n670), .A3(new_n829), .A4(KEYINPUT54), .ZN(new_n830));
  AOI211_X1 g629(.A(new_n822), .B(new_n825), .C1(new_n828), .C2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n680), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT117), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n825), .B1(new_n828), .B2(new_n830), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT55), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(new_n836), .A3(new_n680), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n834), .A2(KEYINPUT55), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n833), .A2(new_n837), .A3(new_n268), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n259), .A2(new_n249), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n244), .A2(new_n247), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n841), .B1(new_n842), .B2(new_n208), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n205), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n264), .A2(new_n265), .A3(new_n248), .A4(new_n206), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n845), .A3(new_n681), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n846), .B(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n701), .B1(new_n840), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n832), .B1(new_n834), .B2(KEYINPUT55), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n838), .B1(new_n850), .B2(new_n836), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n844), .A2(new_n845), .ZN(new_n852));
  AND4_X1   g651(.A1(new_n701), .A2(new_n851), .A3(new_n833), .A4(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n821), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n683), .A2(new_n268), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n527), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n857), .A2(new_n858), .A3(new_n574), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n858), .B1(new_n857), .B2(new_n574), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n556), .ZN(new_n862));
  AOI21_X1  g661(.A(G113gat), .B1(new_n862), .B2(new_n268), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n854), .A2(new_n856), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n865), .B2(new_n456), .ZN(new_n866));
  AOI211_X1 g665(.A(KEYINPUT119), .B(new_n455), .C1(new_n854), .C2(new_n856), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n581), .A2(new_n705), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n580), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n269), .A2(new_n344), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n863), .B1(new_n872), .B2(new_n873), .ZN(G1340gat));
  OAI211_X1 g673(.A(new_n681), .B(new_n870), .C1(new_n866), .C2(new_n867), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(G120gat), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n682), .A2(G120gat), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n581), .B(new_n877), .C1(new_n859), .C2(new_n860), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT121), .ZN(G1341gat));
  NAND2_X1  g679(.A1(new_n335), .A2(new_n336), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n712), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n870), .B(new_n882), .C1(new_n866), .C2(new_n867), .ZN(new_n883));
  XOR2_X1   g682(.A(new_n883), .B(KEYINPUT122), .Z(new_n884));
  AOI21_X1  g683(.A(new_n881), .B1(new_n862), .B2(new_n622), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(G1342gat));
  OAI21_X1  g685(.A(G134gat), .B1(new_n871), .B2(new_n702), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n702), .A2(G134gat), .A3(new_n556), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  OR3_X1    g688(.A1(new_n861), .A2(KEYINPUT56), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT56), .B1(new_n861), .B2(new_n889), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n887), .A2(new_n890), .A3(new_n891), .ZN(G1343gat));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n865), .A2(new_n893), .A3(new_n455), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n701), .A2(new_n851), .A3(new_n833), .A4(new_n852), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n838), .A2(new_n263), .A3(new_n267), .ZN(new_n896));
  AOI22_X1  g695(.A1(new_n896), .A2(new_n850), .B1(new_n681), .B2(new_n852), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n895), .B1(new_n897), .B2(new_n701), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n855), .B1(new_n898), .B2(new_n621), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT57), .B1(new_n899), .B2(new_n456), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n399), .A2(new_n869), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n894), .A2(new_n900), .A3(new_n268), .A4(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n413), .A2(new_n414), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n902), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n857), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n694), .A2(new_n455), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n909), .B1(new_n857), .B2(new_n907), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n269), .A2(G141gat), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n908), .A2(new_n910), .A3(new_n581), .A4(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n903), .B1(new_n902), .B2(new_n905), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n906), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT58), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT58), .B1(new_n902), .B2(new_n905), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n917), .A2(KEYINPUT125), .A3(new_n912), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT125), .B1(new_n917), .B2(new_n912), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n915), .A2(new_n916), .B1(new_n918), .B2(new_n919), .ZN(G1344gat));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n456), .B1(new_n854), .B2(new_n856), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n922), .A2(KEYINPUT57), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n899), .A2(new_n456), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n924), .A2(KEYINPUT57), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n681), .B(new_n901), .C1(new_n923), .C2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n921), .B1(new_n926), .B2(G148gat), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n894), .A2(new_n900), .A3(new_n901), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n928), .A2(new_n682), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n929), .A2(KEYINPUT59), .A3(new_n416), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n908), .A2(new_n581), .A3(new_n910), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n681), .A2(new_n416), .ZN(new_n932));
  OAI22_X1  g731(.A1(new_n927), .A2(new_n930), .B1(new_n931), .B2(new_n932), .ZN(G1345gat));
  OAI21_X1  g732(.A(G155gat), .B1(new_n928), .B2(new_n821), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n622), .A2(new_n420), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n934), .B1(new_n931), .B2(new_n935), .ZN(G1346gat));
  OAI21_X1  g735(.A(G162gat), .B1(new_n928), .B2(new_n702), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n702), .A2(G162gat), .A3(new_n556), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n908), .A2(new_n910), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(G1347gat));
  AND3_X1   g739(.A1(new_n574), .A2(new_n527), .A3(new_n556), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n865), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(G169gat), .B1(new_n943), .B2(new_n268), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n556), .A2(new_n527), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n771), .A2(new_n945), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n868), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n269), .A2(new_n281), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(G1348gat));
  AOI21_X1  g748(.A(new_n282), .B1(new_n947), .B2(new_n681), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n942), .A2(G176gat), .A3(new_n682), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n950), .A2(new_n951), .ZN(G1349gat));
  OAI211_X1 g751(.A(new_n712), .B(new_n946), .C1(new_n866), .C2(new_n867), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G183gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n943), .A2(new_n274), .A3(new_n622), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g756(.A1(new_n943), .A2(new_n277), .A3(new_n701), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n868), .A2(new_n701), .A3(new_n946), .ZN(new_n959));
  NOR2_X1   g758(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n277), .B1(KEYINPUT126), .B2(KEYINPUT61), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n960), .B1(new_n959), .B2(new_n961), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n958), .B1(new_n962), .B2(new_n963), .ZN(G1351gat));
  NOR2_X1   g763(.A1(new_n399), .A2(new_n945), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n965), .B1(new_n923), .B2(new_n925), .ZN(new_n966));
  INV_X1    g765(.A(G197gat), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n966), .A2(new_n967), .A3(new_n269), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n922), .A2(new_n965), .ZN(new_n969));
  AOI21_X1  g768(.A(G197gat), .B1(new_n969), .B2(new_n268), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n968), .A2(new_n970), .ZN(G1352gat));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n682), .A2(G204gat), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n969), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  XOR2_X1   g773(.A(new_n974), .B(KEYINPUT127), .Z(new_n975));
  OAI21_X1  g774(.A(G204gat), .B1(new_n966), .B2(new_n682), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n969), .A2(new_n973), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT62), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n975), .A2(new_n976), .A3(new_n978), .ZN(G1353gat));
  NAND3_X1  g778(.A1(new_n969), .A2(new_n404), .A3(new_n622), .ZN(new_n980));
  OAI211_X1 g779(.A(new_n622), .B(new_n965), .C1(new_n923), .C2(new_n925), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n981), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n982));
  AOI21_X1  g781(.A(KEYINPUT63), .B1(new_n981), .B2(G211gat), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(G1354gat));
  OAI21_X1  g783(.A(G218gat), .B1(new_n966), .B2(new_n702), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n969), .A2(new_n405), .A3(new_n701), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(G1355gat));
endmodule


